module top (\a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \result[0] , \result[1] , \result[2] , \result[3] , \result[4] , \result[5] , \result[6] , \result[7] , \result[8] , \result[9] , \result[10] , \result[11] , \result[12] , \result[13] , \result[14] , \result[15] , \result[16] , \result[17] , \result[18] , \result[19] , \result[20] , \result[21] , \result[22] , \result[23] , \result[24] , \result[25] , \result[26] , \result[27] , \result[28] , \result[29] , \result[30] , \result[31] );
	input \a[0]  ;
	input \a[1]  ;
	input \a[2]  ;
	input \a[3]  ;
	input \a[4]  ;
	input \a[5]  ;
	input \a[6]  ;
	input \a[7]  ;
	input \a[8]  ;
	input \a[9]  ;
	input \a[10]  ;
	input \a[11]  ;
	input \a[12]  ;
	input \a[13]  ;
	input \a[14]  ;
	input \a[15]  ;
	input \a[16]  ;
	input \a[17]  ;
	input \a[18]  ;
	input \a[19]  ;
	input \a[20]  ;
	input \a[21]  ;
	input \a[22]  ;
	input \a[23]  ;
	input \a[24]  ;
	input \a[25]  ;
	input \a[26]  ;
	input \a[27]  ;
	input \a[28]  ;
	input \a[29]  ;
	input \a[30]  ;
	input \a[31]  ;
	output \result[0]  ;
	output \result[1]  ;
	output \result[2]  ;
	output \result[3]  ;
	output \result[4]  ;
	output \result[5]  ;
	output \result[6]  ;
	output \result[7]  ;
	output \result[8]  ;
	output \result[9]  ;
	output \result[10]  ;
	output \result[11]  ;
	output \result[12]  ;
	output \result[13]  ;
	output \result[14]  ;
	output \result[15]  ;
	output \result[16]  ;
	output \result[17]  ;
	output \result[18]  ;
	output \result[19]  ;
	output \result[20]  ;
	output \result[21]  ;
	output \result[22]  ;
	output \result[23]  ;
	output \result[24]  ;
	output \result[25]  ;
	output \result[26]  ;
	output \result[27]  ;
	output \result[28]  ;
	output \result[29]  ;
	output \result[30]  ;
	output \result[31]  ;
	wire _w16192_ ;
	wire _w16191_ ;
	wire _w16190_ ;
	wire _w16189_ ;
	wire _w16188_ ;
	wire _w16187_ ;
	wire _w16186_ ;
	wire _w16185_ ;
	wire _w16184_ ;
	wire _w16183_ ;
	wire _w16182_ ;
	wire _w16181_ ;
	wire _w16180_ ;
	wire _w16179_ ;
	wire _w16178_ ;
	wire _w16177_ ;
	wire _w16176_ ;
	wire _w16175_ ;
	wire _w16174_ ;
	wire _w16173_ ;
	wire _w16172_ ;
	wire _w16171_ ;
	wire _w16170_ ;
	wire _w16169_ ;
	wire _w16168_ ;
	wire _w16167_ ;
	wire _w16166_ ;
	wire _w16165_ ;
	wire _w16164_ ;
	wire _w16163_ ;
	wire _w16162_ ;
	wire _w16161_ ;
	wire _w16160_ ;
	wire _w16159_ ;
	wire _w16158_ ;
	wire _w16157_ ;
	wire _w16156_ ;
	wire _w16155_ ;
	wire _w16154_ ;
	wire _w16153_ ;
	wire _w16152_ ;
	wire _w16151_ ;
	wire _w16150_ ;
	wire _w16149_ ;
	wire _w16148_ ;
	wire _w16147_ ;
	wire _w16146_ ;
	wire _w16145_ ;
	wire _w16144_ ;
	wire _w16143_ ;
	wire _w16142_ ;
	wire _w16141_ ;
	wire _w16140_ ;
	wire _w16139_ ;
	wire _w16138_ ;
	wire _w16137_ ;
	wire _w16136_ ;
	wire _w16135_ ;
	wire _w16134_ ;
	wire _w16133_ ;
	wire _w16132_ ;
	wire _w16131_ ;
	wire _w16130_ ;
	wire _w16129_ ;
	wire _w16128_ ;
	wire _w16127_ ;
	wire _w16126_ ;
	wire _w16125_ ;
	wire _w16124_ ;
	wire _w16123_ ;
	wire _w16122_ ;
	wire _w16121_ ;
	wire _w16120_ ;
	wire _w16119_ ;
	wire _w16118_ ;
	wire _w16117_ ;
	wire _w16116_ ;
	wire _w16115_ ;
	wire _w16114_ ;
	wire _w16113_ ;
	wire _w16112_ ;
	wire _w16111_ ;
	wire _w16110_ ;
	wire _w16109_ ;
	wire _w16108_ ;
	wire _w16107_ ;
	wire _w16106_ ;
	wire _w16105_ ;
	wire _w16104_ ;
	wire _w16103_ ;
	wire _w16102_ ;
	wire _w16101_ ;
	wire _w16100_ ;
	wire _w16099_ ;
	wire _w16098_ ;
	wire _w16097_ ;
	wire _w16096_ ;
	wire _w16095_ ;
	wire _w16094_ ;
	wire _w16093_ ;
	wire _w16092_ ;
	wire _w16091_ ;
	wire _w16090_ ;
	wire _w16089_ ;
	wire _w16088_ ;
	wire _w16087_ ;
	wire _w16086_ ;
	wire _w16085_ ;
	wire _w16084_ ;
	wire _w16083_ ;
	wire _w16082_ ;
	wire _w16081_ ;
	wire _w16080_ ;
	wire _w16079_ ;
	wire _w16078_ ;
	wire _w16077_ ;
	wire _w16076_ ;
	wire _w16075_ ;
	wire _w16074_ ;
	wire _w16073_ ;
	wire _w16072_ ;
	wire _w16071_ ;
	wire _w16070_ ;
	wire _w16069_ ;
	wire _w16068_ ;
	wire _w16067_ ;
	wire _w16066_ ;
	wire _w16065_ ;
	wire _w16064_ ;
	wire _w16063_ ;
	wire _w16062_ ;
	wire _w16061_ ;
	wire _w16060_ ;
	wire _w16059_ ;
	wire _w16058_ ;
	wire _w16057_ ;
	wire _w16056_ ;
	wire _w16055_ ;
	wire _w16054_ ;
	wire _w16053_ ;
	wire _w16052_ ;
	wire _w16051_ ;
	wire _w16050_ ;
	wire _w16049_ ;
	wire _w16048_ ;
	wire _w16047_ ;
	wire _w16046_ ;
	wire _w16045_ ;
	wire _w16044_ ;
	wire _w16043_ ;
	wire _w16042_ ;
	wire _w16041_ ;
	wire _w16040_ ;
	wire _w16039_ ;
	wire _w16038_ ;
	wire _w16037_ ;
	wire _w16036_ ;
	wire _w16035_ ;
	wire _w16034_ ;
	wire _w16033_ ;
	wire _w16032_ ;
	wire _w16031_ ;
	wire _w16030_ ;
	wire _w16029_ ;
	wire _w16028_ ;
	wire _w16027_ ;
	wire _w16026_ ;
	wire _w16025_ ;
	wire _w16024_ ;
	wire _w16023_ ;
	wire _w16022_ ;
	wire _w16021_ ;
	wire _w16020_ ;
	wire _w16019_ ;
	wire _w16018_ ;
	wire _w16017_ ;
	wire _w16016_ ;
	wire _w16015_ ;
	wire _w16014_ ;
	wire _w16013_ ;
	wire _w16012_ ;
	wire _w16011_ ;
	wire _w16010_ ;
	wire _w16009_ ;
	wire _w16008_ ;
	wire _w16007_ ;
	wire _w16006_ ;
	wire _w16005_ ;
	wire _w16004_ ;
	wire _w16003_ ;
	wire _w16002_ ;
	wire _w16001_ ;
	wire _w16000_ ;
	wire _w15999_ ;
	wire _w15998_ ;
	wire _w15997_ ;
	wire _w15996_ ;
	wire _w15995_ ;
	wire _w15994_ ;
	wire _w15993_ ;
	wire _w15992_ ;
	wire _w15991_ ;
	wire _w15990_ ;
	wire _w15989_ ;
	wire _w15988_ ;
	wire _w15987_ ;
	wire _w15986_ ;
	wire _w15985_ ;
	wire _w15984_ ;
	wire _w15983_ ;
	wire _w15982_ ;
	wire _w15981_ ;
	wire _w15980_ ;
	wire _w15979_ ;
	wire _w15978_ ;
	wire _w15977_ ;
	wire _w15976_ ;
	wire _w15975_ ;
	wire _w15974_ ;
	wire _w15973_ ;
	wire _w15972_ ;
	wire _w15971_ ;
	wire _w15970_ ;
	wire _w15969_ ;
	wire _w15968_ ;
	wire _w15967_ ;
	wire _w15966_ ;
	wire _w15965_ ;
	wire _w15964_ ;
	wire _w15963_ ;
	wire _w15962_ ;
	wire _w15961_ ;
	wire _w15960_ ;
	wire _w15959_ ;
	wire _w15958_ ;
	wire _w15957_ ;
	wire _w15956_ ;
	wire _w15955_ ;
	wire _w15954_ ;
	wire _w15953_ ;
	wire _w15952_ ;
	wire _w15951_ ;
	wire _w15950_ ;
	wire _w15949_ ;
	wire _w15948_ ;
	wire _w15947_ ;
	wire _w15946_ ;
	wire _w15945_ ;
	wire _w15944_ ;
	wire _w15943_ ;
	wire _w15942_ ;
	wire _w15941_ ;
	wire _w15940_ ;
	wire _w15939_ ;
	wire _w15938_ ;
	wire _w15937_ ;
	wire _w15936_ ;
	wire _w15935_ ;
	wire _w15934_ ;
	wire _w15933_ ;
	wire _w15932_ ;
	wire _w15931_ ;
	wire _w15930_ ;
	wire _w15929_ ;
	wire _w15928_ ;
	wire _w15927_ ;
	wire _w15926_ ;
	wire _w15925_ ;
	wire _w15924_ ;
	wire _w15923_ ;
	wire _w15922_ ;
	wire _w15921_ ;
	wire _w15920_ ;
	wire _w15919_ ;
	wire _w15918_ ;
	wire _w15917_ ;
	wire _w15916_ ;
	wire _w15915_ ;
	wire _w15914_ ;
	wire _w15913_ ;
	wire _w15912_ ;
	wire _w15911_ ;
	wire _w15910_ ;
	wire _w15909_ ;
	wire _w15908_ ;
	wire _w15907_ ;
	wire _w15906_ ;
	wire _w15905_ ;
	wire _w15904_ ;
	wire _w15903_ ;
	wire _w15902_ ;
	wire _w15901_ ;
	wire _w15900_ ;
	wire _w15899_ ;
	wire _w15898_ ;
	wire _w15897_ ;
	wire _w15896_ ;
	wire _w15895_ ;
	wire _w15894_ ;
	wire _w15893_ ;
	wire _w15892_ ;
	wire _w15891_ ;
	wire _w15890_ ;
	wire _w15889_ ;
	wire _w15888_ ;
	wire _w15887_ ;
	wire _w15886_ ;
	wire _w15885_ ;
	wire _w15884_ ;
	wire _w15883_ ;
	wire _w15882_ ;
	wire _w15881_ ;
	wire _w15880_ ;
	wire _w15879_ ;
	wire _w15878_ ;
	wire _w15877_ ;
	wire _w15876_ ;
	wire _w15875_ ;
	wire _w15874_ ;
	wire _w15873_ ;
	wire _w15872_ ;
	wire _w15871_ ;
	wire _w15870_ ;
	wire _w15869_ ;
	wire _w15868_ ;
	wire _w15867_ ;
	wire _w15866_ ;
	wire _w15865_ ;
	wire _w15864_ ;
	wire _w15863_ ;
	wire _w15862_ ;
	wire _w15861_ ;
	wire _w15860_ ;
	wire _w15859_ ;
	wire _w15858_ ;
	wire _w15857_ ;
	wire _w15856_ ;
	wire _w15855_ ;
	wire _w15854_ ;
	wire _w15853_ ;
	wire _w15852_ ;
	wire _w15851_ ;
	wire _w15850_ ;
	wire _w15849_ ;
	wire _w15848_ ;
	wire _w15847_ ;
	wire _w15846_ ;
	wire _w15845_ ;
	wire _w15844_ ;
	wire _w15843_ ;
	wire _w15842_ ;
	wire _w15841_ ;
	wire _w15840_ ;
	wire _w15839_ ;
	wire _w15838_ ;
	wire _w15837_ ;
	wire _w15836_ ;
	wire _w15835_ ;
	wire _w15834_ ;
	wire _w15833_ ;
	wire _w15832_ ;
	wire _w15831_ ;
	wire _w15830_ ;
	wire _w15829_ ;
	wire _w15828_ ;
	wire _w15827_ ;
	wire _w15826_ ;
	wire _w15825_ ;
	wire _w15824_ ;
	wire _w15823_ ;
	wire _w15822_ ;
	wire _w15821_ ;
	wire _w15820_ ;
	wire _w15819_ ;
	wire _w15818_ ;
	wire _w15817_ ;
	wire _w15816_ ;
	wire _w15815_ ;
	wire _w15814_ ;
	wire _w15813_ ;
	wire _w15812_ ;
	wire _w15811_ ;
	wire _w15810_ ;
	wire _w15809_ ;
	wire _w15808_ ;
	wire _w15807_ ;
	wire _w15806_ ;
	wire _w15805_ ;
	wire _w15804_ ;
	wire _w15803_ ;
	wire _w15802_ ;
	wire _w15801_ ;
	wire _w15800_ ;
	wire _w15799_ ;
	wire _w15798_ ;
	wire _w15797_ ;
	wire _w15796_ ;
	wire _w15795_ ;
	wire _w15794_ ;
	wire _w15793_ ;
	wire _w15792_ ;
	wire _w15791_ ;
	wire _w15790_ ;
	wire _w15789_ ;
	wire _w15788_ ;
	wire _w15787_ ;
	wire _w15786_ ;
	wire _w15785_ ;
	wire _w15784_ ;
	wire _w15783_ ;
	wire _w15782_ ;
	wire _w15781_ ;
	wire _w15780_ ;
	wire _w15779_ ;
	wire _w15778_ ;
	wire _w15777_ ;
	wire _w15776_ ;
	wire _w15775_ ;
	wire _w15774_ ;
	wire _w15773_ ;
	wire _w15772_ ;
	wire _w15771_ ;
	wire _w15770_ ;
	wire _w15769_ ;
	wire _w15768_ ;
	wire _w15767_ ;
	wire _w15766_ ;
	wire _w15765_ ;
	wire _w15764_ ;
	wire _w15763_ ;
	wire _w15762_ ;
	wire _w15761_ ;
	wire _w15760_ ;
	wire _w15759_ ;
	wire _w15758_ ;
	wire _w15757_ ;
	wire _w15756_ ;
	wire _w15755_ ;
	wire _w15754_ ;
	wire _w15753_ ;
	wire _w15752_ ;
	wire _w15751_ ;
	wire _w15750_ ;
	wire _w15749_ ;
	wire _w15748_ ;
	wire _w15747_ ;
	wire _w15746_ ;
	wire _w15745_ ;
	wire _w15744_ ;
	wire _w15743_ ;
	wire _w15742_ ;
	wire _w15741_ ;
	wire _w15740_ ;
	wire _w15739_ ;
	wire _w15738_ ;
	wire _w15737_ ;
	wire _w15736_ ;
	wire _w15735_ ;
	wire _w15734_ ;
	wire _w15733_ ;
	wire _w15732_ ;
	wire _w15731_ ;
	wire _w15730_ ;
	wire _w15729_ ;
	wire _w15728_ ;
	wire _w15727_ ;
	wire _w15726_ ;
	wire _w15725_ ;
	wire _w15724_ ;
	wire _w15723_ ;
	wire _w15722_ ;
	wire _w15721_ ;
	wire _w15720_ ;
	wire _w15719_ ;
	wire _w15718_ ;
	wire _w15717_ ;
	wire _w15716_ ;
	wire _w15715_ ;
	wire _w15714_ ;
	wire _w15713_ ;
	wire _w15712_ ;
	wire _w15711_ ;
	wire _w15710_ ;
	wire _w15709_ ;
	wire _w15708_ ;
	wire _w15707_ ;
	wire _w15706_ ;
	wire _w15705_ ;
	wire _w15704_ ;
	wire _w15703_ ;
	wire _w15702_ ;
	wire _w15701_ ;
	wire _w15700_ ;
	wire _w15699_ ;
	wire _w15698_ ;
	wire _w15697_ ;
	wire _w15696_ ;
	wire _w15695_ ;
	wire _w15694_ ;
	wire _w15693_ ;
	wire _w15692_ ;
	wire _w15691_ ;
	wire _w15690_ ;
	wire _w15689_ ;
	wire _w15688_ ;
	wire _w15687_ ;
	wire _w15686_ ;
	wire _w15685_ ;
	wire _w15684_ ;
	wire _w15683_ ;
	wire _w15682_ ;
	wire _w15681_ ;
	wire _w15680_ ;
	wire _w15679_ ;
	wire _w15678_ ;
	wire _w15677_ ;
	wire _w15676_ ;
	wire _w15675_ ;
	wire _w15674_ ;
	wire _w15673_ ;
	wire _w15672_ ;
	wire _w15671_ ;
	wire _w15670_ ;
	wire _w15669_ ;
	wire _w15668_ ;
	wire _w15667_ ;
	wire _w15666_ ;
	wire _w15665_ ;
	wire _w15664_ ;
	wire _w15663_ ;
	wire _w15662_ ;
	wire _w15661_ ;
	wire _w15660_ ;
	wire _w15659_ ;
	wire _w15658_ ;
	wire _w15657_ ;
	wire _w15656_ ;
	wire _w15655_ ;
	wire _w15654_ ;
	wire _w15653_ ;
	wire _w15652_ ;
	wire _w15651_ ;
	wire _w15650_ ;
	wire _w15649_ ;
	wire _w15648_ ;
	wire _w15647_ ;
	wire _w15646_ ;
	wire _w15645_ ;
	wire _w15644_ ;
	wire _w15643_ ;
	wire _w15642_ ;
	wire _w15641_ ;
	wire _w15640_ ;
	wire _w15639_ ;
	wire _w15638_ ;
	wire _w15637_ ;
	wire _w15636_ ;
	wire _w15635_ ;
	wire _w15634_ ;
	wire _w15633_ ;
	wire _w15632_ ;
	wire _w15631_ ;
	wire _w15630_ ;
	wire _w15629_ ;
	wire _w15628_ ;
	wire _w15627_ ;
	wire _w15626_ ;
	wire _w15625_ ;
	wire _w15624_ ;
	wire _w15623_ ;
	wire _w15622_ ;
	wire _w15621_ ;
	wire _w15620_ ;
	wire _w15619_ ;
	wire _w15618_ ;
	wire _w15617_ ;
	wire _w15616_ ;
	wire _w15615_ ;
	wire _w15614_ ;
	wire _w15613_ ;
	wire _w15612_ ;
	wire _w15611_ ;
	wire _w15610_ ;
	wire _w15609_ ;
	wire _w15608_ ;
	wire _w15607_ ;
	wire _w15606_ ;
	wire _w15605_ ;
	wire _w15604_ ;
	wire _w15603_ ;
	wire _w15602_ ;
	wire _w15601_ ;
	wire _w15600_ ;
	wire _w15599_ ;
	wire _w15598_ ;
	wire _w15597_ ;
	wire _w15596_ ;
	wire _w15595_ ;
	wire _w15594_ ;
	wire _w15593_ ;
	wire _w15592_ ;
	wire _w15591_ ;
	wire _w15590_ ;
	wire _w15589_ ;
	wire _w15588_ ;
	wire _w15587_ ;
	wire _w15586_ ;
	wire _w15585_ ;
	wire _w15584_ ;
	wire _w15583_ ;
	wire _w15582_ ;
	wire _w15581_ ;
	wire _w15580_ ;
	wire _w15579_ ;
	wire _w15578_ ;
	wire _w15577_ ;
	wire _w15576_ ;
	wire _w15575_ ;
	wire _w15574_ ;
	wire _w15573_ ;
	wire _w15572_ ;
	wire _w15571_ ;
	wire _w15570_ ;
	wire _w15569_ ;
	wire _w15568_ ;
	wire _w15567_ ;
	wire _w15566_ ;
	wire _w15565_ ;
	wire _w15564_ ;
	wire _w15563_ ;
	wire _w15562_ ;
	wire _w15561_ ;
	wire _w15560_ ;
	wire _w15559_ ;
	wire _w15558_ ;
	wire _w15557_ ;
	wire _w15556_ ;
	wire _w15555_ ;
	wire _w15554_ ;
	wire _w15553_ ;
	wire _w15552_ ;
	wire _w15551_ ;
	wire _w15550_ ;
	wire _w15549_ ;
	wire _w15548_ ;
	wire _w15547_ ;
	wire _w15546_ ;
	wire _w15545_ ;
	wire _w15544_ ;
	wire _w15543_ ;
	wire _w15542_ ;
	wire _w15541_ ;
	wire _w15540_ ;
	wire _w15539_ ;
	wire _w15538_ ;
	wire _w15537_ ;
	wire _w15536_ ;
	wire _w15535_ ;
	wire _w15534_ ;
	wire _w15533_ ;
	wire _w15532_ ;
	wire _w15531_ ;
	wire _w15530_ ;
	wire _w15529_ ;
	wire _w15528_ ;
	wire _w15527_ ;
	wire _w15526_ ;
	wire _w15525_ ;
	wire _w15524_ ;
	wire _w15523_ ;
	wire _w15522_ ;
	wire _w15521_ ;
	wire _w15520_ ;
	wire _w15519_ ;
	wire _w15518_ ;
	wire _w15517_ ;
	wire _w15516_ ;
	wire _w15515_ ;
	wire _w15514_ ;
	wire _w15513_ ;
	wire _w15512_ ;
	wire _w15511_ ;
	wire _w15510_ ;
	wire _w15509_ ;
	wire _w15508_ ;
	wire _w15507_ ;
	wire _w15506_ ;
	wire _w15505_ ;
	wire _w15504_ ;
	wire _w15503_ ;
	wire _w15502_ ;
	wire _w15501_ ;
	wire _w15500_ ;
	wire _w15499_ ;
	wire _w15498_ ;
	wire _w15497_ ;
	wire _w15496_ ;
	wire _w15495_ ;
	wire _w15494_ ;
	wire _w15493_ ;
	wire _w15492_ ;
	wire _w15491_ ;
	wire _w15490_ ;
	wire _w15489_ ;
	wire _w15488_ ;
	wire _w15487_ ;
	wire _w15486_ ;
	wire _w15485_ ;
	wire _w15484_ ;
	wire _w15483_ ;
	wire _w15482_ ;
	wire _w15481_ ;
	wire _w15480_ ;
	wire _w15479_ ;
	wire _w15478_ ;
	wire _w15477_ ;
	wire _w15476_ ;
	wire _w15475_ ;
	wire _w15474_ ;
	wire _w15473_ ;
	wire _w15472_ ;
	wire _w15471_ ;
	wire _w15470_ ;
	wire _w15469_ ;
	wire _w15468_ ;
	wire _w15467_ ;
	wire _w15466_ ;
	wire _w15465_ ;
	wire _w15464_ ;
	wire _w15463_ ;
	wire _w15462_ ;
	wire _w15461_ ;
	wire _w15460_ ;
	wire _w15459_ ;
	wire _w15458_ ;
	wire _w15457_ ;
	wire _w15456_ ;
	wire _w15455_ ;
	wire _w15454_ ;
	wire _w15453_ ;
	wire _w15452_ ;
	wire _w15451_ ;
	wire _w15450_ ;
	wire _w15449_ ;
	wire _w15448_ ;
	wire _w15447_ ;
	wire _w15446_ ;
	wire _w15445_ ;
	wire _w15444_ ;
	wire _w15443_ ;
	wire _w15442_ ;
	wire _w15441_ ;
	wire _w15440_ ;
	wire _w15439_ ;
	wire _w15438_ ;
	wire _w15437_ ;
	wire _w15436_ ;
	wire _w15435_ ;
	wire _w15434_ ;
	wire _w15433_ ;
	wire _w15432_ ;
	wire _w15431_ ;
	wire _w15430_ ;
	wire _w15429_ ;
	wire _w15428_ ;
	wire _w15427_ ;
	wire _w15426_ ;
	wire _w15425_ ;
	wire _w15424_ ;
	wire _w15423_ ;
	wire _w15422_ ;
	wire _w15421_ ;
	wire _w15420_ ;
	wire _w15419_ ;
	wire _w15418_ ;
	wire _w15417_ ;
	wire _w15416_ ;
	wire _w15415_ ;
	wire _w15414_ ;
	wire _w15413_ ;
	wire _w15412_ ;
	wire _w15411_ ;
	wire _w15410_ ;
	wire _w15409_ ;
	wire _w15408_ ;
	wire _w15407_ ;
	wire _w15406_ ;
	wire _w15405_ ;
	wire _w15404_ ;
	wire _w15403_ ;
	wire _w15402_ ;
	wire _w15401_ ;
	wire _w15400_ ;
	wire _w15399_ ;
	wire _w15398_ ;
	wire _w15397_ ;
	wire _w15396_ ;
	wire _w15395_ ;
	wire _w15394_ ;
	wire _w15393_ ;
	wire _w15392_ ;
	wire _w15391_ ;
	wire _w15390_ ;
	wire _w15389_ ;
	wire _w15388_ ;
	wire _w15387_ ;
	wire _w15386_ ;
	wire _w15385_ ;
	wire _w15384_ ;
	wire _w15383_ ;
	wire _w15382_ ;
	wire _w15381_ ;
	wire _w15380_ ;
	wire _w15379_ ;
	wire _w15378_ ;
	wire _w15377_ ;
	wire _w15376_ ;
	wire _w15375_ ;
	wire _w15374_ ;
	wire _w15373_ ;
	wire _w15372_ ;
	wire _w15371_ ;
	wire _w15370_ ;
	wire _w15369_ ;
	wire _w15368_ ;
	wire _w15367_ ;
	wire _w15366_ ;
	wire _w15365_ ;
	wire _w15364_ ;
	wire _w15363_ ;
	wire _w15362_ ;
	wire _w15361_ ;
	wire _w15360_ ;
	wire _w15359_ ;
	wire _w15358_ ;
	wire _w15357_ ;
	wire _w15356_ ;
	wire _w15355_ ;
	wire _w15354_ ;
	wire _w15353_ ;
	wire _w15352_ ;
	wire _w15351_ ;
	wire _w15350_ ;
	wire _w15349_ ;
	wire _w15348_ ;
	wire _w15347_ ;
	wire _w15346_ ;
	wire _w15345_ ;
	wire _w15344_ ;
	wire _w15343_ ;
	wire _w15342_ ;
	wire _w15341_ ;
	wire _w15340_ ;
	wire _w15339_ ;
	wire _w15338_ ;
	wire _w15337_ ;
	wire _w15336_ ;
	wire _w15335_ ;
	wire _w15334_ ;
	wire _w15333_ ;
	wire _w15332_ ;
	wire _w15331_ ;
	wire _w15330_ ;
	wire _w15329_ ;
	wire _w15328_ ;
	wire _w15327_ ;
	wire _w15326_ ;
	wire _w15325_ ;
	wire _w15324_ ;
	wire _w15323_ ;
	wire _w15322_ ;
	wire _w15321_ ;
	wire _w15320_ ;
	wire _w15319_ ;
	wire _w15318_ ;
	wire _w15317_ ;
	wire _w15316_ ;
	wire _w15315_ ;
	wire _w15314_ ;
	wire _w15313_ ;
	wire _w15312_ ;
	wire _w15311_ ;
	wire _w15310_ ;
	wire _w15309_ ;
	wire _w15308_ ;
	wire _w15307_ ;
	wire _w15306_ ;
	wire _w15305_ ;
	wire _w15304_ ;
	wire _w15303_ ;
	wire _w15302_ ;
	wire _w15301_ ;
	wire _w15300_ ;
	wire _w15299_ ;
	wire _w15298_ ;
	wire _w15297_ ;
	wire _w15296_ ;
	wire _w15295_ ;
	wire _w15294_ ;
	wire _w15293_ ;
	wire _w15292_ ;
	wire _w15291_ ;
	wire _w15290_ ;
	wire _w15289_ ;
	wire _w15288_ ;
	wire _w15287_ ;
	wire _w15286_ ;
	wire _w15285_ ;
	wire _w15284_ ;
	wire _w15283_ ;
	wire _w15282_ ;
	wire _w15281_ ;
	wire _w15280_ ;
	wire _w15279_ ;
	wire _w15278_ ;
	wire _w15277_ ;
	wire _w15276_ ;
	wire _w15275_ ;
	wire _w15274_ ;
	wire _w15273_ ;
	wire _w15272_ ;
	wire _w15271_ ;
	wire _w15270_ ;
	wire _w15269_ ;
	wire _w15268_ ;
	wire _w15267_ ;
	wire _w15266_ ;
	wire _w15265_ ;
	wire _w15264_ ;
	wire _w15263_ ;
	wire _w15262_ ;
	wire _w15261_ ;
	wire _w15260_ ;
	wire _w15259_ ;
	wire _w15258_ ;
	wire _w15257_ ;
	wire _w15256_ ;
	wire _w15255_ ;
	wire _w15254_ ;
	wire _w15253_ ;
	wire _w15252_ ;
	wire _w15251_ ;
	wire _w15250_ ;
	wire _w15249_ ;
	wire _w15248_ ;
	wire _w15247_ ;
	wire _w15246_ ;
	wire _w15245_ ;
	wire _w15244_ ;
	wire _w15243_ ;
	wire _w15242_ ;
	wire _w15241_ ;
	wire _w15240_ ;
	wire _w15239_ ;
	wire _w15238_ ;
	wire _w15237_ ;
	wire _w15236_ ;
	wire _w15235_ ;
	wire _w15234_ ;
	wire _w15233_ ;
	wire _w15232_ ;
	wire _w15231_ ;
	wire _w15230_ ;
	wire _w15229_ ;
	wire _w15228_ ;
	wire _w15227_ ;
	wire _w15226_ ;
	wire _w15225_ ;
	wire _w15224_ ;
	wire _w15223_ ;
	wire _w15222_ ;
	wire _w15221_ ;
	wire _w15220_ ;
	wire _w15219_ ;
	wire _w15218_ ;
	wire _w15217_ ;
	wire _w15216_ ;
	wire _w15215_ ;
	wire _w15214_ ;
	wire _w15213_ ;
	wire _w15212_ ;
	wire _w15211_ ;
	wire _w15210_ ;
	wire _w15209_ ;
	wire _w15208_ ;
	wire _w15207_ ;
	wire _w15206_ ;
	wire _w15205_ ;
	wire _w15204_ ;
	wire _w15203_ ;
	wire _w15202_ ;
	wire _w15201_ ;
	wire _w15200_ ;
	wire _w15199_ ;
	wire _w15198_ ;
	wire _w15197_ ;
	wire _w15196_ ;
	wire _w15195_ ;
	wire _w15194_ ;
	wire _w15193_ ;
	wire _w15192_ ;
	wire _w15191_ ;
	wire _w15190_ ;
	wire _w15189_ ;
	wire _w15188_ ;
	wire _w15187_ ;
	wire _w15186_ ;
	wire _w15185_ ;
	wire _w15184_ ;
	wire _w15183_ ;
	wire _w15182_ ;
	wire _w15181_ ;
	wire _w15180_ ;
	wire _w15179_ ;
	wire _w15178_ ;
	wire _w15177_ ;
	wire _w15176_ ;
	wire _w15175_ ;
	wire _w15174_ ;
	wire _w15173_ ;
	wire _w15172_ ;
	wire _w15171_ ;
	wire _w15170_ ;
	wire _w15169_ ;
	wire _w15168_ ;
	wire _w15167_ ;
	wire _w15166_ ;
	wire _w15165_ ;
	wire _w15164_ ;
	wire _w15163_ ;
	wire _w15162_ ;
	wire _w15161_ ;
	wire _w15160_ ;
	wire _w15159_ ;
	wire _w15158_ ;
	wire _w15157_ ;
	wire _w15156_ ;
	wire _w15155_ ;
	wire _w15154_ ;
	wire _w15153_ ;
	wire _w15152_ ;
	wire _w15151_ ;
	wire _w15150_ ;
	wire _w15149_ ;
	wire _w15148_ ;
	wire _w15147_ ;
	wire _w15146_ ;
	wire _w15145_ ;
	wire _w15144_ ;
	wire _w15143_ ;
	wire _w15142_ ;
	wire _w15141_ ;
	wire _w15140_ ;
	wire _w15139_ ;
	wire _w15138_ ;
	wire _w15137_ ;
	wire _w15136_ ;
	wire _w15135_ ;
	wire _w15134_ ;
	wire _w15133_ ;
	wire _w15132_ ;
	wire _w15131_ ;
	wire _w15130_ ;
	wire _w15129_ ;
	wire _w15128_ ;
	wire _w15127_ ;
	wire _w15126_ ;
	wire _w15125_ ;
	wire _w15124_ ;
	wire _w15123_ ;
	wire _w15122_ ;
	wire _w15121_ ;
	wire _w15120_ ;
	wire _w15119_ ;
	wire _w15118_ ;
	wire _w15117_ ;
	wire _w15116_ ;
	wire _w15115_ ;
	wire _w15114_ ;
	wire _w15113_ ;
	wire _w15112_ ;
	wire _w15111_ ;
	wire _w15110_ ;
	wire _w15109_ ;
	wire _w15108_ ;
	wire _w15107_ ;
	wire _w15106_ ;
	wire _w15105_ ;
	wire _w15104_ ;
	wire _w15103_ ;
	wire _w15102_ ;
	wire _w15101_ ;
	wire _w15100_ ;
	wire _w15099_ ;
	wire _w15098_ ;
	wire _w15097_ ;
	wire _w15096_ ;
	wire _w15095_ ;
	wire _w15094_ ;
	wire _w15093_ ;
	wire _w15092_ ;
	wire _w15091_ ;
	wire _w15090_ ;
	wire _w15089_ ;
	wire _w15088_ ;
	wire _w15087_ ;
	wire _w15086_ ;
	wire _w15085_ ;
	wire _w15084_ ;
	wire _w15083_ ;
	wire _w15082_ ;
	wire _w15081_ ;
	wire _w15080_ ;
	wire _w15079_ ;
	wire _w15078_ ;
	wire _w15077_ ;
	wire _w15076_ ;
	wire _w15075_ ;
	wire _w15074_ ;
	wire _w15073_ ;
	wire _w15072_ ;
	wire _w15071_ ;
	wire _w15070_ ;
	wire _w15069_ ;
	wire _w15068_ ;
	wire _w15067_ ;
	wire _w15066_ ;
	wire _w15065_ ;
	wire _w15064_ ;
	wire _w15063_ ;
	wire _w15062_ ;
	wire _w15061_ ;
	wire _w15060_ ;
	wire _w15059_ ;
	wire _w15058_ ;
	wire _w15057_ ;
	wire _w15056_ ;
	wire _w15055_ ;
	wire _w15054_ ;
	wire _w15053_ ;
	wire _w15052_ ;
	wire _w15051_ ;
	wire _w15050_ ;
	wire _w15049_ ;
	wire _w15048_ ;
	wire _w15047_ ;
	wire _w15046_ ;
	wire _w15045_ ;
	wire _w15044_ ;
	wire _w15043_ ;
	wire _w15042_ ;
	wire _w15041_ ;
	wire _w15040_ ;
	wire _w15039_ ;
	wire _w15038_ ;
	wire _w15037_ ;
	wire _w15036_ ;
	wire _w15035_ ;
	wire _w15034_ ;
	wire _w15033_ ;
	wire _w15032_ ;
	wire _w15031_ ;
	wire _w15030_ ;
	wire _w15029_ ;
	wire _w15028_ ;
	wire _w15027_ ;
	wire _w15026_ ;
	wire _w15025_ ;
	wire _w15024_ ;
	wire _w15023_ ;
	wire _w15022_ ;
	wire _w15021_ ;
	wire _w15020_ ;
	wire _w15019_ ;
	wire _w15018_ ;
	wire _w15017_ ;
	wire _w15016_ ;
	wire _w15015_ ;
	wire _w15014_ ;
	wire _w15013_ ;
	wire _w15012_ ;
	wire _w15011_ ;
	wire _w15010_ ;
	wire _w15009_ ;
	wire _w15008_ ;
	wire _w15007_ ;
	wire _w15006_ ;
	wire _w15005_ ;
	wire _w15004_ ;
	wire _w15003_ ;
	wire _w15002_ ;
	wire _w15001_ ;
	wire _w15000_ ;
	wire _w14999_ ;
	wire _w14998_ ;
	wire _w14997_ ;
	wire _w14996_ ;
	wire _w14995_ ;
	wire _w14994_ ;
	wire _w14993_ ;
	wire _w14992_ ;
	wire _w14991_ ;
	wire _w14990_ ;
	wire _w14989_ ;
	wire _w14988_ ;
	wire _w14987_ ;
	wire _w14986_ ;
	wire _w14985_ ;
	wire _w14984_ ;
	wire _w14983_ ;
	wire _w14982_ ;
	wire _w14981_ ;
	wire _w14980_ ;
	wire _w14979_ ;
	wire _w14978_ ;
	wire _w14977_ ;
	wire _w14976_ ;
	wire _w14975_ ;
	wire _w14974_ ;
	wire _w14973_ ;
	wire _w14972_ ;
	wire _w14971_ ;
	wire _w14970_ ;
	wire _w14969_ ;
	wire _w14968_ ;
	wire _w14967_ ;
	wire _w14966_ ;
	wire _w14965_ ;
	wire _w14964_ ;
	wire _w14963_ ;
	wire _w14962_ ;
	wire _w14961_ ;
	wire _w14960_ ;
	wire _w14959_ ;
	wire _w14958_ ;
	wire _w14957_ ;
	wire _w14956_ ;
	wire _w14955_ ;
	wire _w14954_ ;
	wire _w14953_ ;
	wire _w14952_ ;
	wire _w14951_ ;
	wire _w14950_ ;
	wire _w14949_ ;
	wire _w14948_ ;
	wire _w14947_ ;
	wire _w14946_ ;
	wire _w14945_ ;
	wire _w14944_ ;
	wire _w14943_ ;
	wire _w14942_ ;
	wire _w14941_ ;
	wire _w14940_ ;
	wire _w14939_ ;
	wire _w14938_ ;
	wire _w14937_ ;
	wire _w14936_ ;
	wire _w14935_ ;
	wire _w14934_ ;
	wire _w14933_ ;
	wire _w14932_ ;
	wire _w14931_ ;
	wire _w14930_ ;
	wire _w14929_ ;
	wire _w14928_ ;
	wire _w14927_ ;
	wire _w14926_ ;
	wire _w14925_ ;
	wire _w14924_ ;
	wire _w14923_ ;
	wire _w14922_ ;
	wire _w14921_ ;
	wire _w14920_ ;
	wire _w14919_ ;
	wire _w14918_ ;
	wire _w14917_ ;
	wire _w14916_ ;
	wire _w14915_ ;
	wire _w14914_ ;
	wire _w14913_ ;
	wire _w14912_ ;
	wire _w14911_ ;
	wire _w14910_ ;
	wire _w14909_ ;
	wire _w14908_ ;
	wire _w14907_ ;
	wire _w14906_ ;
	wire _w14905_ ;
	wire _w14904_ ;
	wire _w14903_ ;
	wire _w14902_ ;
	wire _w14901_ ;
	wire _w14900_ ;
	wire _w14899_ ;
	wire _w14898_ ;
	wire _w14897_ ;
	wire _w14896_ ;
	wire _w14895_ ;
	wire _w14894_ ;
	wire _w14893_ ;
	wire _w14892_ ;
	wire _w14891_ ;
	wire _w14890_ ;
	wire _w14889_ ;
	wire _w14888_ ;
	wire _w14887_ ;
	wire _w14886_ ;
	wire _w14885_ ;
	wire _w14884_ ;
	wire _w14883_ ;
	wire _w14882_ ;
	wire _w14881_ ;
	wire _w14880_ ;
	wire _w14879_ ;
	wire _w14878_ ;
	wire _w14877_ ;
	wire _w14876_ ;
	wire _w14875_ ;
	wire _w14874_ ;
	wire _w14873_ ;
	wire _w14872_ ;
	wire _w14871_ ;
	wire _w14870_ ;
	wire _w14869_ ;
	wire _w14868_ ;
	wire _w14867_ ;
	wire _w14866_ ;
	wire _w14865_ ;
	wire _w14864_ ;
	wire _w14863_ ;
	wire _w14862_ ;
	wire _w14861_ ;
	wire _w14860_ ;
	wire _w14859_ ;
	wire _w14858_ ;
	wire _w14857_ ;
	wire _w14856_ ;
	wire _w14855_ ;
	wire _w14854_ ;
	wire _w14853_ ;
	wire _w14852_ ;
	wire _w14851_ ;
	wire _w14850_ ;
	wire _w14849_ ;
	wire _w14848_ ;
	wire _w14847_ ;
	wire _w14846_ ;
	wire _w14845_ ;
	wire _w14844_ ;
	wire _w14843_ ;
	wire _w14842_ ;
	wire _w14841_ ;
	wire _w14840_ ;
	wire _w14839_ ;
	wire _w14838_ ;
	wire _w14837_ ;
	wire _w14836_ ;
	wire _w14835_ ;
	wire _w14834_ ;
	wire _w14833_ ;
	wire _w14832_ ;
	wire _w14831_ ;
	wire _w14830_ ;
	wire _w14829_ ;
	wire _w14828_ ;
	wire _w14827_ ;
	wire _w14826_ ;
	wire _w14825_ ;
	wire _w14824_ ;
	wire _w14823_ ;
	wire _w14822_ ;
	wire _w14821_ ;
	wire _w14820_ ;
	wire _w14819_ ;
	wire _w14818_ ;
	wire _w14817_ ;
	wire _w14816_ ;
	wire _w14815_ ;
	wire _w14814_ ;
	wire _w14813_ ;
	wire _w14812_ ;
	wire _w14811_ ;
	wire _w14810_ ;
	wire _w14809_ ;
	wire _w14808_ ;
	wire _w14807_ ;
	wire _w14806_ ;
	wire _w14805_ ;
	wire _w14804_ ;
	wire _w14803_ ;
	wire _w14802_ ;
	wire _w14801_ ;
	wire _w14800_ ;
	wire _w14799_ ;
	wire _w14798_ ;
	wire _w14797_ ;
	wire _w14796_ ;
	wire _w14795_ ;
	wire _w14794_ ;
	wire _w14793_ ;
	wire _w14792_ ;
	wire _w14791_ ;
	wire _w14790_ ;
	wire _w14789_ ;
	wire _w14788_ ;
	wire _w14787_ ;
	wire _w14786_ ;
	wire _w14785_ ;
	wire _w14784_ ;
	wire _w14783_ ;
	wire _w14782_ ;
	wire _w14781_ ;
	wire _w14780_ ;
	wire _w14779_ ;
	wire _w14778_ ;
	wire _w14777_ ;
	wire _w14776_ ;
	wire _w14775_ ;
	wire _w14774_ ;
	wire _w14773_ ;
	wire _w14772_ ;
	wire _w14771_ ;
	wire _w14770_ ;
	wire _w14769_ ;
	wire _w14768_ ;
	wire _w14767_ ;
	wire _w14766_ ;
	wire _w14765_ ;
	wire _w14764_ ;
	wire _w14763_ ;
	wire _w14762_ ;
	wire _w14761_ ;
	wire _w14760_ ;
	wire _w14759_ ;
	wire _w14758_ ;
	wire _w14757_ ;
	wire _w14756_ ;
	wire _w14755_ ;
	wire _w14754_ ;
	wire _w14753_ ;
	wire _w14752_ ;
	wire _w14751_ ;
	wire _w14750_ ;
	wire _w14749_ ;
	wire _w14748_ ;
	wire _w14747_ ;
	wire _w14746_ ;
	wire _w14745_ ;
	wire _w14744_ ;
	wire _w14743_ ;
	wire _w14742_ ;
	wire _w14741_ ;
	wire _w14740_ ;
	wire _w14739_ ;
	wire _w14738_ ;
	wire _w14737_ ;
	wire _w14736_ ;
	wire _w14735_ ;
	wire _w14734_ ;
	wire _w14733_ ;
	wire _w14732_ ;
	wire _w14731_ ;
	wire _w14730_ ;
	wire _w14729_ ;
	wire _w14728_ ;
	wire _w14727_ ;
	wire _w14726_ ;
	wire _w14725_ ;
	wire _w14724_ ;
	wire _w14723_ ;
	wire _w14722_ ;
	wire _w14721_ ;
	wire _w14720_ ;
	wire _w14719_ ;
	wire _w14718_ ;
	wire _w14717_ ;
	wire _w14716_ ;
	wire _w14715_ ;
	wire _w14714_ ;
	wire _w14713_ ;
	wire _w14712_ ;
	wire _w14711_ ;
	wire _w14710_ ;
	wire _w14709_ ;
	wire _w14708_ ;
	wire _w14707_ ;
	wire _w14706_ ;
	wire _w14705_ ;
	wire _w14704_ ;
	wire _w14703_ ;
	wire _w14702_ ;
	wire _w14701_ ;
	wire _w14700_ ;
	wire _w14699_ ;
	wire _w14698_ ;
	wire _w14697_ ;
	wire _w14696_ ;
	wire _w14695_ ;
	wire _w14694_ ;
	wire _w14693_ ;
	wire _w14692_ ;
	wire _w14691_ ;
	wire _w14690_ ;
	wire _w14689_ ;
	wire _w14688_ ;
	wire _w14687_ ;
	wire _w14686_ ;
	wire _w14685_ ;
	wire _w14684_ ;
	wire _w14683_ ;
	wire _w14682_ ;
	wire _w14681_ ;
	wire _w14680_ ;
	wire _w14679_ ;
	wire _w14678_ ;
	wire _w14677_ ;
	wire _w14676_ ;
	wire _w14675_ ;
	wire _w14674_ ;
	wire _w14673_ ;
	wire _w14672_ ;
	wire _w14671_ ;
	wire _w14670_ ;
	wire _w14669_ ;
	wire _w14668_ ;
	wire _w14667_ ;
	wire _w14666_ ;
	wire _w14665_ ;
	wire _w14664_ ;
	wire _w14663_ ;
	wire _w14662_ ;
	wire _w14661_ ;
	wire _w14660_ ;
	wire _w14659_ ;
	wire _w14658_ ;
	wire _w14657_ ;
	wire _w14656_ ;
	wire _w14655_ ;
	wire _w14654_ ;
	wire _w14653_ ;
	wire _w14652_ ;
	wire _w14651_ ;
	wire _w14650_ ;
	wire _w14649_ ;
	wire _w14648_ ;
	wire _w14647_ ;
	wire _w14646_ ;
	wire _w14645_ ;
	wire _w14644_ ;
	wire _w14643_ ;
	wire _w14642_ ;
	wire _w14641_ ;
	wire _w14640_ ;
	wire _w14639_ ;
	wire _w14638_ ;
	wire _w14637_ ;
	wire _w14636_ ;
	wire _w14635_ ;
	wire _w14634_ ;
	wire _w14633_ ;
	wire _w14632_ ;
	wire _w14631_ ;
	wire _w14630_ ;
	wire _w14629_ ;
	wire _w14628_ ;
	wire _w14627_ ;
	wire _w14626_ ;
	wire _w14625_ ;
	wire _w14624_ ;
	wire _w14623_ ;
	wire _w14622_ ;
	wire _w14621_ ;
	wire _w14620_ ;
	wire _w14619_ ;
	wire _w14618_ ;
	wire _w14617_ ;
	wire _w14616_ ;
	wire _w14615_ ;
	wire _w14614_ ;
	wire _w14613_ ;
	wire _w14612_ ;
	wire _w14611_ ;
	wire _w14610_ ;
	wire _w14609_ ;
	wire _w14608_ ;
	wire _w14607_ ;
	wire _w14606_ ;
	wire _w14605_ ;
	wire _w14604_ ;
	wire _w14603_ ;
	wire _w14602_ ;
	wire _w14601_ ;
	wire _w14600_ ;
	wire _w14599_ ;
	wire _w14598_ ;
	wire _w14597_ ;
	wire _w14596_ ;
	wire _w14595_ ;
	wire _w14594_ ;
	wire _w14593_ ;
	wire _w14592_ ;
	wire _w14591_ ;
	wire _w14590_ ;
	wire _w14589_ ;
	wire _w14588_ ;
	wire _w14587_ ;
	wire _w14586_ ;
	wire _w14585_ ;
	wire _w14584_ ;
	wire _w14583_ ;
	wire _w14582_ ;
	wire _w14581_ ;
	wire _w14580_ ;
	wire _w14579_ ;
	wire _w14578_ ;
	wire _w14577_ ;
	wire _w14576_ ;
	wire _w14575_ ;
	wire _w14574_ ;
	wire _w14573_ ;
	wire _w14572_ ;
	wire _w14571_ ;
	wire _w14570_ ;
	wire _w14569_ ;
	wire _w14568_ ;
	wire _w14567_ ;
	wire _w14566_ ;
	wire _w14565_ ;
	wire _w14564_ ;
	wire _w14563_ ;
	wire _w14562_ ;
	wire _w14561_ ;
	wire _w14560_ ;
	wire _w14559_ ;
	wire _w14558_ ;
	wire _w14557_ ;
	wire _w14556_ ;
	wire _w14555_ ;
	wire _w14554_ ;
	wire _w14553_ ;
	wire _w14552_ ;
	wire _w14551_ ;
	wire _w14550_ ;
	wire _w14549_ ;
	wire _w14548_ ;
	wire _w14547_ ;
	wire _w14546_ ;
	wire _w14545_ ;
	wire _w14544_ ;
	wire _w14543_ ;
	wire _w14542_ ;
	wire _w14541_ ;
	wire _w14540_ ;
	wire _w14539_ ;
	wire _w14538_ ;
	wire _w14537_ ;
	wire _w14536_ ;
	wire _w14535_ ;
	wire _w14534_ ;
	wire _w14533_ ;
	wire _w14532_ ;
	wire _w14531_ ;
	wire _w14530_ ;
	wire _w14529_ ;
	wire _w14528_ ;
	wire _w14527_ ;
	wire _w14526_ ;
	wire _w14525_ ;
	wire _w14524_ ;
	wire _w14523_ ;
	wire _w14522_ ;
	wire _w14521_ ;
	wire _w14520_ ;
	wire _w14519_ ;
	wire _w14518_ ;
	wire _w14517_ ;
	wire _w14516_ ;
	wire _w14515_ ;
	wire _w14514_ ;
	wire _w14513_ ;
	wire _w14512_ ;
	wire _w14511_ ;
	wire _w14510_ ;
	wire _w14509_ ;
	wire _w14508_ ;
	wire _w14507_ ;
	wire _w14506_ ;
	wire _w14505_ ;
	wire _w14504_ ;
	wire _w14503_ ;
	wire _w14502_ ;
	wire _w14501_ ;
	wire _w14500_ ;
	wire _w14499_ ;
	wire _w14498_ ;
	wire _w14497_ ;
	wire _w14496_ ;
	wire _w14495_ ;
	wire _w14494_ ;
	wire _w14493_ ;
	wire _w14492_ ;
	wire _w14491_ ;
	wire _w14490_ ;
	wire _w14489_ ;
	wire _w14488_ ;
	wire _w14487_ ;
	wire _w14486_ ;
	wire _w14485_ ;
	wire _w14484_ ;
	wire _w14483_ ;
	wire _w14482_ ;
	wire _w14481_ ;
	wire _w14480_ ;
	wire _w14479_ ;
	wire _w14478_ ;
	wire _w14477_ ;
	wire _w14476_ ;
	wire _w14475_ ;
	wire _w14474_ ;
	wire _w14473_ ;
	wire _w14472_ ;
	wire _w14471_ ;
	wire _w14470_ ;
	wire _w14469_ ;
	wire _w14468_ ;
	wire _w14467_ ;
	wire _w14466_ ;
	wire _w14465_ ;
	wire _w14464_ ;
	wire _w14463_ ;
	wire _w14462_ ;
	wire _w14461_ ;
	wire _w14460_ ;
	wire _w14459_ ;
	wire _w14458_ ;
	wire _w14457_ ;
	wire _w14456_ ;
	wire _w14455_ ;
	wire _w14454_ ;
	wire _w14453_ ;
	wire _w14452_ ;
	wire _w14451_ ;
	wire _w14450_ ;
	wire _w14449_ ;
	wire _w14448_ ;
	wire _w14447_ ;
	wire _w14446_ ;
	wire _w14445_ ;
	wire _w14444_ ;
	wire _w14443_ ;
	wire _w14442_ ;
	wire _w14441_ ;
	wire _w14440_ ;
	wire _w14439_ ;
	wire _w14438_ ;
	wire _w14437_ ;
	wire _w14436_ ;
	wire _w14435_ ;
	wire _w14434_ ;
	wire _w14433_ ;
	wire _w14432_ ;
	wire _w14431_ ;
	wire _w14430_ ;
	wire _w14429_ ;
	wire _w14428_ ;
	wire _w14427_ ;
	wire _w14426_ ;
	wire _w14425_ ;
	wire _w14424_ ;
	wire _w14423_ ;
	wire _w14422_ ;
	wire _w14421_ ;
	wire _w14420_ ;
	wire _w14419_ ;
	wire _w14418_ ;
	wire _w14417_ ;
	wire _w14416_ ;
	wire _w14415_ ;
	wire _w14414_ ;
	wire _w14413_ ;
	wire _w14412_ ;
	wire _w14411_ ;
	wire _w14410_ ;
	wire _w14409_ ;
	wire _w14408_ ;
	wire _w14407_ ;
	wire _w14406_ ;
	wire _w14405_ ;
	wire _w14404_ ;
	wire _w14403_ ;
	wire _w14402_ ;
	wire _w14401_ ;
	wire _w14400_ ;
	wire _w14399_ ;
	wire _w14398_ ;
	wire _w14397_ ;
	wire _w14396_ ;
	wire _w14395_ ;
	wire _w14394_ ;
	wire _w14393_ ;
	wire _w14392_ ;
	wire _w14391_ ;
	wire _w14390_ ;
	wire _w14389_ ;
	wire _w14388_ ;
	wire _w14387_ ;
	wire _w14386_ ;
	wire _w14385_ ;
	wire _w14384_ ;
	wire _w14383_ ;
	wire _w14382_ ;
	wire _w14381_ ;
	wire _w14380_ ;
	wire _w14379_ ;
	wire _w14378_ ;
	wire _w14377_ ;
	wire _w14376_ ;
	wire _w14375_ ;
	wire _w14374_ ;
	wire _w14373_ ;
	wire _w14372_ ;
	wire _w14371_ ;
	wire _w14370_ ;
	wire _w14369_ ;
	wire _w14368_ ;
	wire _w14367_ ;
	wire _w14366_ ;
	wire _w14365_ ;
	wire _w14364_ ;
	wire _w14363_ ;
	wire _w14362_ ;
	wire _w14361_ ;
	wire _w14360_ ;
	wire _w14359_ ;
	wire _w14358_ ;
	wire _w14357_ ;
	wire _w14356_ ;
	wire _w14355_ ;
	wire _w14354_ ;
	wire _w14353_ ;
	wire _w14352_ ;
	wire _w14351_ ;
	wire _w14350_ ;
	wire _w14349_ ;
	wire _w14348_ ;
	wire _w14347_ ;
	wire _w14346_ ;
	wire _w14345_ ;
	wire _w14344_ ;
	wire _w14343_ ;
	wire _w14342_ ;
	wire _w14341_ ;
	wire _w14340_ ;
	wire _w14339_ ;
	wire _w14338_ ;
	wire _w14337_ ;
	wire _w14336_ ;
	wire _w14335_ ;
	wire _w14334_ ;
	wire _w14333_ ;
	wire _w14332_ ;
	wire _w14331_ ;
	wire _w14330_ ;
	wire _w14329_ ;
	wire _w14328_ ;
	wire _w14327_ ;
	wire _w14326_ ;
	wire _w14325_ ;
	wire _w14324_ ;
	wire _w14323_ ;
	wire _w14322_ ;
	wire _w14321_ ;
	wire _w14320_ ;
	wire _w14319_ ;
	wire _w14318_ ;
	wire _w14317_ ;
	wire _w14316_ ;
	wire _w14315_ ;
	wire _w14314_ ;
	wire _w14313_ ;
	wire _w14312_ ;
	wire _w14311_ ;
	wire _w14310_ ;
	wire _w14309_ ;
	wire _w14308_ ;
	wire _w14307_ ;
	wire _w14306_ ;
	wire _w14305_ ;
	wire _w14304_ ;
	wire _w14303_ ;
	wire _w14302_ ;
	wire _w14301_ ;
	wire _w14300_ ;
	wire _w14299_ ;
	wire _w14298_ ;
	wire _w14297_ ;
	wire _w14296_ ;
	wire _w14295_ ;
	wire _w14294_ ;
	wire _w14293_ ;
	wire _w14292_ ;
	wire _w14291_ ;
	wire _w14290_ ;
	wire _w14289_ ;
	wire _w14288_ ;
	wire _w14287_ ;
	wire _w14286_ ;
	wire _w14285_ ;
	wire _w14284_ ;
	wire _w14283_ ;
	wire _w14282_ ;
	wire _w14281_ ;
	wire _w14280_ ;
	wire _w14279_ ;
	wire _w14278_ ;
	wire _w14277_ ;
	wire _w14276_ ;
	wire _w14275_ ;
	wire _w14274_ ;
	wire _w14273_ ;
	wire _w14272_ ;
	wire _w14271_ ;
	wire _w14270_ ;
	wire _w14269_ ;
	wire _w14268_ ;
	wire _w14267_ ;
	wire _w14266_ ;
	wire _w14265_ ;
	wire _w14264_ ;
	wire _w14263_ ;
	wire _w14262_ ;
	wire _w14261_ ;
	wire _w14260_ ;
	wire _w14259_ ;
	wire _w14258_ ;
	wire _w14257_ ;
	wire _w14256_ ;
	wire _w14255_ ;
	wire _w14254_ ;
	wire _w14253_ ;
	wire _w14252_ ;
	wire _w14251_ ;
	wire _w14250_ ;
	wire _w14249_ ;
	wire _w14248_ ;
	wire _w14247_ ;
	wire _w14246_ ;
	wire _w14245_ ;
	wire _w14244_ ;
	wire _w14243_ ;
	wire _w14242_ ;
	wire _w14241_ ;
	wire _w14240_ ;
	wire _w14239_ ;
	wire _w14238_ ;
	wire _w14237_ ;
	wire _w14236_ ;
	wire _w14235_ ;
	wire _w14234_ ;
	wire _w14233_ ;
	wire _w14232_ ;
	wire _w14231_ ;
	wire _w14230_ ;
	wire _w14229_ ;
	wire _w14228_ ;
	wire _w14227_ ;
	wire _w14226_ ;
	wire _w14225_ ;
	wire _w14224_ ;
	wire _w14223_ ;
	wire _w14222_ ;
	wire _w14221_ ;
	wire _w14220_ ;
	wire _w14219_ ;
	wire _w14218_ ;
	wire _w14217_ ;
	wire _w14216_ ;
	wire _w14215_ ;
	wire _w14214_ ;
	wire _w14213_ ;
	wire _w14212_ ;
	wire _w14211_ ;
	wire _w14210_ ;
	wire _w14209_ ;
	wire _w14208_ ;
	wire _w14207_ ;
	wire _w14206_ ;
	wire _w14205_ ;
	wire _w14204_ ;
	wire _w14203_ ;
	wire _w14202_ ;
	wire _w14201_ ;
	wire _w14200_ ;
	wire _w14199_ ;
	wire _w14198_ ;
	wire _w14197_ ;
	wire _w14196_ ;
	wire _w14195_ ;
	wire _w14194_ ;
	wire _w14193_ ;
	wire _w14192_ ;
	wire _w14191_ ;
	wire _w14190_ ;
	wire _w14189_ ;
	wire _w14188_ ;
	wire _w14187_ ;
	wire _w14186_ ;
	wire _w14185_ ;
	wire _w14184_ ;
	wire _w14183_ ;
	wire _w14182_ ;
	wire _w14181_ ;
	wire _w14180_ ;
	wire _w14179_ ;
	wire _w14178_ ;
	wire _w14177_ ;
	wire _w14176_ ;
	wire _w14175_ ;
	wire _w14174_ ;
	wire _w14173_ ;
	wire _w14172_ ;
	wire _w14171_ ;
	wire _w14170_ ;
	wire _w14169_ ;
	wire _w14168_ ;
	wire _w14167_ ;
	wire _w14166_ ;
	wire _w14165_ ;
	wire _w14164_ ;
	wire _w14163_ ;
	wire _w14162_ ;
	wire _w14161_ ;
	wire _w14160_ ;
	wire _w14159_ ;
	wire _w14158_ ;
	wire _w14157_ ;
	wire _w14156_ ;
	wire _w14155_ ;
	wire _w14154_ ;
	wire _w14153_ ;
	wire _w14152_ ;
	wire _w14151_ ;
	wire _w14150_ ;
	wire _w14149_ ;
	wire _w14148_ ;
	wire _w14147_ ;
	wire _w14146_ ;
	wire _w14145_ ;
	wire _w14144_ ;
	wire _w14143_ ;
	wire _w14142_ ;
	wire _w14141_ ;
	wire _w14140_ ;
	wire _w14139_ ;
	wire _w14138_ ;
	wire _w14137_ ;
	wire _w14136_ ;
	wire _w14135_ ;
	wire _w14134_ ;
	wire _w14133_ ;
	wire _w14132_ ;
	wire _w14131_ ;
	wire _w14130_ ;
	wire _w14129_ ;
	wire _w14128_ ;
	wire _w14127_ ;
	wire _w14126_ ;
	wire _w14125_ ;
	wire _w14124_ ;
	wire _w14123_ ;
	wire _w14122_ ;
	wire _w14121_ ;
	wire _w14120_ ;
	wire _w14119_ ;
	wire _w14118_ ;
	wire _w14117_ ;
	wire _w14116_ ;
	wire _w14115_ ;
	wire _w14114_ ;
	wire _w14113_ ;
	wire _w14112_ ;
	wire _w14111_ ;
	wire _w14110_ ;
	wire _w14109_ ;
	wire _w14108_ ;
	wire _w14107_ ;
	wire _w14106_ ;
	wire _w14105_ ;
	wire _w14104_ ;
	wire _w14103_ ;
	wire _w14102_ ;
	wire _w14101_ ;
	wire _w14100_ ;
	wire _w14099_ ;
	wire _w14098_ ;
	wire _w14097_ ;
	wire _w14096_ ;
	wire _w14095_ ;
	wire _w14094_ ;
	wire _w14093_ ;
	wire _w14092_ ;
	wire _w14091_ ;
	wire _w14090_ ;
	wire _w14089_ ;
	wire _w14088_ ;
	wire _w14087_ ;
	wire _w14086_ ;
	wire _w14085_ ;
	wire _w14084_ ;
	wire _w14083_ ;
	wire _w14082_ ;
	wire _w14081_ ;
	wire _w14080_ ;
	wire _w14079_ ;
	wire _w14078_ ;
	wire _w14077_ ;
	wire _w14076_ ;
	wire _w14075_ ;
	wire _w14074_ ;
	wire _w14073_ ;
	wire _w14072_ ;
	wire _w14071_ ;
	wire _w14070_ ;
	wire _w14069_ ;
	wire _w14068_ ;
	wire _w14067_ ;
	wire _w14066_ ;
	wire _w14065_ ;
	wire _w14064_ ;
	wire _w14063_ ;
	wire _w14062_ ;
	wire _w14061_ ;
	wire _w14060_ ;
	wire _w14059_ ;
	wire _w14058_ ;
	wire _w14057_ ;
	wire _w14056_ ;
	wire _w14055_ ;
	wire _w14054_ ;
	wire _w14053_ ;
	wire _w14052_ ;
	wire _w14051_ ;
	wire _w14050_ ;
	wire _w14049_ ;
	wire _w14048_ ;
	wire _w14047_ ;
	wire _w14046_ ;
	wire _w14045_ ;
	wire _w14044_ ;
	wire _w14043_ ;
	wire _w14042_ ;
	wire _w14041_ ;
	wire _w14040_ ;
	wire _w14039_ ;
	wire _w14038_ ;
	wire _w14037_ ;
	wire _w14036_ ;
	wire _w14035_ ;
	wire _w14034_ ;
	wire _w14033_ ;
	wire _w14032_ ;
	wire _w14031_ ;
	wire _w14030_ ;
	wire _w14029_ ;
	wire _w14028_ ;
	wire _w14027_ ;
	wire _w14026_ ;
	wire _w14025_ ;
	wire _w14024_ ;
	wire _w14023_ ;
	wire _w14022_ ;
	wire _w14021_ ;
	wire _w14020_ ;
	wire _w14019_ ;
	wire _w14018_ ;
	wire _w14017_ ;
	wire _w14016_ ;
	wire _w14015_ ;
	wire _w14014_ ;
	wire _w14013_ ;
	wire _w14012_ ;
	wire _w14011_ ;
	wire _w14010_ ;
	wire _w14009_ ;
	wire _w14008_ ;
	wire _w14007_ ;
	wire _w14006_ ;
	wire _w14005_ ;
	wire _w14004_ ;
	wire _w14003_ ;
	wire _w14002_ ;
	wire _w14001_ ;
	wire _w14000_ ;
	wire _w13999_ ;
	wire _w13998_ ;
	wire _w13997_ ;
	wire _w13996_ ;
	wire _w13995_ ;
	wire _w13994_ ;
	wire _w13993_ ;
	wire _w13992_ ;
	wire _w13991_ ;
	wire _w13990_ ;
	wire _w13989_ ;
	wire _w13988_ ;
	wire _w13987_ ;
	wire _w13986_ ;
	wire _w13985_ ;
	wire _w13984_ ;
	wire _w13983_ ;
	wire _w13982_ ;
	wire _w13981_ ;
	wire _w13980_ ;
	wire _w13979_ ;
	wire _w13978_ ;
	wire _w13977_ ;
	wire _w13976_ ;
	wire _w13975_ ;
	wire _w13974_ ;
	wire _w13973_ ;
	wire _w13972_ ;
	wire _w13971_ ;
	wire _w13970_ ;
	wire _w13969_ ;
	wire _w13968_ ;
	wire _w13967_ ;
	wire _w13966_ ;
	wire _w13965_ ;
	wire _w13964_ ;
	wire _w13963_ ;
	wire _w13962_ ;
	wire _w13961_ ;
	wire _w13960_ ;
	wire _w13959_ ;
	wire _w13958_ ;
	wire _w13957_ ;
	wire _w13956_ ;
	wire _w13955_ ;
	wire _w13954_ ;
	wire _w13953_ ;
	wire _w13952_ ;
	wire _w13951_ ;
	wire _w13950_ ;
	wire _w13949_ ;
	wire _w13948_ ;
	wire _w13947_ ;
	wire _w13946_ ;
	wire _w13945_ ;
	wire _w13944_ ;
	wire _w13943_ ;
	wire _w13942_ ;
	wire _w13941_ ;
	wire _w13940_ ;
	wire _w13939_ ;
	wire _w13938_ ;
	wire _w13937_ ;
	wire _w13936_ ;
	wire _w13935_ ;
	wire _w13934_ ;
	wire _w13933_ ;
	wire _w13932_ ;
	wire _w13931_ ;
	wire _w13930_ ;
	wire _w13929_ ;
	wire _w13928_ ;
	wire _w13927_ ;
	wire _w13926_ ;
	wire _w13925_ ;
	wire _w13924_ ;
	wire _w13923_ ;
	wire _w13922_ ;
	wire _w13921_ ;
	wire _w13920_ ;
	wire _w13919_ ;
	wire _w13918_ ;
	wire _w13917_ ;
	wire _w13916_ ;
	wire _w13915_ ;
	wire _w13914_ ;
	wire _w13913_ ;
	wire _w13912_ ;
	wire _w13911_ ;
	wire _w13910_ ;
	wire _w13909_ ;
	wire _w13908_ ;
	wire _w13907_ ;
	wire _w13906_ ;
	wire _w13905_ ;
	wire _w13904_ ;
	wire _w13903_ ;
	wire _w13902_ ;
	wire _w13901_ ;
	wire _w13900_ ;
	wire _w13899_ ;
	wire _w13898_ ;
	wire _w13897_ ;
	wire _w13896_ ;
	wire _w13895_ ;
	wire _w13894_ ;
	wire _w13893_ ;
	wire _w13892_ ;
	wire _w13891_ ;
	wire _w13890_ ;
	wire _w13889_ ;
	wire _w13888_ ;
	wire _w13887_ ;
	wire _w13886_ ;
	wire _w13885_ ;
	wire _w13884_ ;
	wire _w13883_ ;
	wire _w13882_ ;
	wire _w13881_ ;
	wire _w13880_ ;
	wire _w13879_ ;
	wire _w13878_ ;
	wire _w13877_ ;
	wire _w13876_ ;
	wire _w13875_ ;
	wire _w13874_ ;
	wire _w13873_ ;
	wire _w13872_ ;
	wire _w13871_ ;
	wire _w13870_ ;
	wire _w13869_ ;
	wire _w13868_ ;
	wire _w13867_ ;
	wire _w13866_ ;
	wire _w13865_ ;
	wire _w13864_ ;
	wire _w13863_ ;
	wire _w13862_ ;
	wire _w13861_ ;
	wire _w13860_ ;
	wire _w13859_ ;
	wire _w13858_ ;
	wire _w13857_ ;
	wire _w13856_ ;
	wire _w13855_ ;
	wire _w13854_ ;
	wire _w13853_ ;
	wire _w13852_ ;
	wire _w13851_ ;
	wire _w13850_ ;
	wire _w13849_ ;
	wire _w13848_ ;
	wire _w13847_ ;
	wire _w13846_ ;
	wire _w13845_ ;
	wire _w13844_ ;
	wire _w13843_ ;
	wire _w13842_ ;
	wire _w13841_ ;
	wire _w13840_ ;
	wire _w13839_ ;
	wire _w13838_ ;
	wire _w13837_ ;
	wire _w13836_ ;
	wire _w13835_ ;
	wire _w13834_ ;
	wire _w13833_ ;
	wire _w13832_ ;
	wire _w13831_ ;
	wire _w13830_ ;
	wire _w13829_ ;
	wire _w13828_ ;
	wire _w13827_ ;
	wire _w13826_ ;
	wire _w13825_ ;
	wire _w13824_ ;
	wire _w13823_ ;
	wire _w13822_ ;
	wire _w13821_ ;
	wire _w13820_ ;
	wire _w13819_ ;
	wire _w13818_ ;
	wire _w13817_ ;
	wire _w13816_ ;
	wire _w13815_ ;
	wire _w13814_ ;
	wire _w13813_ ;
	wire _w13812_ ;
	wire _w13811_ ;
	wire _w13810_ ;
	wire _w13809_ ;
	wire _w13808_ ;
	wire _w13807_ ;
	wire _w13806_ ;
	wire _w13805_ ;
	wire _w13804_ ;
	wire _w13803_ ;
	wire _w13802_ ;
	wire _w13801_ ;
	wire _w13800_ ;
	wire _w13799_ ;
	wire _w13798_ ;
	wire _w13797_ ;
	wire _w13796_ ;
	wire _w13795_ ;
	wire _w13794_ ;
	wire _w13793_ ;
	wire _w13792_ ;
	wire _w13791_ ;
	wire _w13790_ ;
	wire _w13789_ ;
	wire _w13788_ ;
	wire _w13787_ ;
	wire _w13786_ ;
	wire _w13785_ ;
	wire _w13784_ ;
	wire _w13783_ ;
	wire _w13782_ ;
	wire _w13781_ ;
	wire _w13780_ ;
	wire _w13779_ ;
	wire _w13778_ ;
	wire _w13777_ ;
	wire _w13776_ ;
	wire _w13775_ ;
	wire _w13774_ ;
	wire _w13773_ ;
	wire _w13772_ ;
	wire _w13771_ ;
	wire _w13770_ ;
	wire _w13769_ ;
	wire _w13768_ ;
	wire _w13767_ ;
	wire _w13766_ ;
	wire _w13765_ ;
	wire _w13764_ ;
	wire _w13763_ ;
	wire _w13762_ ;
	wire _w13761_ ;
	wire _w13760_ ;
	wire _w13759_ ;
	wire _w13758_ ;
	wire _w13757_ ;
	wire _w13756_ ;
	wire _w13755_ ;
	wire _w13754_ ;
	wire _w13753_ ;
	wire _w13752_ ;
	wire _w13751_ ;
	wire _w13750_ ;
	wire _w13749_ ;
	wire _w13748_ ;
	wire _w13747_ ;
	wire _w13746_ ;
	wire _w13745_ ;
	wire _w13744_ ;
	wire _w13743_ ;
	wire _w13742_ ;
	wire _w13741_ ;
	wire _w13740_ ;
	wire _w13739_ ;
	wire _w13738_ ;
	wire _w13737_ ;
	wire _w13736_ ;
	wire _w13735_ ;
	wire _w13734_ ;
	wire _w13733_ ;
	wire _w13732_ ;
	wire _w13731_ ;
	wire _w13730_ ;
	wire _w13729_ ;
	wire _w13728_ ;
	wire _w13727_ ;
	wire _w13726_ ;
	wire _w13725_ ;
	wire _w13724_ ;
	wire _w13723_ ;
	wire _w13722_ ;
	wire _w13721_ ;
	wire _w13720_ ;
	wire _w13719_ ;
	wire _w13718_ ;
	wire _w13717_ ;
	wire _w13716_ ;
	wire _w13715_ ;
	wire _w13714_ ;
	wire _w13713_ ;
	wire _w13712_ ;
	wire _w13711_ ;
	wire _w13710_ ;
	wire _w13709_ ;
	wire _w13708_ ;
	wire _w13707_ ;
	wire _w13706_ ;
	wire _w13705_ ;
	wire _w13704_ ;
	wire _w13703_ ;
	wire _w13702_ ;
	wire _w13701_ ;
	wire _w13700_ ;
	wire _w13699_ ;
	wire _w13698_ ;
	wire _w13697_ ;
	wire _w13696_ ;
	wire _w13695_ ;
	wire _w13694_ ;
	wire _w13693_ ;
	wire _w13692_ ;
	wire _w13691_ ;
	wire _w13690_ ;
	wire _w13689_ ;
	wire _w13688_ ;
	wire _w13687_ ;
	wire _w13686_ ;
	wire _w13685_ ;
	wire _w13684_ ;
	wire _w13683_ ;
	wire _w13682_ ;
	wire _w13681_ ;
	wire _w13680_ ;
	wire _w13679_ ;
	wire _w13678_ ;
	wire _w13677_ ;
	wire _w13676_ ;
	wire _w13675_ ;
	wire _w13674_ ;
	wire _w13673_ ;
	wire _w13672_ ;
	wire _w13671_ ;
	wire _w13670_ ;
	wire _w13669_ ;
	wire _w13668_ ;
	wire _w13667_ ;
	wire _w13666_ ;
	wire _w13665_ ;
	wire _w13664_ ;
	wire _w13663_ ;
	wire _w13662_ ;
	wire _w13661_ ;
	wire _w13660_ ;
	wire _w13659_ ;
	wire _w13658_ ;
	wire _w13657_ ;
	wire _w13656_ ;
	wire _w13655_ ;
	wire _w13654_ ;
	wire _w13653_ ;
	wire _w13652_ ;
	wire _w13651_ ;
	wire _w13650_ ;
	wire _w13649_ ;
	wire _w13648_ ;
	wire _w13647_ ;
	wire _w13646_ ;
	wire _w13645_ ;
	wire _w13644_ ;
	wire _w13643_ ;
	wire _w13642_ ;
	wire _w13641_ ;
	wire _w13640_ ;
	wire _w13639_ ;
	wire _w13638_ ;
	wire _w13637_ ;
	wire _w13636_ ;
	wire _w13635_ ;
	wire _w13634_ ;
	wire _w13633_ ;
	wire _w13632_ ;
	wire _w13631_ ;
	wire _w13630_ ;
	wire _w13629_ ;
	wire _w13628_ ;
	wire _w13627_ ;
	wire _w13626_ ;
	wire _w13625_ ;
	wire _w13624_ ;
	wire _w13623_ ;
	wire _w13622_ ;
	wire _w13621_ ;
	wire _w13620_ ;
	wire _w13619_ ;
	wire _w13618_ ;
	wire _w13617_ ;
	wire _w13616_ ;
	wire _w13615_ ;
	wire _w13614_ ;
	wire _w13613_ ;
	wire _w13612_ ;
	wire _w13611_ ;
	wire _w13610_ ;
	wire _w13609_ ;
	wire _w13608_ ;
	wire _w13607_ ;
	wire _w13606_ ;
	wire _w13605_ ;
	wire _w13604_ ;
	wire _w13603_ ;
	wire _w13602_ ;
	wire _w13601_ ;
	wire _w13600_ ;
	wire _w13599_ ;
	wire _w13598_ ;
	wire _w13597_ ;
	wire _w13596_ ;
	wire _w13595_ ;
	wire _w13594_ ;
	wire _w13593_ ;
	wire _w13592_ ;
	wire _w13591_ ;
	wire _w13590_ ;
	wire _w13589_ ;
	wire _w13588_ ;
	wire _w13587_ ;
	wire _w13586_ ;
	wire _w13585_ ;
	wire _w13584_ ;
	wire _w13583_ ;
	wire _w13582_ ;
	wire _w13581_ ;
	wire _w13580_ ;
	wire _w13579_ ;
	wire _w13578_ ;
	wire _w13577_ ;
	wire _w13576_ ;
	wire _w13575_ ;
	wire _w13574_ ;
	wire _w13573_ ;
	wire _w13572_ ;
	wire _w13571_ ;
	wire _w13570_ ;
	wire _w13569_ ;
	wire _w13568_ ;
	wire _w13567_ ;
	wire _w13566_ ;
	wire _w13565_ ;
	wire _w13564_ ;
	wire _w13563_ ;
	wire _w13562_ ;
	wire _w13561_ ;
	wire _w13560_ ;
	wire _w13559_ ;
	wire _w13558_ ;
	wire _w13557_ ;
	wire _w13556_ ;
	wire _w13555_ ;
	wire _w13554_ ;
	wire _w13553_ ;
	wire _w13552_ ;
	wire _w13551_ ;
	wire _w13550_ ;
	wire _w13549_ ;
	wire _w13548_ ;
	wire _w13547_ ;
	wire _w13546_ ;
	wire _w13545_ ;
	wire _w13544_ ;
	wire _w13543_ ;
	wire _w13542_ ;
	wire _w13541_ ;
	wire _w13540_ ;
	wire _w13539_ ;
	wire _w13538_ ;
	wire _w13537_ ;
	wire _w13536_ ;
	wire _w13535_ ;
	wire _w13534_ ;
	wire _w13533_ ;
	wire _w13532_ ;
	wire _w13531_ ;
	wire _w13530_ ;
	wire _w13529_ ;
	wire _w13528_ ;
	wire _w13527_ ;
	wire _w13526_ ;
	wire _w13525_ ;
	wire _w13524_ ;
	wire _w13523_ ;
	wire _w13522_ ;
	wire _w13521_ ;
	wire _w13520_ ;
	wire _w13519_ ;
	wire _w13518_ ;
	wire _w13517_ ;
	wire _w13516_ ;
	wire _w13515_ ;
	wire _w13514_ ;
	wire _w13513_ ;
	wire _w13512_ ;
	wire _w13511_ ;
	wire _w13510_ ;
	wire _w13509_ ;
	wire _w13508_ ;
	wire _w13507_ ;
	wire _w13506_ ;
	wire _w13505_ ;
	wire _w13504_ ;
	wire _w13503_ ;
	wire _w13502_ ;
	wire _w13501_ ;
	wire _w13500_ ;
	wire _w13499_ ;
	wire _w13498_ ;
	wire _w13497_ ;
	wire _w13496_ ;
	wire _w13495_ ;
	wire _w13494_ ;
	wire _w13493_ ;
	wire _w13492_ ;
	wire _w13491_ ;
	wire _w13490_ ;
	wire _w13489_ ;
	wire _w13488_ ;
	wire _w13487_ ;
	wire _w13486_ ;
	wire _w13485_ ;
	wire _w13484_ ;
	wire _w13483_ ;
	wire _w13482_ ;
	wire _w13481_ ;
	wire _w13480_ ;
	wire _w13479_ ;
	wire _w13478_ ;
	wire _w13477_ ;
	wire _w13476_ ;
	wire _w13475_ ;
	wire _w13474_ ;
	wire _w13473_ ;
	wire _w13472_ ;
	wire _w13471_ ;
	wire _w13470_ ;
	wire _w13469_ ;
	wire _w13468_ ;
	wire _w13467_ ;
	wire _w13466_ ;
	wire _w13465_ ;
	wire _w13464_ ;
	wire _w13463_ ;
	wire _w13462_ ;
	wire _w13461_ ;
	wire _w13460_ ;
	wire _w13459_ ;
	wire _w13458_ ;
	wire _w13457_ ;
	wire _w13456_ ;
	wire _w13455_ ;
	wire _w13454_ ;
	wire _w13453_ ;
	wire _w13452_ ;
	wire _w13451_ ;
	wire _w13450_ ;
	wire _w13449_ ;
	wire _w13448_ ;
	wire _w13447_ ;
	wire _w13446_ ;
	wire _w13445_ ;
	wire _w13444_ ;
	wire _w13443_ ;
	wire _w13442_ ;
	wire _w13441_ ;
	wire _w13440_ ;
	wire _w13439_ ;
	wire _w13438_ ;
	wire _w13437_ ;
	wire _w13436_ ;
	wire _w13435_ ;
	wire _w13434_ ;
	wire _w13433_ ;
	wire _w13432_ ;
	wire _w13431_ ;
	wire _w13430_ ;
	wire _w13429_ ;
	wire _w13428_ ;
	wire _w13427_ ;
	wire _w13426_ ;
	wire _w13425_ ;
	wire _w13424_ ;
	wire _w13423_ ;
	wire _w13422_ ;
	wire _w13421_ ;
	wire _w13420_ ;
	wire _w13419_ ;
	wire _w13418_ ;
	wire _w13417_ ;
	wire _w13416_ ;
	wire _w13415_ ;
	wire _w13414_ ;
	wire _w13413_ ;
	wire _w13412_ ;
	wire _w13411_ ;
	wire _w13410_ ;
	wire _w13409_ ;
	wire _w13408_ ;
	wire _w13407_ ;
	wire _w13406_ ;
	wire _w13405_ ;
	wire _w13404_ ;
	wire _w13403_ ;
	wire _w13402_ ;
	wire _w13401_ ;
	wire _w13400_ ;
	wire _w13399_ ;
	wire _w13398_ ;
	wire _w13397_ ;
	wire _w13396_ ;
	wire _w13395_ ;
	wire _w13394_ ;
	wire _w13393_ ;
	wire _w13392_ ;
	wire _w13391_ ;
	wire _w13390_ ;
	wire _w13389_ ;
	wire _w13388_ ;
	wire _w13387_ ;
	wire _w13386_ ;
	wire _w13385_ ;
	wire _w13384_ ;
	wire _w13383_ ;
	wire _w13382_ ;
	wire _w13381_ ;
	wire _w13380_ ;
	wire _w13379_ ;
	wire _w13378_ ;
	wire _w13377_ ;
	wire _w13376_ ;
	wire _w13375_ ;
	wire _w13374_ ;
	wire _w13373_ ;
	wire _w13372_ ;
	wire _w13371_ ;
	wire _w13370_ ;
	wire _w13369_ ;
	wire _w13368_ ;
	wire _w13367_ ;
	wire _w13366_ ;
	wire _w13365_ ;
	wire _w13364_ ;
	wire _w13363_ ;
	wire _w13362_ ;
	wire _w13361_ ;
	wire _w13360_ ;
	wire _w13359_ ;
	wire _w13358_ ;
	wire _w13357_ ;
	wire _w13356_ ;
	wire _w13355_ ;
	wire _w13354_ ;
	wire _w13353_ ;
	wire _w13352_ ;
	wire _w13351_ ;
	wire _w13350_ ;
	wire _w13349_ ;
	wire _w13348_ ;
	wire _w13347_ ;
	wire _w13346_ ;
	wire _w13345_ ;
	wire _w13344_ ;
	wire _w13343_ ;
	wire _w13342_ ;
	wire _w13341_ ;
	wire _w13340_ ;
	wire _w13339_ ;
	wire _w13338_ ;
	wire _w13337_ ;
	wire _w13336_ ;
	wire _w13335_ ;
	wire _w13334_ ;
	wire _w13333_ ;
	wire _w13332_ ;
	wire _w13331_ ;
	wire _w13330_ ;
	wire _w13329_ ;
	wire _w13328_ ;
	wire _w13327_ ;
	wire _w13326_ ;
	wire _w13325_ ;
	wire _w13324_ ;
	wire _w13323_ ;
	wire _w13322_ ;
	wire _w13321_ ;
	wire _w13320_ ;
	wire _w13319_ ;
	wire _w13318_ ;
	wire _w13317_ ;
	wire _w13316_ ;
	wire _w13315_ ;
	wire _w13314_ ;
	wire _w13313_ ;
	wire _w13312_ ;
	wire _w13311_ ;
	wire _w13310_ ;
	wire _w13309_ ;
	wire _w13308_ ;
	wire _w13307_ ;
	wire _w13306_ ;
	wire _w13305_ ;
	wire _w13304_ ;
	wire _w13303_ ;
	wire _w13302_ ;
	wire _w13301_ ;
	wire _w13300_ ;
	wire _w13299_ ;
	wire _w13298_ ;
	wire _w13297_ ;
	wire _w13296_ ;
	wire _w13295_ ;
	wire _w13294_ ;
	wire _w13293_ ;
	wire _w13292_ ;
	wire _w13291_ ;
	wire _w13290_ ;
	wire _w13289_ ;
	wire _w13288_ ;
	wire _w13287_ ;
	wire _w13286_ ;
	wire _w13285_ ;
	wire _w13284_ ;
	wire _w13283_ ;
	wire _w13282_ ;
	wire _w13281_ ;
	wire _w13280_ ;
	wire _w13279_ ;
	wire _w13278_ ;
	wire _w13277_ ;
	wire _w13276_ ;
	wire _w13275_ ;
	wire _w13274_ ;
	wire _w13273_ ;
	wire _w13272_ ;
	wire _w13271_ ;
	wire _w13270_ ;
	wire _w13269_ ;
	wire _w13268_ ;
	wire _w13267_ ;
	wire _w13266_ ;
	wire _w13265_ ;
	wire _w13264_ ;
	wire _w13263_ ;
	wire _w13262_ ;
	wire _w13261_ ;
	wire _w13260_ ;
	wire _w13259_ ;
	wire _w13258_ ;
	wire _w13257_ ;
	wire _w13256_ ;
	wire _w13255_ ;
	wire _w13254_ ;
	wire _w13253_ ;
	wire _w13252_ ;
	wire _w13251_ ;
	wire _w13250_ ;
	wire _w13249_ ;
	wire _w13248_ ;
	wire _w13247_ ;
	wire _w13246_ ;
	wire _w13245_ ;
	wire _w13244_ ;
	wire _w13243_ ;
	wire _w13242_ ;
	wire _w13241_ ;
	wire _w13240_ ;
	wire _w13239_ ;
	wire _w13238_ ;
	wire _w13237_ ;
	wire _w13236_ ;
	wire _w13235_ ;
	wire _w13234_ ;
	wire _w13233_ ;
	wire _w13232_ ;
	wire _w13231_ ;
	wire _w13230_ ;
	wire _w13229_ ;
	wire _w13228_ ;
	wire _w13227_ ;
	wire _w13226_ ;
	wire _w13225_ ;
	wire _w13224_ ;
	wire _w13223_ ;
	wire _w13222_ ;
	wire _w13221_ ;
	wire _w13220_ ;
	wire _w13219_ ;
	wire _w13218_ ;
	wire _w13217_ ;
	wire _w13216_ ;
	wire _w13215_ ;
	wire _w13214_ ;
	wire _w13213_ ;
	wire _w13212_ ;
	wire _w13211_ ;
	wire _w13210_ ;
	wire _w13209_ ;
	wire _w13208_ ;
	wire _w13207_ ;
	wire _w13206_ ;
	wire _w13205_ ;
	wire _w13204_ ;
	wire _w13203_ ;
	wire _w13202_ ;
	wire _w13201_ ;
	wire _w13200_ ;
	wire _w13199_ ;
	wire _w13198_ ;
	wire _w13197_ ;
	wire _w13196_ ;
	wire _w13195_ ;
	wire _w13194_ ;
	wire _w13193_ ;
	wire _w13192_ ;
	wire _w13191_ ;
	wire _w13190_ ;
	wire _w13189_ ;
	wire _w13188_ ;
	wire _w13187_ ;
	wire _w13186_ ;
	wire _w13185_ ;
	wire _w13184_ ;
	wire _w13183_ ;
	wire _w13182_ ;
	wire _w13181_ ;
	wire _w13180_ ;
	wire _w13179_ ;
	wire _w13178_ ;
	wire _w13177_ ;
	wire _w13176_ ;
	wire _w13175_ ;
	wire _w13174_ ;
	wire _w13173_ ;
	wire _w13172_ ;
	wire _w13171_ ;
	wire _w13170_ ;
	wire _w13169_ ;
	wire _w13168_ ;
	wire _w13167_ ;
	wire _w13166_ ;
	wire _w13165_ ;
	wire _w13164_ ;
	wire _w13163_ ;
	wire _w13162_ ;
	wire _w13161_ ;
	wire _w13160_ ;
	wire _w13159_ ;
	wire _w13158_ ;
	wire _w13157_ ;
	wire _w13156_ ;
	wire _w13155_ ;
	wire _w13154_ ;
	wire _w13153_ ;
	wire _w13152_ ;
	wire _w13151_ ;
	wire _w13150_ ;
	wire _w13149_ ;
	wire _w13148_ ;
	wire _w13147_ ;
	wire _w13146_ ;
	wire _w13145_ ;
	wire _w13144_ ;
	wire _w13143_ ;
	wire _w13142_ ;
	wire _w13141_ ;
	wire _w13140_ ;
	wire _w13139_ ;
	wire _w13138_ ;
	wire _w13137_ ;
	wire _w13136_ ;
	wire _w13135_ ;
	wire _w13134_ ;
	wire _w13133_ ;
	wire _w13132_ ;
	wire _w13131_ ;
	wire _w13130_ ;
	wire _w13129_ ;
	wire _w13128_ ;
	wire _w13127_ ;
	wire _w13126_ ;
	wire _w13125_ ;
	wire _w13124_ ;
	wire _w13123_ ;
	wire _w13122_ ;
	wire _w13121_ ;
	wire _w13120_ ;
	wire _w13119_ ;
	wire _w13118_ ;
	wire _w13117_ ;
	wire _w13116_ ;
	wire _w13115_ ;
	wire _w13114_ ;
	wire _w13113_ ;
	wire _w13112_ ;
	wire _w13111_ ;
	wire _w13110_ ;
	wire _w13109_ ;
	wire _w13108_ ;
	wire _w13107_ ;
	wire _w13106_ ;
	wire _w13105_ ;
	wire _w13104_ ;
	wire _w13103_ ;
	wire _w13102_ ;
	wire _w13101_ ;
	wire _w13100_ ;
	wire _w13099_ ;
	wire _w13098_ ;
	wire _w13097_ ;
	wire _w13096_ ;
	wire _w13095_ ;
	wire _w13094_ ;
	wire _w13093_ ;
	wire _w13092_ ;
	wire _w13091_ ;
	wire _w13090_ ;
	wire _w13089_ ;
	wire _w13088_ ;
	wire _w13087_ ;
	wire _w13086_ ;
	wire _w13085_ ;
	wire _w13084_ ;
	wire _w13083_ ;
	wire _w13082_ ;
	wire _w13081_ ;
	wire _w13080_ ;
	wire _w13079_ ;
	wire _w13078_ ;
	wire _w13077_ ;
	wire _w13076_ ;
	wire _w13075_ ;
	wire _w13074_ ;
	wire _w13073_ ;
	wire _w13072_ ;
	wire _w13071_ ;
	wire _w13070_ ;
	wire _w13069_ ;
	wire _w13068_ ;
	wire _w13067_ ;
	wire _w13066_ ;
	wire _w13065_ ;
	wire _w13064_ ;
	wire _w13063_ ;
	wire _w13062_ ;
	wire _w13061_ ;
	wire _w13060_ ;
	wire _w13059_ ;
	wire _w13058_ ;
	wire _w13057_ ;
	wire _w13056_ ;
	wire _w13055_ ;
	wire _w13054_ ;
	wire _w13053_ ;
	wire _w13052_ ;
	wire _w13051_ ;
	wire _w13050_ ;
	wire _w13049_ ;
	wire _w13048_ ;
	wire _w13047_ ;
	wire _w13046_ ;
	wire _w13045_ ;
	wire _w13044_ ;
	wire _w13043_ ;
	wire _w13042_ ;
	wire _w13041_ ;
	wire _w13040_ ;
	wire _w13039_ ;
	wire _w13038_ ;
	wire _w13037_ ;
	wire _w13036_ ;
	wire _w13035_ ;
	wire _w13034_ ;
	wire _w13033_ ;
	wire _w13032_ ;
	wire _w13031_ ;
	wire _w13030_ ;
	wire _w13029_ ;
	wire _w13028_ ;
	wire _w13027_ ;
	wire _w13026_ ;
	wire _w13025_ ;
	wire _w13024_ ;
	wire _w13023_ ;
	wire _w13022_ ;
	wire _w13021_ ;
	wire _w13020_ ;
	wire _w13019_ ;
	wire _w13018_ ;
	wire _w13017_ ;
	wire _w13016_ ;
	wire _w13015_ ;
	wire _w13014_ ;
	wire _w13013_ ;
	wire _w13012_ ;
	wire _w13011_ ;
	wire _w13010_ ;
	wire _w13009_ ;
	wire _w13008_ ;
	wire _w13007_ ;
	wire _w13006_ ;
	wire _w13005_ ;
	wire _w13004_ ;
	wire _w13003_ ;
	wire _w13002_ ;
	wire _w13001_ ;
	wire _w13000_ ;
	wire _w12999_ ;
	wire _w12998_ ;
	wire _w12997_ ;
	wire _w12996_ ;
	wire _w12995_ ;
	wire _w12994_ ;
	wire _w12993_ ;
	wire _w12992_ ;
	wire _w12991_ ;
	wire _w12990_ ;
	wire _w12989_ ;
	wire _w12988_ ;
	wire _w12987_ ;
	wire _w12986_ ;
	wire _w12985_ ;
	wire _w12984_ ;
	wire _w12983_ ;
	wire _w12982_ ;
	wire _w12981_ ;
	wire _w12980_ ;
	wire _w12979_ ;
	wire _w12978_ ;
	wire _w12977_ ;
	wire _w12976_ ;
	wire _w12975_ ;
	wire _w12974_ ;
	wire _w12973_ ;
	wire _w12972_ ;
	wire _w12971_ ;
	wire _w12970_ ;
	wire _w12969_ ;
	wire _w12968_ ;
	wire _w12967_ ;
	wire _w12966_ ;
	wire _w12965_ ;
	wire _w12964_ ;
	wire _w12963_ ;
	wire _w12962_ ;
	wire _w12961_ ;
	wire _w12960_ ;
	wire _w12959_ ;
	wire _w12958_ ;
	wire _w12957_ ;
	wire _w12956_ ;
	wire _w12955_ ;
	wire _w12954_ ;
	wire _w12953_ ;
	wire _w12952_ ;
	wire _w12951_ ;
	wire _w12950_ ;
	wire _w12949_ ;
	wire _w12948_ ;
	wire _w12947_ ;
	wire _w12946_ ;
	wire _w12945_ ;
	wire _w12944_ ;
	wire _w12943_ ;
	wire _w12942_ ;
	wire _w12941_ ;
	wire _w12940_ ;
	wire _w12939_ ;
	wire _w12938_ ;
	wire _w12937_ ;
	wire _w12936_ ;
	wire _w12935_ ;
	wire _w12934_ ;
	wire _w12933_ ;
	wire _w12932_ ;
	wire _w12931_ ;
	wire _w12930_ ;
	wire _w12929_ ;
	wire _w12928_ ;
	wire _w12927_ ;
	wire _w12926_ ;
	wire _w12925_ ;
	wire _w12924_ ;
	wire _w12923_ ;
	wire _w12922_ ;
	wire _w12921_ ;
	wire _w12920_ ;
	wire _w12919_ ;
	wire _w12918_ ;
	wire _w12917_ ;
	wire _w12916_ ;
	wire _w12915_ ;
	wire _w12914_ ;
	wire _w12913_ ;
	wire _w12912_ ;
	wire _w12911_ ;
	wire _w12910_ ;
	wire _w12909_ ;
	wire _w12908_ ;
	wire _w12907_ ;
	wire _w12906_ ;
	wire _w12905_ ;
	wire _w12904_ ;
	wire _w12903_ ;
	wire _w12902_ ;
	wire _w12901_ ;
	wire _w12900_ ;
	wire _w12899_ ;
	wire _w12898_ ;
	wire _w12897_ ;
	wire _w12896_ ;
	wire _w12895_ ;
	wire _w12894_ ;
	wire _w12893_ ;
	wire _w12892_ ;
	wire _w12891_ ;
	wire _w12890_ ;
	wire _w12889_ ;
	wire _w12888_ ;
	wire _w12887_ ;
	wire _w12886_ ;
	wire _w12885_ ;
	wire _w12884_ ;
	wire _w12883_ ;
	wire _w12882_ ;
	wire _w12881_ ;
	wire _w12880_ ;
	wire _w12879_ ;
	wire _w12878_ ;
	wire _w12877_ ;
	wire _w12876_ ;
	wire _w12875_ ;
	wire _w12874_ ;
	wire _w12873_ ;
	wire _w12872_ ;
	wire _w12871_ ;
	wire _w12870_ ;
	wire _w12869_ ;
	wire _w12868_ ;
	wire _w12867_ ;
	wire _w12866_ ;
	wire _w12865_ ;
	wire _w12864_ ;
	wire _w12863_ ;
	wire _w12862_ ;
	wire _w12861_ ;
	wire _w12860_ ;
	wire _w12859_ ;
	wire _w12858_ ;
	wire _w12857_ ;
	wire _w12856_ ;
	wire _w12855_ ;
	wire _w12854_ ;
	wire _w12853_ ;
	wire _w12852_ ;
	wire _w12851_ ;
	wire _w12850_ ;
	wire _w12849_ ;
	wire _w12848_ ;
	wire _w12847_ ;
	wire _w12846_ ;
	wire _w12845_ ;
	wire _w12844_ ;
	wire _w12843_ ;
	wire _w12842_ ;
	wire _w12841_ ;
	wire _w12840_ ;
	wire _w12839_ ;
	wire _w12838_ ;
	wire _w12837_ ;
	wire _w12836_ ;
	wire _w12835_ ;
	wire _w12834_ ;
	wire _w12833_ ;
	wire _w12832_ ;
	wire _w12831_ ;
	wire _w12830_ ;
	wire _w12829_ ;
	wire _w12828_ ;
	wire _w12827_ ;
	wire _w12826_ ;
	wire _w12825_ ;
	wire _w12824_ ;
	wire _w12823_ ;
	wire _w12822_ ;
	wire _w12821_ ;
	wire _w12820_ ;
	wire _w12819_ ;
	wire _w12818_ ;
	wire _w12817_ ;
	wire _w12816_ ;
	wire _w12815_ ;
	wire _w12814_ ;
	wire _w12813_ ;
	wire _w12812_ ;
	wire _w12811_ ;
	wire _w12810_ ;
	wire _w12809_ ;
	wire _w12808_ ;
	wire _w12807_ ;
	wire _w12806_ ;
	wire _w12805_ ;
	wire _w12804_ ;
	wire _w12803_ ;
	wire _w12802_ ;
	wire _w12801_ ;
	wire _w12800_ ;
	wire _w12799_ ;
	wire _w12798_ ;
	wire _w12797_ ;
	wire _w12796_ ;
	wire _w12795_ ;
	wire _w12794_ ;
	wire _w12793_ ;
	wire _w12792_ ;
	wire _w12791_ ;
	wire _w12790_ ;
	wire _w12789_ ;
	wire _w12788_ ;
	wire _w12787_ ;
	wire _w12786_ ;
	wire _w12785_ ;
	wire _w12784_ ;
	wire _w12783_ ;
	wire _w12782_ ;
	wire _w12781_ ;
	wire _w12780_ ;
	wire _w12779_ ;
	wire _w12778_ ;
	wire _w12777_ ;
	wire _w12776_ ;
	wire _w12775_ ;
	wire _w12774_ ;
	wire _w12773_ ;
	wire _w12772_ ;
	wire _w12771_ ;
	wire _w12770_ ;
	wire _w12769_ ;
	wire _w12768_ ;
	wire _w12767_ ;
	wire _w12766_ ;
	wire _w12765_ ;
	wire _w12764_ ;
	wire _w12763_ ;
	wire _w12762_ ;
	wire _w12761_ ;
	wire _w12760_ ;
	wire _w12759_ ;
	wire _w12758_ ;
	wire _w12757_ ;
	wire _w12756_ ;
	wire _w12755_ ;
	wire _w12754_ ;
	wire _w12753_ ;
	wire _w12752_ ;
	wire _w12751_ ;
	wire _w12750_ ;
	wire _w12749_ ;
	wire _w12748_ ;
	wire _w12747_ ;
	wire _w12746_ ;
	wire _w12745_ ;
	wire _w12744_ ;
	wire _w12743_ ;
	wire _w12742_ ;
	wire _w12741_ ;
	wire _w12740_ ;
	wire _w12739_ ;
	wire _w12738_ ;
	wire _w12737_ ;
	wire _w12736_ ;
	wire _w12735_ ;
	wire _w12734_ ;
	wire _w12733_ ;
	wire _w12732_ ;
	wire _w12731_ ;
	wire _w12730_ ;
	wire _w12729_ ;
	wire _w12728_ ;
	wire _w12727_ ;
	wire _w12726_ ;
	wire _w12725_ ;
	wire _w12724_ ;
	wire _w12723_ ;
	wire _w12722_ ;
	wire _w12721_ ;
	wire _w12720_ ;
	wire _w12719_ ;
	wire _w12718_ ;
	wire _w12717_ ;
	wire _w12716_ ;
	wire _w12715_ ;
	wire _w12714_ ;
	wire _w12713_ ;
	wire _w12712_ ;
	wire _w12711_ ;
	wire _w12710_ ;
	wire _w12709_ ;
	wire _w12708_ ;
	wire _w12707_ ;
	wire _w12706_ ;
	wire _w12705_ ;
	wire _w12704_ ;
	wire _w12703_ ;
	wire _w12702_ ;
	wire _w12701_ ;
	wire _w12700_ ;
	wire _w12699_ ;
	wire _w12698_ ;
	wire _w12697_ ;
	wire _w12696_ ;
	wire _w12695_ ;
	wire _w12694_ ;
	wire _w12693_ ;
	wire _w12692_ ;
	wire _w12691_ ;
	wire _w12690_ ;
	wire _w12689_ ;
	wire _w12688_ ;
	wire _w12687_ ;
	wire _w12686_ ;
	wire _w12685_ ;
	wire _w12684_ ;
	wire _w12683_ ;
	wire _w12682_ ;
	wire _w12681_ ;
	wire _w12680_ ;
	wire _w12679_ ;
	wire _w12678_ ;
	wire _w12677_ ;
	wire _w12676_ ;
	wire _w12675_ ;
	wire _w12674_ ;
	wire _w12673_ ;
	wire _w12672_ ;
	wire _w12671_ ;
	wire _w12670_ ;
	wire _w12669_ ;
	wire _w12668_ ;
	wire _w12667_ ;
	wire _w12666_ ;
	wire _w12665_ ;
	wire _w12664_ ;
	wire _w12663_ ;
	wire _w12662_ ;
	wire _w12661_ ;
	wire _w12660_ ;
	wire _w12659_ ;
	wire _w12658_ ;
	wire _w12657_ ;
	wire _w12656_ ;
	wire _w12655_ ;
	wire _w12654_ ;
	wire _w12653_ ;
	wire _w12652_ ;
	wire _w12651_ ;
	wire _w12650_ ;
	wire _w12649_ ;
	wire _w12648_ ;
	wire _w12647_ ;
	wire _w12646_ ;
	wire _w12645_ ;
	wire _w12644_ ;
	wire _w12643_ ;
	wire _w12642_ ;
	wire _w12641_ ;
	wire _w12640_ ;
	wire _w12639_ ;
	wire _w12638_ ;
	wire _w12637_ ;
	wire _w12636_ ;
	wire _w12635_ ;
	wire _w12634_ ;
	wire _w12633_ ;
	wire _w12632_ ;
	wire _w12631_ ;
	wire _w12630_ ;
	wire _w12629_ ;
	wire _w12628_ ;
	wire _w12627_ ;
	wire _w12626_ ;
	wire _w12625_ ;
	wire _w12624_ ;
	wire _w12623_ ;
	wire _w12622_ ;
	wire _w12621_ ;
	wire _w12620_ ;
	wire _w12619_ ;
	wire _w12618_ ;
	wire _w12617_ ;
	wire _w12616_ ;
	wire _w12615_ ;
	wire _w12614_ ;
	wire _w12613_ ;
	wire _w12612_ ;
	wire _w12611_ ;
	wire _w12610_ ;
	wire _w12609_ ;
	wire _w12608_ ;
	wire _w12607_ ;
	wire _w12606_ ;
	wire _w12605_ ;
	wire _w12604_ ;
	wire _w12603_ ;
	wire _w12602_ ;
	wire _w12601_ ;
	wire _w12600_ ;
	wire _w12599_ ;
	wire _w12598_ ;
	wire _w12597_ ;
	wire _w12596_ ;
	wire _w12595_ ;
	wire _w12594_ ;
	wire _w12593_ ;
	wire _w12592_ ;
	wire _w12591_ ;
	wire _w12590_ ;
	wire _w12589_ ;
	wire _w12588_ ;
	wire _w12587_ ;
	wire _w12586_ ;
	wire _w12585_ ;
	wire _w12584_ ;
	wire _w12583_ ;
	wire _w12582_ ;
	wire _w12581_ ;
	wire _w12580_ ;
	wire _w12579_ ;
	wire _w12578_ ;
	wire _w12577_ ;
	wire _w12576_ ;
	wire _w12575_ ;
	wire _w12574_ ;
	wire _w12573_ ;
	wire _w12572_ ;
	wire _w12571_ ;
	wire _w12570_ ;
	wire _w12569_ ;
	wire _w12568_ ;
	wire _w12567_ ;
	wire _w12566_ ;
	wire _w12565_ ;
	wire _w12564_ ;
	wire _w12563_ ;
	wire _w12562_ ;
	wire _w12561_ ;
	wire _w12560_ ;
	wire _w12559_ ;
	wire _w12558_ ;
	wire _w12557_ ;
	wire _w12556_ ;
	wire _w12555_ ;
	wire _w12554_ ;
	wire _w12553_ ;
	wire _w12552_ ;
	wire _w12551_ ;
	wire _w12550_ ;
	wire _w12549_ ;
	wire _w12548_ ;
	wire _w12547_ ;
	wire _w12546_ ;
	wire _w12545_ ;
	wire _w12544_ ;
	wire _w12543_ ;
	wire _w12542_ ;
	wire _w12541_ ;
	wire _w12540_ ;
	wire _w12539_ ;
	wire _w12538_ ;
	wire _w12537_ ;
	wire _w12536_ ;
	wire _w12535_ ;
	wire _w12534_ ;
	wire _w12533_ ;
	wire _w12532_ ;
	wire _w12531_ ;
	wire _w12530_ ;
	wire _w12529_ ;
	wire _w12528_ ;
	wire _w12527_ ;
	wire _w12526_ ;
	wire _w12525_ ;
	wire _w12524_ ;
	wire _w12523_ ;
	wire _w12522_ ;
	wire _w12521_ ;
	wire _w12520_ ;
	wire _w12519_ ;
	wire _w12518_ ;
	wire _w12517_ ;
	wire _w12516_ ;
	wire _w12515_ ;
	wire _w12514_ ;
	wire _w12513_ ;
	wire _w12512_ ;
	wire _w12511_ ;
	wire _w12510_ ;
	wire _w12509_ ;
	wire _w12508_ ;
	wire _w12507_ ;
	wire _w12506_ ;
	wire _w12505_ ;
	wire _w12504_ ;
	wire _w12503_ ;
	wire _w12502_ ;
	wire _w12501_ ;
	wire _w12500_ ;
	wire _w12499_ ;
	wire _w12498_ ;
	wire _w12497_ ;
	wire _w12496_ ;
	wire _w12495_ ;
	wire _w12494_ ;
	wire _w12493_ ;
	wire _w12492_ ;
	wire _w12491_ ;
	wire _w12490_ ;
	wire _w12489_ ;
	wire _w12488_ ;
	wire _w12487_ ;
	wire _w12486_ ;
	wire _w12485_ ;
	wire _w12484_ ;
	wire _w12483_ ;
	wire _w12482_ ;
	wire _w12481_ ;
	wire _w12480_ ;
	wire _w12479_ ;
	wire _w12478_ ;
	wire _w12477_ ;
	wire _w12476_ ;
	wire _w12475_ ;
	wire _w12474_ ;
	wire _w12473_ ;
	wire _w12472_ ;
	wire _w12471_ ;
	wire _w12470_ ;
	wire _w12469_ ;
	wire _w12468_ ;
	wire _w12467_ ;
	wire _w12466_ ;
	wire _w12465_ ;
	wire _w12464_ ;
	wire _w12463_ ;
	wire _w12462_ ;
	wire _w12461_ ;
	wire _w12460_ ;
	wire _w12459_ ;
	wire _w12458_ ;
	wire _w12457_ ;
	wire _w12456_ ;
	wire _w12455_ ;
	wire _w12454_ ;
	wire _w12453_ ;
	wire _w12452_ ;
	wire _w12451_ ;
	wire _w12450_ ;
	wire _w12449_ ;
	wire _w12448_ ;
	wire _w12447_ ;
	wire _w12446_ ;
	wire _w12445_ ;
	wire _w12444_ ;
	wire _w12443_ ;
	wire _w12442_ ;
	wire _w12441_ ;
	wire _w12440_ ;
	wire _w12439_ ;
	wire _w12438_ ;
	wire _w12437_ ;
	wire _w12436_ ;
	wire _w12435_ ;
	wire _w12434_ ;
	wire _w12433_ ;
	wire _w12432_ ;
	wire _w12431_ ;
	wire _w12430_ ;
	wire _w12429_ ;
	wire _w12428_ ;
	wire _w12427_ ;
	wire _w12426_ ;
	wire _w12425_ ;
	wire _w12424_ ;
	wire _w12423_ ;
	wire _w12422_ ;
	wire _w12421_ ;
	wire _w12420_ ;
	wire _w12419_ ;
	wire _w12418_ ;
	wire _w12417_ ;
	wire _w12416_ ;
	wire _w12415_ ;
	wire _w12414_ ;
	wire _w12413_ ;
	wire _w12412_ ;
	wire _w12411_ ;
	wire _w12410_ ;
	wire _w12409_ ;
	wire _w12408_ ;
	wire _w12407_ ;
	wire _w12406_ ;
	wire _w12405_ ;
	wire _w12404_ ;
	wire _w12403_ ;
	wire _w12402_ ;
	wire _w12401_ ;
	wire _w12400_ ;
	wire _w12399_ ;
	wire _w12398_ ;
	wire _w12397_ ;
	wire _w12396_ ;
	wire _w12395_ ;
	wire _w12394_ ;
	wire _w12393_ ;
	wire _w12392_ ;
	wire _w12391_ ;
	wire _w12390_ ;
	wire _w12389_ ;
	wire _w12388_ ;
	wire _w12387_ ;
	wire _w12386_ ;
	wire _w12385_ ;
	wire _w12384_ ;
	wire _w12383_ ;
	wire _w12382_ ;
	wire _w12381_ ;
	wire _w12380_ ;
	wire _w12379_ ;
	wire _w12378_ ;
	wire _w12377_ ;
	wire _w12376_ ;
	wire _w12375_ ;
	wire _w12374_ ;
	wire _w12373_ ;
	wire _w12372_ ;
	wire _w12371_ ;
	wire _w12370_ ;
	wire _w12369_ ;
	wire _w12368_ ;
	wire _w12367_ ;
	wire _w12366_ ;
	wire _w12365_ ;
	wire _w12364_ ;
	wire _w12363_ ;
	wire _w12362_ ;
	wire _w12361_ ;
	wire _w12360_ ;
	wire _w12359_ ;
	wire _w12358_ ;
	wire _w12357_ ;
	wire _w12356_ ;
	wire _w12355_ ;
	wire _w12354_ ;
	wire _w12353_ ;
	wire _w12352_ ;
	wire _w12351_ ;
	wire _w12350_ ;
	wire _w12349_ ;
	wire _w12348_ ;
	wire _w12347_ ;
	wire _w12346_ ;
	wire _w12345_ ;
	wire _w12344_ ;
	wire _w12343_ ;
	wire _w12342_ ;
	wire _w12341_ ;
	wire _w12340_ ;
	wire _w12339_ ;
	wire _w12338_ ;
	wire _w12337_ ;
	wire _w12336_ ;
	wire _w12335_ ;
	wire _w12334_ ;
	wire _w12333_ ;
	wire _w12332_ ;
	wire _w12331_ ;
	wire _w12330_ ;
	wire _w12329_ ;
	wire _w12328_ ;
	wire _w12327_ ;
	wire _w12326_ ;
	wire _w12325_ ;
	wire _w12324_ ;
	wire _w12323_ ;
	wire _w12322_ ;
	wire _w12321_ ;
	wire _w12320_ ;
	wire _w12319_ ;
	wire _w12318_ ;
	wire _w12317_ ;
	wire _w12316_ ;
	wire _w12315_ ;
	wire _w12314_ ;
	wire _w12313_ ;
	wire _w12312_ ;
	wire _w12311_ ;
	wire _w12310_ ;
	wire _w12309_ ;
	wire _w12308_ ;
	wire _w12307_ ;
	wire _w12306_ ;
	wire _w12305_ ;
	wire _w12304_ ;
	wire _w12303_ ;
	wire _w12302_ ;
	wire _w12301_ ;
	wire _w12300_ ;
	wire _w12299_ ;
	wire _w12298_ ;
	wire _w12297_ ;
	wire _w12296_ ;
	wire _w12295_ ;
	wire _w12294_ ;
	wire _w12293_ ;
	wire _w12292_ ;
	wire _w12291_ ;
	wire _w12290_ ;
	wire _w12289_ ;
	wire _w12288_ ;
	wire _w12287_ ;
	wire _w12286_ ;
	wire _w12285_ ;
	wire _w12284_ ;
	wire _w12283_ ;
	wire _w12282_ ;
	wire _w12281_ ;
	wire _w12280_ ;
	wire _w12279_ ;
	wire _w12278_ ;
	wire _w12277_ ;
	wire _w12276_ ;
	wire _w12275_ ;
	wire _w12274_ ;
	wire _w12273_ ;
	wire _w12272_ ;
	wire _w12271_ ;
	wire _w12270_ ;
	wire _w12269_ ;
	wire _w12268_ ;
	wire _w12267_ ;
	wire _w12266_ ;
	wire _w12265_ ;
	wire _w12264_ ;
	wire _w12263_ ;
	wire _w12262_ ;
	wire _w12261_ ;
	wire _w12260_ ;
	wire _w12259_ ;
	wire _w12258_ ;
	wire _w12257_ ;
	wire _w12256_ ;
	wire _w12255_ ;
	wire _w12254_ ;
	wire _w12253_ ;
	wire _w12252_ ;
	wire _w12251_ ;
	wire _w12250_ ;
	wire _w12249_ ;
	wire _w12248_ ;
	wire _w12247_ ;
	wire _w12246_ ;
	wire _w12245_ ;
	wire _w12244_ ;
	wire _w12243_ ;
	wire _w12242_ ;
	wire _w12241_ ;
	wire _w12240_ ;
	wire _w12239_ ;
	wire _w12238_ ;
	wire _w12237_ ;
	wire _w12236_ ;
	wire _w12235_ ;
	wire _w12234_ ;
	wire _w12233_ ;
	wire _w12232_ ;
	wire _w12231_ ;
	wire _w12230_ ;
	wire _w12229_ ;
	wire _w12228_ ;
	wire _w12227_ ;
	wire _w12226_ ;
	wire _w12225_ ;
	wire _w12224_ ;
	wire _w12223_ ;
	wire _w12222_ ;
	wire _w12221_ ;
	wire _w12220_ ;
	wire _w12219_ ;
	wire _w12218_ ;
	wire _w12217_ ;
	wire _w12216_ ;
	wire _w12215_ ;
	wire _w12214_ ;
	wire _w12213_ ;
	wire _w12212_ ;
	wire _w12211_ ;
	wire _w12210_ ;
	wire _w12209_ ;
	wire _w12208_ ;
	wire _w12207_ ;
	wire _w12206_ ;
	wire _w12205_ ;
	wire _w12204_ ;
	wire _w12203_ ;
	wire _w12202_ ;
	wire _w12201_ ;
	wire _w12200_ ;
	wire _w12199_ ;
	wire _w12198_ ;
	wire _w12197_ ;
	wire _w12196_ ;
	wire _w12195_ ;
	wire _w12194_ ;
	wire _w12193_ ;
	wire _w12192_ ;
	wire _w12191_ ;
	wire _w12190_ ;
	wire _w12189_ ;
	wire _w12188_ ;
	wire _w12187_ ;
	wire _w12186_ ;
	wire _w12185_ ;
	wire _w12184_ ;
	wire _w12183_ ;
	wire _w12182_ ;
	wire _w12181_ ;
	wire _w12180_ ;
	wire _w12179_ ;
	wire _w12178_ ;
	wire _w12177_ ;
	wire _w12176_ ;
	wire _w12175_ ;
	wire _w12174_ ;
	wire _w12173_ ;
	wire _w12172_ ;
	wire _w12171_ ;
	wire _w12170_ ;
	wire _w12169_ ;
	wire _w12168_ ;
	wire _w12167_ ;
	wire _w12166_ ;
	wire _w12165_ ;
	wire _w12164_ ;
	wire _w12163_ ;
	wire _w12162_ ;
	wire _w12161_ ;
	wire _w12160_ ;
	wire _w12159_ ;
	wire _w12158_ ;
	wire _w12157_ ;
	wire _w12156_ ;
	wire _w12155_ ;
	wire _w12154_ ;
	wire _w12153_ ;
	wire _w12152_ ;
	wire _w12151_ ;
	wire _w12150_ ;
	wire _w12149_ ;
	wire _w12148_ ;
	wire _w12147_ ;
	wire _w12146_ ;
	wire _w12145_ ;
	wire _w12144_ ;
	wire _w12143_ ;
	wire _w12142_ ;
	wire _w12141_ ;
	wire _w12140_ ;
	wire _w12139_ ;
	wire _w12138_ ;
	wire _w12137_ ;
	wire _w12136_ ;
	wire _w12135_ ;
	wire _w12134_ ;
	wire _w12133_ ;
	wire _w12132_ ;
	wire _w12131_ ;
	wire _w12130_ ;
	wire _w12129_ ;
	wire _w12128_ ;
	wire _w12127_ ;
	wire _w12126_ ;
	wire _w12125_ ;
	wire _w12124_ ;
	wire _w12123_ ;
	wire _w12122_ ;
	wire _w12121_ ;
	wire _w12120_ ;
	wire _w12119_ ;
	wire _w12118_ ;
	wire _w12117_ ;
	wire _w12116_ ;
	wire _w12115_ ;
	wire _w12114_ ;
	wire _w12113_ ;
	wire _w12112_ ;
	wire _w12111_ ;
	wire _w12110_ ;
	wire _w12109_ ;
	wire _w12108_ ;
	wire _w12107_ ;
	wire _w12106_ ;
	wire _w12105_ ;
	wire _w12104_ ;
	wire _w12103_ ;
	wire _w12102_ ;
	wire _w12101_ ;
	wire _w12100_ ;
	wire _w12099_ ;
	wire _w12098_ ;
	wire _w12097_ ;
	wire _w12096_ ;
	wire _w12095_ ;
	wire _w12094_ ;
	wire _w12093_ ;
	wire _w12092_ ;
	wire _w12091_ ;
	wire _w12090_ ;
	wire _w12089_ ;
	wire _w12088_ ;
	wire _w12087_ ;
	wire _w12086_ ;
	wire _w12085_ ;
	wire _w12084_ ;
	wire _w12083_ ;
	wire _w12082_ ;
	wire _w12081_ ;
	wire _w12080_ ;
	wire _w12079_ ;
	wire _w12078_ ;
	wire _w12077_ ;
	wire _w12076_ ;
	wire _w12075_ ;
	wire _w12074_ ;
	wire _w12073_ ;
	wire _w12072_ ;
	wire _w12071_ ;
	wire _w12070_ ;
	wire _w12069_ ;
	wire _w12068_ ;
	wire _w12067_ ;
	wire _w12066_ ;
	wire _w12065_ ;
	wire _w12064_ ;
	wire _w12063_ ;
	wire _w12062_ ;
	wire _w12061_ ;
	wire _w12060_ ;
	wire _w12059_ ;
	wire _w12058_ ;
	wire _w12057_ ;
	wire _w12056_ ;
	wire _w12055_ ;
	wire _w12054_ ;
	wire _w12053_ ;
	wire _w12052_ ;
	wire _w12051_ ;
	wire _w12050_ ;
	wire _w12049_ ;
	wire _w12048_ ;
	wire _w12047_ ;
	wire _w12046_ ;
	wire _w12045_ ;
	wire _w12044_ ;
	wire _w12043_ ;
	wire _w12042_ ;
	wire _w12041_ ;
	wire _w12040_ ;
	wire _w12039_ ;
	wire _w12038_ ;
	wire _w12037_ ;
	wire _w12036_ ;
	wire _w12035_ ;
	wire _w12034_ ;
	wire _w12033_ ;
	wire _w12032_ ;
	wire _w12031_ ;
	wire _w12030_ ;
	wire _w12029_ ;
	wire _w12028_ ;
	wire _w12027_ ;
	wire _w12026_ ;
	wire _w12025_ ;
	wire _w12024_ ;
	wire _w12023_ ;
	wire _w12022_ ;
	wire _w12021_ ;
	wire _w12020_ ;
	wire _w12019_ ;
	wire _w12018_ ;
	wire _w12017_ ;
	wire _w12016_ ;
	wire _w12015_ ;
	wire _w12014_ ;
	wire _w12013_ ;
	wire _w12012_ ;
	wire _w12011_ ;
	wire _w12010_ ;
	wire _w12009_ ;
	wire _w12008_ ;
	wire _w12007_ ;
	wire _w12006_ ;
	wire _w12005_ ;
	wire _w12004_ ;
	wire _w12003_ ;
	wire _w12002_ ;
	wire _w12001_ ;
	wire _w12000_ ;
	wire _w11999_ ;
	wire _w11998_ ;
	wire _w11997_ ;
	wire _w11996_ ;
	wire _w11995_ ;
	wire _w11994_ ;
	wire _w11993_ ;
	wire _w11992_ ;
	wire _w11991_ ;
	wire _w11990_ ;
	wire _w11989_ ;
	wire _w11988_ ;
	wire _w11987_ ;
	wire _w11986_ ;
	wire _w11985_ ;
	wire _w11984_ ;
	wire _w11983_ ;
	wire _w11982_ ;
	wire _w11981_ ;
	wire _w11980_ ;
	wire _w11979_ ;
	wire _w11978_ ;
	wire _w11977_ ;
	wire _w11976_ ;
	wire _w11975_ ;
	wire _w11974_ ;
	wire _w11973_ ;
	wire _w11972_ ;
	wire _w11971_ ;
	wire _w11970_ ;
	wire _w11969_ ;
	wire _w11968_ ;
	wire _w11967_ ;
	wire _w11966_ ;
	wire _w11965_ ;
	wire _w11964_ ;
	wire _w11963_ ;
	wire _w11962_ ;
	wire _w11961_ ;
	wire _w11960_ ;
	wire _w11959_ ;
	wire _w11958_ ;
	wire _w11957_ ;
	wire _w11956_ ;
	wire _w11955_ ;
	wire _w11954_ ;
	wire _w11953_ ;
	wire _w11952_ ;
	wire _w11951_ ;
	wire _w11950_ ;
	wire _w11949_ ;
	wire _w11948_ ;
	wire _w11947_ ;
	wire _w11946_ ;
	wire _w11945_ ;
	wire _w11944_ ;
	wire _w11943_ ;
	wire _w11942_ ;
	wire _w11941_ ;
	wire _w11940_ ;
	wire _w11939_ ;
	wire _w11938_ ;
	wire _w11937_ ;
	wire _w11936_ ;
	wire _w11935_ ;
	wire _w11934_ ;
	wire _w11933_ ;
	wire _w11932_ ;
	wire _w11931_ ;
	wire _w11930_ ;
	wire _w11929_ ;
	wire _w11928_ ;
	wire _w11927_ ;
	wire _w11926_ ;
	wire _w11925_ ;
	wire _w11924_ ;
	wire _w11923_ ;
	wire _w11922_ ;
	wire _w11921_ ;
	wire _w11920_ ;
	wire _w11919_ ;
	wire _w11918_ ;
	wire _w11917_ ;
	wire _w11916_ ;
	wire _w11915_ ;
	wire _w11914_ ;
	wire _w11913_ ;
	wire _w11912_ ;
	wire _w11911_ ;
	wire _w11910_ ;
	wire _w11909_ ;
	wire _w11908_ ;
	wire _w11907_ ;
	wire _w11906_ ;
	wire _w11905_ ;
	wire _w11904_ ;
	wire _w11903_ ;
	wire _w11902_ ;
	wire _w11901_ ;
	wire _w11900_ ;
	wire _w11899_ ;
	wire _w11898_ ;
	wire _w11897_ ;
	wire _w11896_ ;
	wire _w11895_ ;
	wire _w11894_ ;
	wire _w11893_ ;
	wire _w11892_ ;
	wire _w11891_ ;
	wire _w11890_ ;
	wire _w11889_ ;
	wire _w11888_ ;
	wire _w11887_ ;
	wire _w11886_ ;
	wire _w11885_ ;
	wire _w11884_ ;
	wire _w11883_ ;
	wire _w11882_ ;
	wire _w11881_ ;
	wire _w11880_ ;
	wire _w11879_ ;
	wire _w11878_ ;
	wire _w11877_ ;
	wire _w11876_ ;
	wire _w11875_ ;
	wire _w11874_ ;
	wire _w11873_ ;
	wire _w11872_ ;
	wire _w11871_ ;
	wire _w11870_ ;
	wire _w11869_ ;
	wire _w11868_ ;
	wire _w11867_ ;
	wire _w11866_ ;
	wire _w11865_ ;
	wire _w11864_ ;
	wire _w11863_ ;
	wire _w11862_ ;
	wire _w11861_ ;
	wire _w11860_ ;
	wire _w11859_ ;
	wire _w11858_ ;
	wire _w11857_ ;
	wire _w11856_ ;
	wire _w11855_ ;
	wire _w11854_ ;
	wire _w11853_ ;
	wire _w11852_ ;
	wire _w11851_ ;
	wire _w11850_ ;
	wire _w11849_ ;
	wire _w11848_ ;
	wire _w11847_ ;
	wire _w11846_ ;
	wire _w11845_ ;
	wire _w11844_ ;
	wire _w11843_ ;
	wire _w11842_ ;
	wire _w11841_ ;
	wire _w11840_ ;
	wire _w11839_ ;
	wire _w11838_ ;
	wire _w11837_ ;
	wire _w11836_ ;
	wire _w11835_ ;
	wire _w11834_ ;
	wire _w11833_ ;
	wire _w11832_ ;
	wire _w11831_ ;
	wire _w11830_ ;
	wire _w11829_ ;
	wire _w11828_ ;
	wire _w11827_ ;
	wire _w11826_ ;
	wire _w11825_ ;
	wire _w11824_ ;
	wire _w11823_ ;
	wire _w11822_ ;
	wire _w11821_ ;
	wire _w11820_ ;
	wire _w11819_ ;
	wire _w11818_ ;
	wire _w11817_ ;
	wire _w11816_ ;
	wire _w11815_ ;
	wire _w11814_ ;
	wire _w11813_ ;
	wire _w11812_ ;
	wire _w11811_ ;
	wire _w11810_ ;
	wire _w11809_ ;
	wire _w11808_ ;
	wire _w11807_ ;
	wire _w11806_ ;
	wire _w11805_ ;
	wire _w11804_ ;
	wire _w11803_ ;
	wire _w11802_ ;
	wire _w11801_ ;
	wire _w11800_ ;
	wire _w11799_ ;
	wire _w11798_ ;
	wire _w11797_ ;
	wire _w11796_ ;
	wire _w11795_ ;
	wire _w11794_ ;
	wire _w11793_ ;
	wire _w11792_ ;
	wire _w11791_ ;
	wire _w11790_ ;
	wire _w11789_ ;
	wire _w11788_ ;
	wire _w11787_ ;
	wire _w11786_ ;
	wire _w11785_ ;
	wire _w11784_ ;
	wire _w11783_ ;
	wire _w11782_ ;
	wire _w11781_ ;
	wire _w11780_ ;
	wire _w11779_ ;
	wire _w11778_ ;
	wire _w11777_ ;
	wire _w11776_ ;
	wire _w11775_ ;
	wire _w11774_ ;
	wire _w11773_ ;
	wire _w11772_ ;
	wire _w11771_ ;
	wire _w11770_ ;
	wire _w11769_ ;
	wire _w11768_ ;
	wire _w11767_ ;
	wire _w11766_ ;
	wire _w11765_ ;
	wire _w11764_ ;
	wire _w11763_ ;
	wire _w11762_ ;
	wire _w11761_ ;
	wire _w11760_ ;
	wire _w11759_ ;
	wire _w11758_ ;
	wire _w11757_ ;
	wire _w11756_ ;
	wire _w11755_ ;
	wire _w11754_ ;
	wire _w11753_ ;
	wire _w11752_ ;
	wire _w11751_ ;
	wire _w11750_ ;
	wire _w11749_ ;
	wire _w11748_ ;
	wire _w11747_ ;
	wire _w11746_ ;
	wire _w11745_ ;
	wire _w11744_ ;
	wire _w11743_ ;
	wire _w11742_ ;
	wire _w11741_ ;
	wire _w11740_ ;
	wire _w11739_ ;
	wire _w11738_ ;
	wire _w11737_ ;
	wire _w11736_ ;
	wire _w11735_ ;
	wire _w11734_ ;
	wire _w11733_ ;
	wire _w11732_ ;
	wire _w11731_ ;
	wire _w11730_ ;
	wire _w11729_ ;
	wire _w11728_ ;
	wire _w11727_ ;
	wire _w11726_ ;
	wire _w11725_ ;
	wire _w11724_ ;
	wire _w11723_ ;
	wire _w11722_ ;
	wire _w11721_ ;
	wire _w11720_ ;
	wire _w11719_ ;
	wire _w11718_ ;
	wire _w11717_ ;
	wire _w11716_ ;
	wire _w11715_ ;
	wire _w11714_ ;
	wire _w11713_ ;
	wire _w11712_ ;
	wire _w11711_ ;
	wire _w11710_ ;
	wire _w11709_ ;
	wire _w11708_ ;
	wire _w11707_ ;
	wire _w11706_ ;
	wire _w11705_ ;
	wire _w11704_ ;
	wire _w11703_ ;
	wire _w11702_ ;
	wire _w11701_ ;
	wire _w11700_ ;
	wire _w11699_ ;
	wire _w11698_ ;
	wire _w11697_ ;
	wire _w11696_ ;
	wire _w11695_ ;
	wire _w11694_ ;
	wire _w11693_ ;
	wire _w11692_ ;
	wire _w11691_ ;
	wire _w11690_ ;
	wire _w11689_ ;
	wire _w11688_ ;
	wire _w11687_ ;
	wire _w11686_ ;
	wire _w11685_ ;
	wire _w11684_ ;
	wire _w11683_ ;
	wire _w11682_ ;
	wire _w11681_ ;
	wire _w11680_ ;
	wire _w11679_ ;
	wire _w11678_ ;
	wire _w11677_ ;
	wire _w11676_ ;
	wire _w11675_ ;
	wire _w11674_ ;
	wire _w11673_ ;
	wire _w11672_ ;
	wire _w11671_ ;
	wire _w11670_ ;
	wire _w11669_ ;
	wire _w11668_ ;
	wire _w11667_ ;
	wire _w11666_ ;
	wire _w11665_ ;
	wire _w11664_ ;
	wire _w11663_ ;
	wire _w11662_ ;
	wire _w11661_ ;
	wire _w11660_ ;
	wire _w11659_ ;
	wire _w11658_ ;
	wire _w11657_ ;
	wire _w11656_ ;
	wire _w11655_ ;
	wire _w11654_ ;
	wire _w11653_ ;
	wire _w11652_ ;
	wire _w11651_ ;
	wire _w11650_ ;
	wire _w11649_ ;
	wire _w11648_ ;
	wire _w11647_ ;
	wire _w11646_ ;
	wire _w11645_ ;
	wire _w11644_ ;
	wire _w11643_ ;
	wire _w11642_ ;
	wire _w11641_ ;
	wire _w11640_ ;
	wire _w11639_ ;
	wire _w11638_ ;
	wire _w11637_ ;
	wire _w11636_ ;
	wire _w11635_ ;
	wire _w11634_ ;
	wire _w11633_ ;
	wire _w11632_ ;
	wire _w11631_ ;
	wire _w11630_ ;
	wire _w11629_ ;
	wire _w11628_ ;
	wire _w11627_ ;
	wire _w11626_ ;
	wire _w11625_ ;
	wire _w11624_ ;
	wire _w11623_ ;
	wire _w11622_ ;
	wire _w11621_ ;
	wire _w11620_ ;
	wire _w11619_ ;
	wire _w11618_ ;
	wire _w11617_ ;
	wire _w11616_ ;
	wire _w11615_ ;
	wire _w11614_ ;
	wire _w11613_ ;
	wire _w11612_ ;
	wire _w11611_ ;
	wire _w11610_ ;
	wire _w11609_ ;
	wire _w11608_ ;
	wire _w11607_ ;
	wire _w11606_ ;
	wire _w11605_ ;
	wire _w11604_ ;
	wire _w11603_ ;
	wire _w11602_ ;
	wire _w11601_ ;
	wire _w11600_ ;
	wire _w11599_ ;
	wire _w11598_ ;
	wire _w11597_ ;
	wire _w11596_ ;
	wire _w11595_ ;
	wire _w11594_ ;
	wire _w11593_ ;
	wire _w11592_ ;
	wire _w11591_ ;
	wire _w11590_ ;
	wire _w11589_ ;
	wire _w11588_ ;
	wire _w11587_ ;
	wire _w11586_ ;
	wire _w11585_ ;
	wire _w11584_ ;
	wire _w11583_ ;
	wire _w11582_ ;
	wire _w11581_ ;
	wire _w11580_ ;
	wire _w11579_ ;
	wire _w11578_ ;
	wire _w11577_ ;
	wire _w11576_ ;
	wire _w11575_ ;
	wire _w11574_ ;
	wire _w11573_ ;
	wire _w11572_ ;
	wire _w11571_ ;
	wire _w11570_ ;
	wire _w11569_ ;
	wire _w11568_ ;
	wire _w11567_ ;
	wire _w11566_ ;
	wire _w11565_ ;
	wire _w11564_ ;
	wire _w11563_ ;
	wire _w11562_ ;
	wire _w11561_ ;
	wire _w11560_ ;
	wire _w11559_ ;
	wire _w11558_ ;
	wire _w11557_ ;
	wire _w11556_ ;
	wire _w11555_ ;
	wire _w11554_ ;
	wire _w11553_ ;
	wire _w11552_ ;
	wire _w11551_ ;
	wire _w11550_ ;
	wire _w11549_ ;
	wire _w11548_ ;
	wire _w11547_ ;
	wire _w11546_ ;
	wire _w11545_ ;
	wire _w11544_ ;
	wire _w11543_ ;
	wire _w11542_ ;
	wire _w11541_ ;
	wire _w11540_ ;
	wire _w11539_ ;
	wire _w11538_ ;
	wire _w11537_ ;
	wire _w11536_ ;
	wire _w11535_ ;
	wire _w11534_ ;
	wire _w11533_ ;
	wire _w11532_ ;
	wire _w11531_ ;
	wire _w11530_ ;
	wire _w11529_ ;
	wire _w11528_ ;
	wire _w11527_ ;
	wire _w11526_ ;
	wire _w11525_ ;
	wire _w11524_ ;
	wire _w11523_ ;
	wire _w11522_ ;
	wire _w11521_ ;
	wire _w11520_ ;
	wire _w11519_ ;
	wire _w11518_ ;
	wire _w11517_ ;
	wire _w11516_ ;
	wire _w11515_ ;
	wire _w11514_ ;
	wire _w11513_ ;
	wire _w11512_ ;
	wire _w11511_ ;
	wire _w11510_ ;
	wire _w11509_ ;
	wire _w11508_ ;
	wire _w11507_ ;
	wire _w11506_ ;
	wire _w11505_ ;
	wire _w11504_ ;
	wire _w11503_ ;
	wire _w11502_ ;
	wire _w11501_ ;
	wire _w11500_ ;
	wire _w11499_ ;
	wire _w11498_ ;
	wire _w11497_ ;
	wire _w11496_ ;
	wire _w11495_ ;
	wire _w11494_ ;
	wire _w11493_ ;
	wire _w11492_ ;
	wire _w11491_ ;
	wire _w11490_ ;
	wire _w11489_ ;
	wire _w11488_ ;
	wire _w11487_ ;
	wire _w11486_ ;
	wire _w11485_ ;
	wire _w11484_ ;
	wire _w11483_ ;
	wire _w11482_ ;
	wire _w11481_ ;
	wire _w11480_ ;
	wire _w11479_ ;
	wire _w11478_ ;
	wire _w11477_ ;
	wire _w11476_ ;
	wire _w11475_ ;
	wire _w11474_ ;
	wire _w11473_ ;
	wire _w11472_ ;
	wire _w11471_ ;
	wire _w11470_ ;
	wire _w11469_ ;
	wire _w11468_ ;
	wire _w11467_ ;
	wire _w11466_ ;
	wire _w11465_ ;
	wire _w11464_ ;
	wire _w11463_ ;
	wire _w11462_ ;
	wire _w11461_ ;
	wire _w11460_ ;
	wire _w11459_ ;
	wire _w11458_ ;
	wire _w11457_ ;
	wire _w11456_ ;
	wire _w11455_ ;
	wire _w11454_ ;
	wire _w11453_ ;
	wire _w11452_ ;
	wire _w11451_ ;
	wire _w11450_ ;
	wire _w11449_ ;
	wire _w11448_ ;
	wire _w11447_ ;
	wire _w11446_ ;
	wire _w11445_ ;
	wire _w11444_ ;
	wire _w11443_ ;
	wire _w11442_ ;
	wire _w11441_ ;
	wire _w11440_ ;
	wire _w11439_ ;
	wire _w11438_ ;
	wire _w11437_ ;
	wire _w11436_ ;
	wire _w11435_ ;
	wire _w11434_ ;
	wire _w11433_ ;
	wire _w11432_ ;
	wire _w11431_ ;
	wire _w11430_ ;
	wire _w11429_ ;
	wire _w11428_ ;
	wire _w11427_ ;
	wire _w11426_ ;
	wire _w11425_ ;
	wire _w11424_ ;
	wire _w11423_ ;
	wire _w11422_ ;
	wire _w11421_ ;
	wire _w11420_ ;
	wire _w11419_ ;
	wire _w11418_ ;
	wire _w11417_ ;
	wire _w11416_ ;
	wire _w11415_ ;
	wire _w11414_ ;
	wire _w11413_ ;
	wire _w11412_ ;
	wire _w11411_ ;
	wire _w11410_ ;
	wire _w11409_ ;
	wire _w11408_ ;
	wire _w11407_ ;
	wire _w11406_ ;
	wire _w11405_ ;
	wire _w11404_ ;
	wire _w11403_ ;
	wire _w11402_ ;
	wire _w11401_ ;
	wire _w11400_ ;
	wire _w11399_ ;
	wire _w11398_ ;
	wire _w11397_ ;
	wire _w11396_ ;
	wire _w11395_ ;
	wire _w11394_ ;
	wire _w11393_ ;
	wire _w11392_ ;
	wire _w11391_ ;
	wire _w11390_ ;
	wire _w11389_ ;
	wire _w11388_ ;
	wire _w11387_ ;
	wire _w11386_ ;
	wire _w11385_ ;
	wire _w11384_ ;
	wire _w11383_ ;
	wire _w11382_ ;
	wire _w11381_ ;
	wire _w11380_ ;
	wire _w11379_ ;
	wire _w11378_ ;
	wire _w11377_ ;
	wire _w11376_ ;
	wire _w11375_ ;
	wire _w11374_ ;
	wire _w11373_ ;
	wire _w11372_ ;
	wire _w11371_ ;
	wire _w11370_ ;
	wire _w11369_ ;
	wire _w11368_ ;
	wire _w11367_ ;
	wire _w11366_ ;
	wire _w11365_ ;
	wire _w11364_ ;
	wire _w11363_ ;
	wire _w11362_ ;
	wire _w11361_ ;
	wire _w11360_ ;
	wire _w11359_ ;
	wire _w11358_ ;
	wire _w11357_ ;
	wire _w11356_ ;
	wire _w11355_ ;
	wire _w11354_ ;
	wire _w11353_ ;
	wire _w11352_ ;
	wire _w11351_ ;
	wire _w11350_ ;
	wire _w11349_ ;
	wire _w11348_ ;
	wire _w11347_ ;
	wire _w11346_ ;
	wire _w11345_ ;
	wire _w11344_ ;
	wire _w11343_ ;
	wire _w11342_ ;
	wire _w11341_ ;
	wire _w11340_ ;
	wire _w11339_ ;
	wire _w11338_ ;
	wire _w11337_ ;
	wire _w11336_ ;
	wire _w11335_ ;
	wire _w11334_ ;
	wire _w11333_ ;
	wire _w11332_ ;
	wire _w11331_ ;
	wire _w11330_ ;
	wire _w11329_ ;
	wire _w11328_ ;
	wire _w11327_ ;
	wire _w11326_ ;
	wire _w11325_ ;
	wire _w11324_ ;
	wire _w11323_ ;
	wire _w11322_ ;
	wire _w11321_ ;
	wire _w11320_ ;
	wire _w11319_ ;
	wire _w11318_ ;
	wire _w11317_ ;
	wire _w11316_ ;
	wire _w11315_ ;
	wire _w11314_ ;
	wire _w11313_ ;
	wire _w11312_ ;
	wire _w11311_ ;
	wire _w11310_ ;
	wire _w11309_ ;
	wire _w11308_ ;
	wire _w11307_ ;
	wire _w11306_ ;
	wire _w11305_ ;
	wire _w11304_ ;
	wire _w11303_ ;
	wire _w11302_ ;
	wire _w11301_ ;
	wire _w11300_ ;
	wire _w11299_ ;
	wire _w11298_ ;
	wire _w11297_ ;
	wire _w11296_ ;
	wire _w11295_ ;
	wire _w11294_ ;
	wire _w11293_ ;
	wire _w11292_ ;
	wire _w11291_ ;
	wire _w11290_ ;
	wire _w11289_ ;
	wire _w11288_ ;
	wire _w11287_ ;
	wire _w11286_ ;
	wire _w11285_ ;
	wire _w11284_ ;
	wire _w11283_ ;
	wire _w11282_ ;
	wire _w11281_ ;
	wire _w11280_ ;
	wire _w11279_ ;
	wire _w11278_ ;
	wire _w11277_ ;
	wire _w11276_ ;
	wire _w11275_ ;
	wire _w11274_ ;
	wire _w11273_ ;
	wire _w11272_ ;
	wire _w11271_ ;
	wire _w11270_ ;
	wire _w11269_ ;
	wire _w11268_ ;
	wire _w11267_ ;
	wire _w11266_ ;
	wire _w11265_ ;
	wire _w11264_ ;
	wire _w11263_ ;
	wire _w11262_ ;
	wire _w11261_ ;
	wire _w11260_ ;
	wire _w11259_ ;
	wire _w11258_ ;
	wire _w11257_ ;
	wire _w11256_ ;
	wire _w11255_ ;
	wire _w11254_ ;
	wire _w11253_ ;
	wire _w11252_ ;
	wire _w11251_ ;
	wire _w11250_ ;
	wire _w11249_ ;
	wire _w11248_ ;
	wire _w11247_ ;
	wire _w11246_ ;
	wire _w11245_ ;
	wire _w11244_ ;
	wire _w11243_ ;
	wire _w11242_ ;
	wire _w11241_ ;
	wire _w11240_ ;
	wire _w11239_ ;
	wire _w11238_ ;
	wire _w11237_ ;
	wire _w11236_ ;
	wire _w11235_ ;
	wire _w11234_ ;
	wire _w11233_ ;
	wire _w11232_ ;
	wire _w11231_ ;
	wire _w11230_ ;
	wire _w11229_ ;
	wire _w11228_ ;
	wire _w11227_ ;
	wire _w11226_ ;
	wire _w11225_ ;
	wire _w11224_ ;
	wire _w11223_ ;
	wire _w11222_ ;
	wire _w11221_ ;
	wire _w11220_ ;
	wire _w11219_ ;
	wire _w11218_ ;
	wire _w11217_ ;
	wire _w11216_ ;
	wire _w11215_ ;
	wire _w11214_ ;
	wire _w11213_ ;
	wire _w11212_ ;
	wire _w11211_ ;
	wire _w11210_ ;
	wire _w11209_ ;
	wire _w11208_ ;
	wire _w11207_ ;
	wire _w11206_ ;
	wire _w11205_ ;
	wire _w11204_ ;
	wire _w11203_ ;
	wire _w11202_ ;
	wire _w11201_ ;
	wire _w11200_ ;
	wire _w11199_ ;
	wire _w11198_ ;
	wire _w11197_ ;
	wire _w11196_ ;
	wire _w11195_ ;
	wire _w11194_ ;
	wire _w11193_ ;
	wire _w11192_ ;
	wire _w11191_ ;
	wire _w11190_ ;
	wire _w11189_ ;
	wire _w11188_ ;
	wire _w11187_ ;
	wire _w11186_ ;
	wire _w11185_ ;
	wire _w11184_ ;
	wire _w11183_ ;
	wire _w11182_ ;
	wire _w11181_ ;
	wire _w11180_ ;
	wire _w11179_ ;
	wire _w11178_ ;
	wire _w11177_ ;
	wire _w11176_ ;
	wire _w11175_ ;
	wire _w11174_ ;
	wire _w11173_ ;
	wire _w11172_ ;
	wire _w11171_ ;
	wire _w11170_ ;
	wire _w11169_ ;
	wire _w11168_ ;
	wire _w11167_ ;
	wire _w11166_ ;
	wire _w11165_ ;
	wire _w11164_ ;
	wire _w11163_ ;
	wire _w11162_ ;
	wire _w11161_ ;
	wire _w11160_ ;
	wire _w11159_ ;
	wire _w11158_ ;
	wire _w11157_ ;
	wire _w11156_ ;
	wire _w11155_ ;
	wire _w11154_ ;
	wire _w11153_ ;
	wire _w11152_ ;
	wire _w11151_ ;
	wire _w11150_ ;
	wire _w11149_ ;
	wire _w11148_ ;
	wire _w11147_ ;
	wire _w11146_ ;
	wire _w11145_ ;
	wire _w11144_ ;
	wire _w11143_ ;
	wire _w11142_ ;
	wire _w11141_ ;
	wire _w11140_ ;
	wire _w11139_ ;
	wire _w11138_ ;
	wire _w11137_ ;
	wire _w11136_ ;
	wire _w11135_ ;
	wire _w11134_ ;
	wire _w11133_ ;
	wire _w11132_ ;
	wire _w11131_ ;
	wire _w11130_ ;
	wire _w11129_ ;
	wire _w11128_ ;
	wire _w11127_ ;
	wire _w11126_ ;
	wire _w11125_ ;
	wire _w11124_ ;
	wire _w11123_ ;
	wire _w11122_ ;
	wire _w11121_ ;
	wire _w11120_ ;
	wire _w11119_ ;
	wire _w11118_ ;
	wire _w11117_ ;
	wire _w11116_ ;
	wire _w11115_ ;
	wire _w11114_ ;
	wire _w11113_ ;
	wire _w11112_ ;
	wire _w11111_ ;
	wire _w11110_ ;
	wire _w11109_ ;
	wire _w11108_ ;
	wire _w11107_ ;
	wire _w11106_ ;
	wire _w11105_ ;
	wire _w11104_ ;
	wire _w11103_ ;
	wire _w11102_ ;
	wire _w11101_ ;
	wire _w11100_ ;
	wire _w11099_ ;
	wire _w11098_ ;
	wire _w11097_ ;
	wire _w11096_ ;
	wire _w11095_ ;
	wire _w11094_ ;
	wire _w11093_ ;
	wire _w11092_ ;
	wire _w11091_ ;
	wire _w11090_ ;
	wire _w11089_ ;
	wire _w11088_ ;
	wire _w11087_ ;
	wire _w11086_ ;
	wire _w11085_ ;
	wire _w11084_ ;
	wire _w11083_ ;
	wire _w11082_ ;
	wire _w11081_ ;
	wire _w11080_ ;
	wire _w11079_ ;
	wire _w11078_ ;
	wire _w11077_ ;
	wire _w11076_ ;
	wire _w11075_ ;
	wire _w11074_ ;
	wire _w11073_ ;
	wire _w11072_ ;
	wire _w11071_ ;
	wire _w11070_ ;
	wire _w11069_ ;
	wire _w11068_ ;
	wire _w11067_ ;
	wire _w11066_ ;
	wire _w11065_ ;
	wire _w11064_ ;
	wire _w11063_ ;
	wire _w11062_ ;
	wire _w11061_ ;
	wire _w11060_ ;
	wire _w11059_ ;
	wire _w11058_ ;
	wire _w11057_ ;
	wire _w11056_ ;
	wire _w11055_ ;
	wire _w11054_ ;
	wire _w11053_ ;
	wire _w11052_ ;
	wire _w11051_ ;
	wire _w11050_ ;
	wire _w11049_ ;
	wire _w11048_ ;
	wire _w11047_ ;
	wire _w11046_ ;
	wire _w11045_ ;
	wire _w11044_ ;
	wire _w11043_ ;
	wire _w11042_ ;
	wire _w11041_ ;
	wire _w11040_ ;
	wire _w11039_ ;
	wire _w11038_ ;
	wire _w11037_ ;
	wire _w11036_ ;
	wire _w11035_ ;
	wire _w11034_ ;
	wire _w11033_ ;
	wire _w11032_ ;
	wire _w11031_ ;
	wire _w11030_ ;
	wire _w11029_ ;
	wire _w11028_ ;
	wire _w11027_ ;
	wire _w11026_ ;
	wire _w11025_ ;
	wire _w11024_ ;
	wire _w11023_ ;
	wire _w11022_ ;
	wire _w11021_ ;
	wire _w11020_ ;
	wire _w11019_ ;
	wire _w11018_ ;
	wire _w11017_ ;
	wire _w11016_ ;
	wire _w11015_ ;
	wire _w11014_ ;
	wire _w11013_ ;
	wire _w11012_ ;
	wire _w11011_ ;
	wire _w11010_ ;
	wire _w11009_ ;
	wire _w11008_ ;
	wire _w11007_ ;
	wire _w11006_ ;
	wire _w11005_ ;
	wire _w11004_ ;
	wire _w11003_ ;
	wire _w11002_ ;
	wire _w11001_ ;
	wire _w11000_ ;
	wire _w10999_ ;
	wire _w10998_ ;
	wire _w10997_ ;
	wire _w10996_ ;
	wire _w10995_ ;
	wire _w10994_ ;
	wire _w10993_ ;
	wire _w10992_ ;
	wire _w10991_ ;
	wire _w10990_ ;
	wire _w10989_ ;
	wire _w10988_ ;
	wire _w10987_ ;
	wire _w10986_ ;
	wire _w10985_ ;
	wire _w10984_ ;
	wire _w10983_ ;
	wire _w10982_ ;
	wire _w10981_ ;
	wire _w10980_ ;
	wire _w10979_ ;
	wire _w10978_ ;
	wire _w10977_ ;
	wire _w10976_ ;
	wire _w10975_ ;
	wire _w10974_ ;
	wire _w10973_ ;
	wire _w10972_ ;
	wire _w10971_ ;
	wire _w10970_ ;
	wire _w10969_ ;
	wire _w10968_ ;
	wire _w10967_ ;
	wire _w10966_ ;
	wire _w10965_ ;
	wire _w10964_ ;
	wire _w10963_ ;
	wire _w10962_ ;
	wire _w10961_ ;
	wire _w10960_ ;
	wire _w10959_ ;
	wire _w10958_ ;
	wire _w10957_ ;
	wire _w10956_ ;
	wire _w10955_ ;
	wire _w10954_ ;
	wire _w10953_ ;
	wire _w10952_ ;
	wire _w10951_ ;
	wire _w10950_ ;
	wire _w10949_ ;
	wire _w10948_ ;
	wire _w10947_ ;
	wire _w10946_ ;
	wire _w10945_ ;
	wire _w10944_ ;
	wire _w10943_ ;
	wire _w10942_ ;
	wire _w10941_ ;
	wire _w10940_ ;
	wire _w10939_ ;
	wire _w10938_ ;
	wire _w10937_ ;
	wire _w10936_ ;
	wire _w10935_ ;
	wire _w10934_ ;
	wire _w10933_ ;
	wire _w10932_ ;
	wire _w10931_ ;
	wire _w10930_ ;
	wire _w10929_ ;
	wire _w10928_ ;
	wire _w10927_ ;
	wire _w10926_ ;
	wire _w10925_ ;
	wire _w10924_ ;
	wire _w10923_ ;
	wire _w10922_ ;
	wire _w10921_ ;
	wire _w10920_ ;
	wire _w10919_ ;
	wire _w10918_ ;
	wire _w10917_ ;
	wire _w10916_ ;
	wire _w10915_ ;
	wire _w10914_ ;
	wire _w10913_ ;
	wire _w10912_ ;
	wire _w10911_ ;
	wire _w10910_ ;
	wire _w10909_ ;
	wire _w10908_ ;
	wire _w10907_ ;
	wire _w10906_ ;
	wire _w10905_ ;
	wire _w10904_ ;
	wire _w10903_ ;
	wire _w10902_ ;
	wire _w10901_ ;
	wire _w10900_ ;
	wire _w10899_ ;
	wire _w10898_ ;
	wire _w10897_ ;
	wire _w10896_ ;
	wire _w10895_ ;
	wire _w10894_ ;
	wire _w10893_ ;
	wire _w10892_ ;
	wire _w10891_ ;
	wire _w10890_ ;
	wire _w10889_ ;
	wire _w10888_ ;
	wire _w10887_ ;
	wire _w10886_ ;
	wire _w10885_ ;
	wire _w10884_ ;
	wire _w10883_ ;
	wire _w10882_ ;
	wire _w10881_ ;
	wire _w10880_ ;
	wire _w10879_ ;
	wire _w10878_ ;
	wire _w10877_ ;
	wire _w10876_ ;
	wire _w10875_ ;
	wire _w10874_ ;
	wire _w10873_ ;
	wire _w10872_ ;
	wire _w10871_ ;
	wire _w10870_ ;
	wire _w10869_ ;
	wire _w10868_ ;
	wire _w10867_ ;
	wire _w10866_ ;
	wire _w10865_ ;
	wire _w10864_ ;
	wire _w10863_ ;
	wire _w10862_ ;
	wire _w10861_ ;
	wire _w10860_ ;
	wire _w10859_ ;
	wire _w10858_ ;
	wire _w10857_ ;
	wire _w10856_ ;
	wire _w10855_ ;
	wire _w10854_ ;
	wire _w10853_ ;
	wire _w10852_ ;
	wire _w10851_ ;
	wire _w10850_ ;
	wire _w10849_ ;
	wire _w10848_ ;
	wire _w10847_ ;
	wire _w10846_ ;
	wire _w10845_ ;
	wire _w10844_ ;
	wire _w10843_ ;
	wire _w10842_ ;
	wire _w10841_ ;
	wire _w10840_ ;
	wire _w10839_ ;
	wire _w10838_ ;
	wire _w10837_ ;
	wire _w10836_ ;
	wire _w10835_ ;
	wire _w10834_ ;
	wire _w10833_ ;
	wire _w10832_ ;
	wire _w10831_ ;
	wire _w10830_ ;
	wire _w10829_ ;
	wire _w10828_ ;
	wire _w10827_ ;
	wire _w10826_ ;
	wire _w10825_ ;
	wire _w10824_ ;
	wire _w10823_ ;
	wire _w10822_ ;
	wire _w10821_ ;
	wire _w10820_ ;
	wire _w10819_ ;
	wire _w10818_ ;
	wire _w10817_ ;
	wire _w10816_ ;
	wire _w10815_ ;
	wire _w10814_ ;
	wire _w10813_ ;
	wire _w10812_ ;
	wire _w10811_ ;
	wire _w10810_ ;
	wire _w10809_ ;
	wire _w10808_ ;
	wire _w10807_ ;
	wire _w10806_ ;
	wire _w10805_ ;
	wire _w10804_ ;
	wire _w10803_ ;
	wire _w10802_ ;
	wire _w10801_ ;
	wire _w10800_ ;
	wire _w10799_ ;
	wire _w10798_ ;
	wire _w10797_ ;
	wire _w10796_ ;
	wire _w10795_ ;
	wire _w10794_ ;
	wire _w10793_ ;
	wire _w10792_ ;
	wire _w10791_ ;
	wire _w10790_ ;
	wire _w10789_ ;
	wire _w10788_ ;
	wire _w10787_ ;
	wire _w10786_ ;
	wire _w10785_ ;
	wire _w10784_ ;
	wire _w10783_ ;
	wire _w10782_ ;
	wire _w10781_ ;
	wire _w10780_ ;
	wire _w10779_ ;
	wire _w10778_ ;
	wire _w10777_ ;
	wire _w10776_ ;
	wire _w10775_ ;
	wire _w10774_ ;
	wire _w10773_ ;
	wire _w10772_ ;
	wire _w10771_ ;
	wire _w10770_ ;
	wire _w10769_ ;
	wire _w10768_ ;
	wire _w10767_ ;
	wire _w10766_ ;
	wire _w10765_ ;
	wire _w10764_ ;
	wire _w10763_ ;
	wire _w10762_ ;
	wire _w10761_ ;
	wire _w10760_ ;
	wire _w10759_ ;
	wire _w10758_ ;
	wire _w10757_ ;
	wire _w10756_ ;
	wire _w10755_ ;
	wire _w10754_ ;
	wire _w10753_ ;
	wire _w10752_ ;
	wire _w10751_ ;
	wire _w10750_ ;
	wire _w10749_ ;
	wire _w10748_ ;
	wire _w10747_ ;
	wire _w10746_ ;
	wire _w10745_ ;
	wire _w10744_ ;
	wire _w10743_ ;
	wire _w10742_ ;
	wire _w10741_ ;
	wire _w10740_ ;
	wire _w10739_ ;
	wire _w10738_ ;
	wire _w10737_ ;
	wire _w10736_ ;
	wire _w10735_ ;
	wire _w10734_ ;
	wire _w10733_ ;
	wire _w10732_ ;
	wire _w10731_ ;
	wire _w10730_ ;
	wire _w10729_ ;
	wire _w10728_ ;
	wire _w10727_ ;
	wire _w10726_ ;
	wire _w10725_ ;
	wire _w10724_ ;
	wire _w10723_ ;
	wire _w10722_ ;
	wire _w10721_ ;
	wire _w10720_ ;
	wire _w10719_ ;
	wire _w10718_ ;
	wire _w10717_ ;
	wire _w10716_ ;
	wire _w10715_ ;
	wire _w10714_ ;
	wire _w10713_ ;
	wire _w10712_ ;
	wire _w10711_ ;
	wire _w10710_ ;
	wire _w10709_ ;
	wire _w10708_ ;
	wire _w10707_ ;
	wire _w10706_ ;
	wire _w10705_ ;
	wire _w10704_ ;
	wire _w10703_ ;
	wire _w10702_ ;
	wire _w10701_ ;
	wire _w10700_ ;
	wire _w10699_ ;
	wire _w10698_ ;
	wire _w10697_ ;
	wire _w10696_ ;
	wire _w10695_ ;
	wire _w10694_ ;
	wire _w10693_ ;
	wire _w10692_ ;
	wire _w10691_ ;
	wire _w10690_ ;
	wire _w10689_ ;
	wire _w10688_ ;
	wire _w10687_ ;
	wire _w10686_ ;
	wire _w10685_ ;
	wire _w10684_ ;
	wire _w10683_ ;
	wire _w10682_ ;
	wire _w10681_ ;
	wire _w10680_ ;
	wire _w10679_ ;
	wire _w10678_ ;
	wire _w10677_ ;
	wire _w10676_ ;
	wire _w10675_ ;
	wire _w10674_ ;
	wire _w10673_ ;
	wire _w10672_ ;
	wire _w10671_ ;
	wire _w10670_ ;
	wire _w10669_ ;
	wire _w10668_ ;
	wire _w10667_ ;
	wire _w10666_ ;
	wire _w10665_ ;
	wire _w10664_ ;
	wire _w10663_ ;
	wire _w10662_ ;
	wire _w10661_ ;
	wire _w10660_ ;
	wire _w10659_ ;
	wire _w10658_ ;
	wire _w10657_ ;
	wire _w10656_ ;
	wire _w10655_ ;
	wire _w10654_ ;
	wire _w10653_ ;
	wire _w10652_ ;
	wire _w10651_ ;
	wire _w10650_ ;
	wire _w10649_ ;
	wire _w10648_ ;
	wire _w10647_ ;
	wire _w10646_ ;
	wire _w10645_ ;
	wire _w10644_ ;
	wire _w10643_ ;
	wire _w10642_ ;
	wire _w10641_ ;
	wire _w10640_ ;
	wire _w10639_ ;
	wire _w10638_ ;
	wire _w10637_ ;
	wire _w10636_ ;
	wire _w10635_ ;
	wire _w10634_ ;
	wire _w10633_ ;
	wire _w10632_ ;
	wire _w10631_ ;
	wire _w10630_ ;
	wire _w10629_ ;
	wire _w10628_ ;
	wire _w10627_ ;
	wire _w10626_ ;
	wire _w10625_ ;
	wire _w10624_ ;
	wire _w10623_ ;
	wire _w10622_ ;
	wire _w10621_ ;
	wire _w10620_ ;
	wire _w10619_ ;
	wire _w10618_ ;
	wire _w10617_ ;
	wire _w10616_ ;
	wire _w10615_ ;
	wire _w10614_ ;
	wire _w10613_ ;
	wire _w10612_ ;
	wire _w10611_ ;
	wire _w10610_ ;
	wire _w10609_ ;
	wire _w10608_ ;
	wire _w10607_ ;
	wire _w10606_ ;
	wire _w10605_ ;
	wire _w10604_ ;
	wire _w10603_ ;
	wire _w10602_ ;
	wire _w10601_ ;
	wire _w10600_ ;
	wire _w10599_ ;
	wire _w10598_ ;
	wire _w10597_ ;
	wire _w10596_ ;
	wire _w10595_ ;
	wire _w10594_ ;
	wire _w10593_ ;
	wire _w10592_ ;
	wire _w10591_ ;
	wire _w10590_ ;
	wire _w10589_ ;
	wire _w10588_ ;
	wire _w10587_ ;
	wire _w10586_ ;
	wire _w10585_ ;
	wire _w10584_ ;
	wire _w10583_ ;
	wire _w10582_ ;
	wire _w10581_ ;
	wire _w10580_ ;
	wire _w10579_ ;
	wire _w10578_ ;
	wire _w10577_ ;
	wire _w10576_ ;
	wire _w10575_ ;
	wire _w10574_ ;
	wire _w10573_ ;
	wire _w10572_ ;
	wire _w10571_ ;
	wire _w10570_ ;
	wire _w10569_ ;
	wire _w10568_ ;
	wire _w10567_ ;
	wire _w10566_ ;
	wire _w10565_ ;
	wire _w10564_ ;
	wire _w10563_ ;
	wire _w10562_ ;
	wire _w10561_ ;
	wire _w10560_ ;
	wire _w10559_ ;
	wire _w10558_ ;
	wire _w10557_ ;
	wire _w10556_ ;
	wire _w10555_ ;
	wire _w10554_ ;
	wire _w10553_ ;
	wire _w10552_ ;
	wire _w10551_ ;
	wire _w10550_ ;
	wire _w10549_ ;
	wire _w10548_ ;
	wire _w10547_ ;
	wire _w10546_ ;
	wire _w10545_ ;
	wire _w10544_ ;
	wire _w10543_ ;
	wire _w10542_ ;
	wire _w10541_ ;
	wire _w10540_ ;
	wire _w10539_ ;
	wire _w10538_ ;
	wire _w10537_ ;
	wire _w10536_ ;
	wire _w10535_ ;
	wire _w10534_ ;
	wire _w10533_ ;
	wire _w10532_ ;
	wire _w10531_ ;
	wire _w10530_ ;
	wire _w10529_ ;
	wire _w10528_ ;
	wire _w10527_ ;
	wire _w10526_ ;
	wire _w10525_ ;
	wire _w10524_ ;
	wire _w10523_ ;
	wire _w10522_ ;
	wire _w10521_ ;
	wire _w10520_ ;
	wire _w10519_ ;
	wire _w10518_ ;
	wire _w10517_ ;
	wire _w10516_ ;
	wire _w10515_ ;
	wire _w10514_ ;
	wire _w10513_ ;
	wire _w10512_ ;
	wire _w10511_ ;
	wire _w10510_ ;
	wire _w10509_ ;
	wire _w10508_ ;
	wire _w10507_ ;
	wire _w10506_ ;
	wire _w10505_ ;
	wire _w10504_ ;
	wire _w10503_ ;
	wire _w10502_ ;
	wire _w10501_ ;
	wire _w10500_ ;
	wire _w10499_ ;
	wire _w10498_ ;
	wire _w10497_ ;
	wire _w10496_ ;
	wire _w10495_ ;
	wire _w10494_ ;
	wire _w10493_ ;
	wire _w10492_ ;
	wire _w10491_ ;
	wire _w10490_ ;
	wire _w10489_ ;
	wire _w10488_ ;
	wire _w10487_ ;
	wire _w10486_ ;
	wire _w10485_ ;
	wire _w10484_ ;
	wire _w10483_ ;
	wire _w10482_ ;
	wire _w10481_ ;
	wire _w10480_ ;
	wire _w10479_ ;
	wire _w10478_ ;
	wire _w10477_ ;
	wire _w10476_ ;
	wire _w10475_ ;
	wire _w10474_ ;
	wire _w10473_ ;
	wire _w10472_ ;
	wire _w10471_ ;
	wire _w10470_ ;
	wire _w10469_ ;
	wire _w10468_ ;
	wire _w10467_ ;
	wire _w10466_ ;
	wire _w10465_ ;
	wire _w10464_ ;
	wire _w10463_ ;
	wire _w10462_ ;
	wire _w10461_ ;
	wire _w10460_ ;
	wire _w10459_ ;
	wire _w10458_ ;
	wire _w10457_ ;
	wire _w10456_ ;
	wire _w10455_ ;
	wire _w10454_ ;
	wire _w10453_ ;
	wire _w10452_ ;
	wire _w10451_ ;
	wire _w10450_ ;
	wire _w10449_ ;
	wire _w10448_ ;
	wire _w10447_ ;
	wire _w10446_ ;
	wire _w10445_ ;
	wire _w10444_ ;
	wire _w10443_ ;
	wire _w10442_ ;
	wire _w10441_ ;
	wire _w10440_ ;
	wire _w10439_ ;
	wire _w10438_ ;
	wire _w10437_ ;
	wire _w10436_ ;
	wire _w10435_ ;
	wire _w10434_ ;
	wire _w10433_ ;
	wire _w10432_ ;
	wire _w10431_ ;
	wire _w10430_ ;
	wire _w10429_ ;
	wire _w10428_ ;
	wire _w10427_ ;
	wire _w10426_ ;
	wire _w10425_ ;
	wire _w10424_ ;
	wire _w10423_ ;
	wire _w10422_ ;
	wire _w10421_ ;
	wire _w10420_ ;
	wire _w10419_ ;
	wire _w10418_ ;
	wire _w10417_ ;
	wire _w10416_ ;
	wire _w10415_ ;
	wire _w10414_ ;
	wire _w10413_ ;
	wire _w10412_ ;
	wire _w10411_ ;
	wire _w10410_ ;
	wire _w10409_ ;
	wire _w10408_ ;
	wire _w10407_ ;
	wire _w10406_ ;
	wire _w10405_ ;
	wire _w10404_ ;
	wire _w10403_ ;
	wire _w10402_ ;
	wire _w10401_ ;
	wire _w10400_ ;
	wire _w10399_ ;
	wire _w10398_ ;
	wire _w10397_ ;
	wire _w10396_ ;
	wire _w10395_ ;
	wire _w10394_ ;
	wire _w10393_ ;
	wire _w10392_ ;
	wire _w10391_ ;
	wire _w10390_ ;
	wire _w10389_ ;
	wire _w10388_ ;
	wire _w10387_ ;
	wire _w10386_ ;
	wire _w10385_ ;
	wire _w10384_ ;
	wire _w10383_ ;
	wire _w10382_ ;
	wire _w10381_ ;
	wire _w10380_ ;
	wire _w10379_ ;
	wire _w10378_ ;
	wire _w10377_ ;
	wire _w10376_ ;
	wire _w10375_ ;
	wire _w10374_ ;
	wire _w10373_ ;
	wire _w10372_ ;
	wire _w10371_ ;
	wire _w10370_ ;
	wire _w10369_ ;
	wire _w10368_ ;
	wire _w10367_ ;
	wire _w10366_ ;
	wire _w10365_ ;
	wire _w10364_ ;
	wire _w10363_ ;
	wire _w10362_ ;
	wire _w10361_ ;
	wire _w10360_ ;
	wire _w10359_ ;
	wire _w10358_ ;
	wire _w10357_ ;
	wire _w10356_ ;
	wire _w10355_ ;
	wire _w10354_ ;
	wire _w10353_ ;
	wire _w10352_ ;
	wire _w10351_ ;
	wire _w10350_ ;
	wire _w10349_ ;
	wire _w10348_ ;
	wire _w10347_ ;
	wire _w10346_ ;
	wire _w10345_ ;
	wire _w10344_ ;
	wire _w10343_ ;
	wire _w10342_ ;
	wire _w10341_ ;
	wire _w10340_ ;
	wire _w10339_ ;
	wire _w10338_ ;
	wire _w10337_ ;
	wire _w10336_ ;
	wire _w10335_ ;
	wire _w10334_ ;
	wire _w10333_ ;
	wire _w10332_ ;
	wire _w10331_ ;
	wire _w10330_ ;
	wire _w10329_ ;
	wire _w10328_ ;
	wire _w10327_ ;
	wire _w10326_ ;
	wire _w10325_ ;
	wire _w10324_ ;
	wire _w10323_ ;
	wire _w10322_ ;
	wire _w10321_ ;
	wire _w10320_ ;
	wire _w10319_ ;
	wire _w10318_ ;
	wire _w10317_ ;
	wire _w10316_ ;
	wire _w10315_ ;
	wire _w10314_ ;
	wire _w10313_ ;
	wire _w10312_ ;
	wire _w10311_ ;
	wire _w10310_ ;
	wire _w10309_ ;
	wire _w10308_ ;
	wire _w10307_ ;
	wire _w5120_ ;
	wire _w5119_ ;
	wire _w5118_ ;
	wire _w5117_ ;
	wire _w5116_ ;
	wire _w5115_ ;
	wire _w5114_ ;
	wire _w5113_ ;
	wire _w5112_ ;
	wire _w5111_ ;
	wire _w5110_ ;
	wire _w5109_ ;
	wire _w5108_ ;
	wire _w5107_ ;
	wire _w5106_ ;
	wire _w5105_ ;
	wire _w5104_ ;
	wire _w5103_ ;
	wire _w5102_ ;
	wire _w5101_ ;
	wire _w5100_ ;
	wire _w5099_ ;
	wire _w5098_ ;
	wire _w5097_ ;
	wire _w5096_ ;
	wire _w5095_ ;
	wire _w5094_ ;
	wire _w5093_ ;
	wire _w5092_ ;
	wire _w5091_ ;
	wire _w5090_ ;
	wire _w5089_ ;
	wire _w5088_ ;
	wire _w5087_ ;
	wire _w5086_ ;
	wire _w5085_ ;
	wire _w5084_ ;
	wire _w5083_ ;
	wire _w5082_ ;
	wire _w5081_ ;
	wire _w5080_ ;
	wire _w5079_ ;
	wire _w5078_ ;
	wire _w5077_ ;
	wire _w5076_ ;
	wire _w5075_ ;
	wire _w5074_ ;
	wire _w5073_ ;
	wire _w5072_ ;
	wire _w5071_ ;
	wire _w5070_ ;
	wire _w5069_ ;
	wire _w5068_ ;
	wire _w5067_ ;
	wire _w5066_ ;
	wire _w5065_ ;
	wire _w5064_ ;
	wire _w5063_ ;
	wire _w5062_ ;
	wire _w5061_ ;
	wire _w5060_ ;
	wire _w5059_ ;
	wire _w5058_ ;
	wire _w5057_ ;
	wire _w5056_ ;
	wire _w5055_ ;
	wire _w5054_ ;
	wire _w5053_ ;
	wire _w5052_ ;
	wire _w5051_ ;
	wire _w5050_ ;
	wire _w5049_ ;
	wire _w5048_ ;
	wire _w5047_ ;
	wire _w5046_ ;
	wire _w5045_ ;
	wire _w5044_ ;
	wire _w5043_ ;
	wire _w5042_ ;
	wire _w5041_ ;
	wire _w5040_ ;
	wire _w5039_ ;
	wire _w5038_ ;
	wire _w5037_ ;
	wire _w5036_ ;
	wire _w5035_ ;
	wire _w5034_ ;
	wire _w5033_ ;
	wire _w5032_ ;
	wire _w5031_ ;
	wire _w5030_ ;
	wire _w5029_ ;
	wire _w5028_ ;
	wire _w5027_ ;
	wire _w5026_ ;
	wire _w5025_ ;
	wire _w5024_ ;
	wire _w5023_ ;
	wire _w5022_ ;
	wire _w5021_ ;
	wire _w5020_ ;
	wire _w5019_ ;
	wire _w5018_ ;
	wire _w5017_ ;
	wire _w5016_ ;
	wire _w5015_ ;
	wire _w5014_ ;
	wire _w5013_ ;
	wire _w5012_ ;
	wire _w5011_ ;
	wire _w5010_ ;
	wire _w5009_ ;
	wire _w5008_ ;
	wire _w5007_ ;
	wire _w5006_ ;
	wire _w5005_ ;
	wire _w5004_ ;
	wire _w5003_ ;
	wire _w5002_ ;
	wire _w5001_ ;
	wire _w5000_ ;
	wire _w4999_ ;
	wire _w4998_ ;
	wire _w4997_ ;
	wire _w4996_ ;
	wire _w4995_ ;
	wire _w4994_ ;
	wire _w4993_ ;
	wire _w4992_ ;
	wire _w4991_ ;
	wire _w4990_ ;
	wire _w4989_ ;
	wire _w4988_ ;
	wire _w4987_ ;
	wire _w4986_ ;
	wire _w4985_ ;
	wire _w4984_ ;
	wire _w4983_ ;
	wire _w4982_ ;
	wire _w4981_ ;
	wire _w4980_ ;
	wire _w4979_ ;
	wire _w4978_ ;
	wire _w4977_ ;
	wire _w4976_ ;
	wire _w4975_ ;
	wire _w4974_ ;
	wire _w4973_ ;
	wire _w4972_ ;
	wire _w4971_ ;
	wire _w4970_ ;
	wire _w4969_ ;
	wire _w4968_ ;
	wire _w4967_ ;
	wire _w4966_ ;
	wire _w4965_ ;
	wire _w4964_ ;
	wire _w4963_ ;
	wire _w4962_ ;
	wire _w4961_ ;
	wire _w4960_ ;
	wire _w4959_ ;
	wire _w4958_ ;
	wire _w4957_ ;
	wire _w4956_ ;
	wire _w4955_ ;
	wire _w4954_ ;
	wire _w4953_ ;
	wire _w4952_ ;
	wire _w4951_ ;
	wire _w4950_ ;
	wire _w4949_ ;
	wire _w4948_ ;
	wire _w4947_ ;
	wire _w4946_ ;
	wire _w4945_ ;
	wire _w4944_ ;
	wire _w4943_ ;
	wire _w4942_ ;
	wire _w4941_ ;
	wire _w4940_ ;
	wire _w4939_ ;
	wire _w4938_ ;
	wire _w4937_ ;
	wire _w4936_ ;
	wire _w4935_ ;
	wire _w4934_ ;
	wire _w4933_ ;
	wire _w4932_ ;
	wire _w4931_ ;
	wire _w4930_ ;
	wire _w4929_ ;
	wire _w4928_ ;
	wire _w4927_ ;
	wire _w4926_ ;
	wire _w4925_ ;
	wire _w4924_ ;
	wire _w4923_ ;
	wire _w4922_ ;
	wire _w4921_ ;
	wire _w4920_ ;
	wire _w4919_ ;
	wire _w4918_ ;
	wire _w4917_ ;
	wire _w4916_ ;
	wire _w4915_ ;
	wire _w4914_ ;
	wire _w4913_ ;
	wire _w4912_ ;
	wire _w4911_ ;
	wire _w4910_ ;
	wire _w4909_ ;
	wire _w4908_ ;
	wire _w4907_ ;
	wire _w4906_ ;
	wire _w4905_ ;
	wire _w4904_ ;
	wire _w4903_ ;
	wire _w4902_ ;
	wire _w4901_ ;
	wire _w4900_ ;
	wire _w4899_ ;
	wire _w4898_ ;
	wire _w4897_ ;
	wire _w4896_ ;
	wire _w4895_ ;
	wire _w4894_ ;
	wire _w4893_ ;
	wire _w4892_ ;
	wire _w4891_ ;
	wire _w4890_ ;
	wire _w4889_ ;
	wire _w4888_ ;
	wire _w4887_ ;
	wire _w4886_ ;
	wire _w4885_ ;
	wire _w4884_ ;
	wire _w4883_ ;
	wire _w4882_ ;
	wire _w4881_ ;
	wire _w4880_ ;
	wire _w4879_ ;
	wire _w4878_ ;
	wire _w4877_ ;
	wire _w4876_ ;
	wire _w4875_ ;
	wire _w4874_ ;
	wire _w4873_ ;
	wire _w4872_ ;
	wire _w4871_ ;
	wire _w4870_ ;
	wire _w4869_ ;
	wire _w4868_ ;
	wire _w4867_ ;
	wire _w4866_ ;
	wire _w4865_ ;
	wire _w4864_ ;
	wire _w4863_ ;
	wire _w4862_ ;
	wire _w4861_ ;
	wire _w4860_ ;
	wire _w4859_ ;
	wire _w4858_ ;
	wire _w4857_ ;
	wire _w4856_ ;
	wire _w4855_ ;
	wire _w4854_ ;
	wire _w4853_ ;
	wire _w4852_ ;
	wire _w4851_ ;
	wire _w4850_ ;
	wire _w4849_ ;
	wire _w4848_ ;
	wire _w4847_ ;
	wire _w4846_ ;
	wire _w4845_ ;
	wire _w4844_ ;
	wire _w4843_ ;
	wire _w4842_ ;
	wire _w4841_ ;
	wire _w4840_ ;
	wire _w4839_ ;
	wire _w4838_ ;
	wire _w4837_ ;
	wire _w4836_ ;
	wire _w4835_ ;
	wire _w4834_ ;
	wire _w4833_ ;
	wire _w4832_ ;
	wire _w4831_ ;
	wire _w4830_ ;
	wire _w4829_ ;
	wire _w4828_ ;
	wire _w4827_ ;
	wire _w4826_ ;
	wire _w4825_ ;
	wire _w4824_ ;
	wire _w4823_ ;
	wire _w4822_ ;
	wire _w4821_ ;
	wire _w4820_ ;
	wire _w4819_ ;
	wire _w4818_ ;
	wire _w4817_ ;
	wire _w4816_ ;
	wire _w4815_ ;
	wire _w4814_ ;
	wire _w4813_ ;
	wire _w4812_ ;
	wire _w4811_ ;
	wire _w4810_ ;
	wire _w4809_ ;
	wire _w4808_ ;
	wire _w4807_ ;
	wire _w4806_ ;
	wire _w4805_ ;
	wire _w4804_ ;
	wire _w4803_ ;
	wire _w4802_ ;
	wire _w4801_ ;
	wire _w4800_ ;
	wire _w4799_ ;
	wire _w4798_ ;
	wire _w4797_ ;
	wire _w4796_ ;
	wire _w4795_ ;
	wire _w4794_ ;
	wire _w4793_ ;
	wire _w4792_ ;
	wire _w4791_ ;
	wire _w4790_ ;
	wire _w4789_ ;
	wire _w4788_ ;
	wire _w4787_ ;
	wire _w4786_ ;
	wire _w4785_ ;
	wire _w4784_ ;
	wire _w4783_ ;
	wire _w4782_ ;
	wire _w4781_ ;
	wire _w4780_ ;
	wire _w4779_ ;
	wire _w4778_ ;
	wire _w4777_ ;
	wire _w4776_ ;
	wire _w4775_ ;
	wire _w4774_ ;
	wire _w4773_ ;
	wire _w4772_ ;
	wire _w4771_ ;
	wire _w4770_ ;
	wire _w4769_ ;
	wire _w4768_ ;
	wire _w4767_ ;
	wire _w4766_ ;
	wire _w4765_ ;
	wire _w4764_ ;
	wire _w4763_ ;
	wire _w4762_ ;
	wire _w4761_ ;
	wire _w4760_ ;
	wire _w4759_ ;
	wire _w4758_ ;
	wire _w4757_ ;
	wire _w4756_ ;
	wire _w4755_ ;
	wire _w4754_ ;
	wire _w4753_ ;
	wire _w4752_ ;
	wire _w4751_ ;
	wire _w4750_ ;
	wire _w4749_ ;
	wire _w4748_ ;
	wire _w4747_ ;
	wire _w4746_ ;
	wire _w4745_ ;
	wire _w4744_ ;
	wire _w4743_ ;
	wire _w4742_ ;
	wire _w4741_ ;
	wire _w4740_ ;
	wire _w4739_ ;
	wire _w4738_ ;
	wire _w4737_ ;
	wire _w4736_ ;
	wire _w4735_ ;
	wire _w4734_ ;
	wire _w4733_ ;
	wire _w4732_ ;
	wire _w4731_ ;
	wire _w4730_ ;
	wire _w4729_ ;
	wire _w4728_ ;
	wire _w4727_ ;
	wire _w4726_ ;
	wire _w4725_ ;
	wire _w4724_ ;
	wire _w4723_ ;
	wire _w4722_ ;
	wire _w4721_ ;
	wire _w4720_ ;
	wire _w4719_ ;
	wire _w4718_ ;
	wire _w4717_ ;
	wire _w4716_ ;
	wire _w4715_ ;
	wire _w4714_ ;
	wire _w4713_ ;
	wire _w4712_ ;
	wire _w4711_ ;
	wire _w4710_ ;
	wire _w4709_ ;
	wire _w4708_ ;
	wire _w4707_ ;
	wire _w4706_ ;
	wire _w4705_ ;
	wire _w4704_ ;
	wire _w4703_ ;
	wire _w4702_ ;
	wire _w4701_ ;
	wire _w4700_ ;
	wire _w4699_ ;
	wire _w4698_ ;
	wire _w4697_ ;
	wire _w4696_ ;
	wire _w4695_ ;
	wire _w4694_ ;
	wire _w4693_ ;
	wire _w4692_ ;
	wire _w4691_ ;
	wire _w4690_ ;
	wire _w4689_ ;
	wire _w4688_ ;
	wire _w4687_ ;
	wire _w4686_ ;
	wire _w4685_ ;
	wire _w4684_ ;
	wire _w4683_ ;
	wire _w4682_ ;
	wire _w4681_ ;
	wire _w4680_ ;
	wire _w4679_ ;
	wire _w4678_ ;
	wire _w4677_ ;
	wire _w4676_ ;
	wire _w4675_ ;
	wire _w4674_ ;
	wire _w4673_ ;
	wire _w4672_ ;
	wire _w4671_ ;
	wire _w4670_ ;
	wire _w4669_ ;
	wire _w4668_ ;
	wire _w4667_ ;
	wire _w4666_ ;
	wire _w4665_ ;
	wire _w4664_ ;
	wire _w4663_ ;
	wire _w4662_ ;
	wire _w4661_ ;
	wire _w4660_ ;
	wire _w4659_ ;
	wire _w4658_ ;
	wire _w4657_ ;
	wire _w4656_ ;
	wire _w4655_ ;
	wire _w4654_ ;
	wire _w4653_ ;
	wire _w4652_ ;
	wire _w4651_ ;
	wire _w4650_ ;
	wire _w4649_ ;
	wire _w4648_ ;
	wire _w4647_ ;
	wire _w4646_ ;
	wire _w4645_ ;
	wire _w4644_ ;
	wire _w4643_ ;
	wire _w4642_ ;
	wire _w4641_ ;
	wire _w4640_ ;
	wire _w4639_ ;
	wire _w4638_ ;
	wire _w4637_ ;
	wire _w4636_ ;
	wire _w4635_ ;
	wire _w4634_ ;
	wire _w4633_ ;
	wire _w4632_ ;
	wire _w4631_ ;
	wire _w4630_ ;
	wire _w4629_ ;
	wire _w4628_ ;
	wire _w4627_ ;
	wire _w4626_ ;
	wire _w4625_ ;
	wire _w4624_ ;
	wire _w4623_ ;
	wire _w4622_ ;
	wire _w4621_ ;
	wire _w4620_ ;
	wire _w4619_ ;
	wire _w4618_ ;
	wire _w4617_ ;
	wire _w4616_ ;
	wire _w4615_ ;
	wire _w4614_ ;
	wire _w4613_ ;
	wire _w4612_ ;
	wire _w4611_ ;
	wire _w4610_ ;
	wire _w4609_ ;
	wire _w4608_ ;
	wire _w4607_ ;
	wire _w4606_ ;
	wire _w4605_ ;
	wire _w4604_ ;
	wire _w4603_ ;
	wire _w4602_ ;
	wire _w4601_ ;
	wire _w4600_ ;
	wire _w4599_ ;
	wire _w4598_ ;
	wire _w4597_ ;
	wire _w4596_ ;
	wire _w4595_ ;
	wire _w4594_ ;
	wire _w4593_ ;
	wire _w4592_ ;
	wire _w4591_ ;
	wire _w4590_ ;
	wire _w4589_ ;
	wire _w4588_ ;
	wire _w4587_ ;
	wire _w4586_ ;
	wire _w4585_ ;
	wire _w4584_ ;
	wire _w4583_ ;
	wire _w4582_ ;
	wire _w4581_ ;
	wire _w4580_ ;
	wire _w4579_ ;
	wire _w4578_ ;
	wire _w4577_ ;
	wire _w4576_ ;
	wire _w4575_ ;
	wire _w4574_ ;
	wire _w4573_ ;
	wire _w4572_ ;
	wire _w4571_ ;
	wire _w4570_ ;
	wire _w4569_ ;
	wire _w4568_ ;
	wire _w4567_ ;
	wire _w4566_ ;
	wire _w4565_ ;
	wire _w4564_ ;
	wire _w4563_ ;
	wire _w4562_ ;
	wire _w4561_ ;
	wire _w4560_ ;
	wire _w4559_ ;
	wire _w4558_ ;
	wire _w4557_ ;
	wire _w4556_ ;
	wire _w4555_ ;
	wire _w4554_ ;
	wire _w4553_ ;
	wire _w4552_ ;
	wire _w4551_ ;
	wire _w4550_ ;
	wire _w4549_ ;
	wire _w4548_ ;
	wire _w4547_ ;
	wire _w4546_ ;
	wire _w4545_ ;
	wire _w4544_ ;
	wire _w4543_ ;
	wire _w4542_ ;
	wire _w4541_ ;
	wire _w4540_ ;
	wire _w4539_ ;
	wire _w4538_ ;
	wire _w4537_ ;
	wire _w4536_ ;
	wire _w4535_ ;
	wire _w4534_ ;
	wire _w4533_ ;
	wire _w4532_ ;
	wire _w4531_ ;
	wire _w4530_ ;
	wire _w4529_ ;
	wire _w4528_ ;
	wire _w4527_ ;
	wire _w4526_ ;
	wire _w4525_ ;
	wire _w4524_ ;
	wire _w4523_ ;
	wire _w4522_ ;
	wire _w4521_ ;
	wire _w4520_ ;
	wire _w4519_ ;
	wire _w4518_ ;
	wire _w4517_ ;
	wire _w4516_ ;
	wire _w4515_ ;
	wire _w4514_ ;
	wire _w4513_ ;
	wire _w4512_ ;
	wire _w4511_ ;
	wire _w4510_ ;
	wire _w4509_ ;
	wire _w4508_ ;
	wire _w4507_ ;
	wire _w4506_ ;
	wire _w4505_ ;
	wire _w4504_ ;
	wire _w4503_ ;
	wire _w4502_ ;
	wire _w4501_ ;
	wire _w4500_ ;
	wire _w4499_ ;
	wire _w4498_ ;
	wire _w4497_ ;
	wire _w4496_ ;
	wire _w4495_ ;
	wire _w4494_ ;
	wire _w4493_ ;
	wire _w4492_ ;
	wire _w4491_ ;
	wire _w4490_ ;
	wire _w4489_ ;
	wire _w4488_ ;
	wire _w4487_ ;
	wire _w4486_ ;
	wire _w4485_ ;
	wire _w4484_ ;
	wire _w4483_ ;
	wire _w4482_ ;
	wire _w4481_ ;
	wire _w4480_ ;
	wire _w4479_ ;
	wire _w4478_ ;
	wire _w4477_ ;
	wire _w4476_ ;
	wire _w4475_ ;
	wire _w4474_ ;
	wire _w4473_ ;
	wire _w4472_ ;
	wire _w4471_ ;
	wire _w4470_ ;
	wire _w4469_ ;
	wire _w4468_ ;
	wire _w4467_ ;
	wire _w4466_ ;
	wire _w4465_ ;
	wire _w4464_ ;
	wire _w4463_ ;
	wire _w4462_ ;
	wire _w4461_ ;
	wire _w4460_ ;
	wire _w4459_ ;
	wire _w4458_ ;
	wire _w4457_ ;
	wire _w4456_ ;
	wire _w4455_ ;
	wire _w4454_ ;
	wire _w4453_ ;
	wire _w4452_ ;
	wire _w4451_ ;
	wire _w4450_ ;
	wire _w4449_ ;
	wire _w4448_ ;
	wire _w4447_ ;
	wire _w4446_ ;
	wire _w4445_ ;
	wire _w4444_ ;
	wire _w4443_ ;
	wire _w4442_ ;
	wire _w4441_ ;
	wire _w4440_ ;
	wire _w4439_ ;
	wire _w4438_ ;
	wire _w4437_ ;
	wire _w4436_ ;
	wire _w4435_ ;
	wire _w4434_ ;
	wire _w4433_ ;
	wire _w4432_ ;
	wire _w4431_ ;
	wire _w4430_ ;
	wire _w4429_ ;
	wire _w4428_ ;
	wire _w4427_ ;
	wire _w4426_ ;
	wire _w4425_ ;
	wire _w4424_ ;
	wire _w4423_ ;
	wire _w4422_ ;
	wire _w4421_ ;
	wire _w4420_ ;
	wire _w4419_ ;
	wire _w4418_ ;
	wire _w4417_ ;
	wire _w4416_ ;
	wire _w4415_ ;
	wire _w4414_ ;
	wire _w4413_ ;
	wire _w4412_ ;
	wire _w4411_ ;
	wire _w4410_ ;
	wire _w4409_ ;
	wire _w4408_ ;
	wire _w4407_ ;
	wire _w4406_ ;
	wire _w4405_ ;
	wire _w4404_ ;
	wire _w4403_ ;
	wire _w4402_ ;
	wire _w4401_ ;
	wire _w4400_ ;
	wire _w4399_ ;
	wire _w4398_ ;
	wire _w4397_ ;
	wire _w4396_ ;
	wire _w4395_ ;
	wire _w4394_ ;
	wire _w4393_ ;
	wire _w4392_ ;
	wire _w4391_ ;
	wire _w4390_ ;
	wire _w4389_ ;
	wire _w4388_ ;
	wire _w4387_ ;
	wire _w4386_ ;
	wire _w4385_ ;
	wire _w4384_ ;
	wire _w4383_ ;
	wire _w4382_ ;
	wire _w4381_ ;
	wire _w4380_ ;
	wire _w4379_ ;
	wire _w4378_ ;
	wire _w4377_ ;
	wire _w4376_ ;
	wire _w4375_ ;
	wire _w4374_ ;
	wire _w4373_ ;
	wire _w4372_ ;
	wire _w4371_ ;
	wire _w4370_ ;
	wire _w4369_ ;
	wire _w4368_ ;
	wire _w4367_ ;
	wire _w4366_ ;
	wire _w4365_ ;
	wire _w4364_ ;
	wire _w4363_ ;
	wire _w4362_ ;
	wire _w4361_ ;
	wire _w4360_ ;
	wire _w4359_ ;
	wire _w4358_ ;
	wire _w4357_ ;
	wire _w4356_ ;
	wire _w4355_ ;
	wire _w4354_ ;
	wire _w4353_ ;
	wire _w4352_ ;
	wire _w4351_ ;
	wire _w4350_ ;
	wire _w4349_ ;
	wire _w4348_ ;
	wire _w4347_ ;
	wire _w4346_ ;
	wire _w4345_ ;
	wire _w4344_ ;
	wire _w4343_ ;
	wire _w4342_ ;
	wire _w4341_ ;
	wire _w4340_ ;
	wire _w4339_ ;
	wire _w4338_ ;
	wire _w4337_ ;
	wire _w4336_ ;
	wire _w4335_ ;
	wire _w4334_ ;
	wire _w4333_ ;
	wire _w4332_ ;
	wire _w4331_ ;
	wire _w4330_ ;
	wire _w4329_ ;
	wire _w4328_ ;
	wire _w4327_ ;
	wire _w4326_ ;
	wire _w4325_ ;
	wire _w4324_ ;
	wire _w4323_ ;
	wire _w4322_ ;
	wire _w4321_ ;
	wire _w4320_ ;
	wire _w4319_ ;
	wire _w4318_ ;
	wire _w4317_ ;
	wire _w4316_ ;
	wire _w4315_ ;
	wire _w4314_ ;
	wire _w4313_ ;
	wire _w4312_ ;
	wire _w4311_ ;
	wire _w4310_ ;
	wire _w4309_ ;
	wire _w4308_ ;
	wire _w4307_ ;
	wire _w4306_ ;
	wire _w4305_ ;
	wire _w4304_ ;
	wire _w4303_ ;
	wire _w4302_ ;
	wire _w4301_ ;
	wire _w4300_ ;
	wire _w4299_ ;
	wire _w4298_ ;
	wire _w4297_ ;
	wire _w4296_ ;
	wire _w4295_ ;
	wire _w4294_ ;
	wire _w4293_ ;
	wire _w4292_ ;
	wire _w4291_ ;
	wire _w4290_ ;
	wire _w4289_ ;
	wire _w4288_ ;
	wire _w4287_ ;
	wire _w4286_ ;
	wire _w4285_ ;
	wire _w4284_ ;
	wire _w4283_ ;
	wire _w4282_ ;
	wire _w4281_ ;
	wire _w4280_ ;
	wire _w4279_ ;
	wire _w4278_ ;
	wire _w4277_ ;
	wire _w4276_ ;
	wire _w4275_ ;
	wire _w4274_ ;
	wire _w4273_ ;
	wire _w4272_ ;
	wire _w4271_ ;
	wire _w4270_ ;
	wire _w4269_ ;
	wire _w4268_ ;
	wire _w4267_ ;
	wire _w4266_ ;
	wire _w4265_ ;
	wire _w4264_ ;
	wire _w4263_ ;
	wire _w4262_ ;
	wire _w4261_ ;
	wire _w4260_ ;
	wire _w4259_ ;
	wire _w4258_ ;
	wire _w4257_ ;
	wire _w4256_ ;
	wire _w4255_ ;
	wire _w4254_ ;
	wire _w4253_ ;
	wire _w4252_ ;
	wire _w4251_ ;
	wire _w4250_ ;
	wire _w4249_ ;
	wire _w4248_ ;
	wire _w4247_ ;
	wire _w4246_ ;
	wire _w4245_ ;
	wire _w4244_ ;
	wire _w4243_ ;
	wire _w4242_ ;
	wire _w4241_ ;
	wire _w4240_ ;
	wire _w4239_ ;
	wire _w4238_ ;
	wire _w4237_ ;
	wire _w4236_ ;
	wire _w4235_ ;
	wire _w4234_ ;
	wire _w4233_ ;
	wire _w4232_ ;
	wire _w4231_ ;
	wire _w4230_ ;
	wire _w4229_ ;
	wire _w4228_ ;
	wire _w4227_ ;
	wire _w4226_ ;
	wire _w4225_ ;
	wire _w4224_ ;
	wire _w4223_ ;
	wire _w4222_ ;
	wire _w4221_ ;
	wire _w4220_ ;
	wire _w4219_ ;
	wire _w4218_ ;
	wire _w4217_ ;
	wire _w4216_ ;
	wire _w4215_ ;
	wire _w4214_ ;
	wire _w4213_ ;
	wire _w4212_ ;
	wire _w4211_ ;
	wire _w4210_ ;
	wire _w4209_ ;
	wire _w4208_ ;
	wire _w4207_ ;
	wire _w4206_ ;
	wire _w4205_ ;
	wire _w4204_ ;
	wire _w4203_ ;
	wire _w4202_ ;
	wire _w4201_ ;
	wire _w4200_ ;
	wire _w4199_ ;
	wire _w4198_ ;
	wire _w4197_ ;
	wire _w4196_ ;
	wire _w4195_ ;
	wire _w4194_ ;
	wire _w4193_ ;
	wire _w4192_ ;
	wire _w4191_ ;
	wire _w4190_ ;
	wire _w4189_ ;
	wire _w4188_ ;
	wire _w4187_ ;
	wire _w4186_ ;
	wire _w4185_ ;
	wire _w4184_ ;
	wire _w4183_ ;
	wire _w4182_ ;
	wire _w4181_ ;
	wire _w4180_ ;
	wire _w4179_ ;
	wire _w4178_ ;
	wire _w4177_ ;
	wire _w4176_ ;
	wire _w4175_ ;
	wire _w4174_ ;
	wire _w4173_ ;
	wire _w4172_ ;
	wire _w4171_ ;
	wire _w4170_ ;
	wire _w4169_ ;
	wire _w4168_ ;
	wire _w4167_ ;
	wire _w4166_ ;
	wire _w4165_ ;
	wire _w4164_ ;
	wire _w4163_ ;
	wire _w4162_ ;
	wire _w4161_ ;
	wire _w4160_ ;
	wire _w4159_ ;
	wire _w4158_ ;
	wire _w4157_ ;
	wire _w4156_ ;
	wire _w4155_ ;
	wire _w4154_ ;
	wire _w4153_ ;
	wire _w4152_ ;
	wire _w4151_ ;
	wire _w4150_ ;
	wire _w4149_ ;
	wire _w4148_ ;
	wire _w4147_ ;
	wire _w4146_ ;
	wire _w4145_ ;
	wire _w4144_ ;
	wire _w4143_ ;
	wire _w4142_ ;
	wire _w4141_ ;
	wire _w4140_ ;
	wire _w4139_ ;
	wire _w4138_ ;
	wire _w4137_ ;
	wire _w4136_ ;
	wire _w4135_ ;
	wire _w4134_ ;
	wire _w4133_ ;
	wire _w4132_ ;
	wire _w4131_ ;
	wire _w4130_ ;
	wire _w4129_ ;
	wire _w4128_ ;
	wire _w4127_ ;
	wire _w4126_ ;
	wire _w4125_ ;
	wire _w4124_ ;
	wire _w4123_ ;
	wire _w4122_ ;
	wire _w4121_ ;
	wire _w4120_ ;
	wire _w4119_ ;
	wire _w4118_ ;
	wire _w4117_ ;
	wire _w4116_ ;
	wire _w4115_ ;
	wire _w4114_ ;
	wire _w4113_ ;
	wire _w4112_ ;
	wire _w4111_ ;
	wire _w4110_ ;
	wire _w4109_ ;
	wire _w4108_ ;
	wire _w4107_ ;
	wire _w4106_ ;
	wire _w4105_ ;
	wire _w4104_ ;
	wire _w4103_ ;
	wire _w4102_ ;
	wire _w4101_ ;
	wire _w4100_ ;
	wire _w4099_ ;
	wire _w4098_ ;
	wire _w4097_ ;
	wire _w4096_ ;
	wire _w4095_ ;
	wire _w4094_ ;
	wire _w4093_ ;
	wire _w4092_ ;
	wire _w4091_ ;
	wire _w4090_ ;
	wire _w4089_ ;
	wire _w4088_ ;
	wire _w4087_ ;
	wire _w4086_ ;
	wire _w4085_ ;
	wire _w4084_ ;
	wire _w4083_ ;
	wire _w4082_ ;
	wire _w4081_ ;
	wire _w4080_ ;
	wire _w4079_ ;
	wire _w4078_ ;
	wire _w4077_ ;
	wire _w4076_ ;
	wire _w4075_ ;
	wire _w4074_ ;
	wire _w4073_ ;
	wire _w4072_ ;
	wire _w4071_ ;
	wire _w4070_ ;
	wire _w4069_ ;
	wire _w4068_ ;
	wire _w4067_ ;
	wire _w4066_ ;
	wire _w4065_ ;
	wire _w4064_ ;
	wire _w4063_ ;
	wire _w4062_ ;
	wire _w4061_ ;
	wire _w4060_ ;
	wire _w4059_ ;
	wire _w4058_ ;
	wire _w4057_ ;
	wire _w4056_ ;
	wire _w4055_ ;
	wire _w4054_ ;
	wire _w4053_ ;
	wire _w4052_ ;
	wire _w4051_ ;
	wire _w4050_ ;
	wire _w4049_ ;
	wire _w4048_ ;
	wire _w4047_ ;
	wire _w4046_ ;
	wire _w4045_ ;
	wire _w4044_ ;
	wire _w4043_ ;
	wire _w4042_ ;
	wire _w4041_ ;
	wire _w4040_ ;
	wire _w4039_ ;
	wire _w4038_ ;
	wire _w4037_ ;
	wire _w4036_ ;
	wire _w4035_ ;
	wire _w4034_ ;
	wire _w4033_ ;
	wire _w4032_ ;
	wire _w4031_ ;
	wire _w4030_ ;
	wire _w4029_ ;
	wire _w4028_ ;
	wire _w4027_ ;
	wire _w4026_ ;
	wire _w4025_ ;
	wire _w4024_ ;
	wire _w4023_ ;
	wire _w4022_ ;
	wire _w4021_ ;
	wire _w4020_ ;
	wire _w4019_ ;
	wire _w4018_ ;
	wire _w4017_ ;
	wire _w4016_ ;
	wire _w4015_ ;
	wire _w4014_ ;
	wire _w4013_ ;
	wire _w4012_ ;
	wire _w4011_ ;
	wire _w4010_ ;
	wire _w4009_ ;
	wire _w4008_ ;
	wire _w4007_ ;
	wire _w4006_ ;
	wire _w4005_ ;
	wire _w4004_ ;
	wire _w4003_ ;
	wire _w4002_ ;
	wire _w4001_ ;
	wire _w4000_ ;
	wire _w3999_ ;
	wire _w3998_ ;
	wire _w3997_ ;
	wire _w3996_ ;
	wire _w3995_ ;
	wire _w3994_ ;
	wire _w3993_ ;
	wire _w3992_ ;
	wire _w3991_ ;
	wire _w3990_ ;
	wire _w3989_ ;
	wire _w3988_ ;
	wire _w3987_ ;
	wire _w3986_ ;
	wire _w3985_ ;
	wire _w3984_ ;
	wire _w3983_ ;
	wire _w3982_ ;
	wire _w3981_ ;
	wire _w3980_ ;
	wire _w3979_ ;
	wire _w3978_ ;
	wire _w3977_ ;
	wire _w3976_ ;
	wire _w3975_ ;
	wire _w3974_ ;
	wire _w3973_ ;
	wire _w3972_ ;
	wire _w3971_ ;
	wire _w3970_ ;
	wire _w3969_ ;
	wire _w3968_ ;
	wire _w3967_ ;
	wire _w3966_ ;
	wire _w3965_ ;
	wire _w3964_ ;
	wire _w3963_ ;
	wire _w3962_ ;
	wire _w3961_ ;
	wire _w3960_ ;
	wire _w3959_ ;
	wire _w3958_ ;
	wire _w3957_ ;
	wire _w3956_ ;
	wire _w3955_ ;
	wire _w3954_ ;
	wire _w3953_ ;
	wire _w3952_ ;
	wire _w3951_ ;
	wire _w3950_ ;
	wire _w3949_ ;
	wire _w3948_ ;
	wire _w3947_ ;
	wire _w3946_ ;
	wire _w3945_ ;
	wire _w3944_ ;
	wire _w3943_ ;
	wire _w3942_ ;
	wire _w3941_ ;
	wire _w3940_ ;
	wire _w3939_ ;
	wire _w3938_ ;
	wire _w3937_ ;
	wire _w3936_ ;
	wire _w3935_ ;
	wire _w3934_ ;
	wire _w3933_ ;
	wire _w3932_ ;
	wire _w3931_ ;
	wire _w3930_ ;
	wire _w3929_ ;
	wire _w3928_ ;
	wire _w3927_ ;
	wire _w3926_ ;
	wire _w3925_ ;
	wire _w3924_ ;
	wire _w3923_ ;
	wire _w3922_ ;
	wire _w3921_ ;
	wire _w3920_ ;
	wire _w3919_ ;
	wire _w3918_ ;
	wire _w3917_ ;
	wire _w3916_ ;
	wire _w3915_ ;
	wire _w3914_ ;
	wire _w3913_ ;
	wire _w3912_ ;
	wire _w3911_ ;
	wire _w3910_ ;
	wire _w3909_ ;
	wire _w3908_ ;
	wire _w3907_ ;
	wire _w3906_ ;
	wire _w3905_ ;
	wire _w3904_ ;
	wire _w3903_ ;
	wire _w3902_ ;
	wire _w3901_ ;
	wire _w3900_ ;
	wire _w3899_ ;
	wire _w3898_ ;
	wire _w3897_ ;
	wire _w3896_ ;
	wire _w3895_ ;
	wire _w3894_ ;
	wire _w3893_ ;
	wire _w3892_ ;
	wire _w3891_ ;
	wire _w3890_ ;
	wire _w3889_ ;
	wire _w3888_ ;
	wire _w3887_ ;
	wire _w3886_ ;
	wire _w3885_ ;
	wire _w3884_ ;
	wire _w3883_ ;
	wire _w3882_ ;
	wire _w3881_ ;
	wire _w3880_ ;
	wire _w3879_ ;
	wire _w3878_ ;
	wire _w3877_ ;
	wire _w3876_ ;
	wire _w3875_ ;
	wire _w3874_ ;
	wire _w3873_ ;
	wire _w3872_ ;
	wire _w3871_ ;
	wire _w3870_ ;
	wire _w3869_ ;
	wire _w3868_ ;
	wire _w3867_ ;
	wire _w3866_ ;
	wire _w3865_ ;
	wire _w3864_ ;
	wire _w3863_ ;
	wire _w3862_ ;
	wire _w3861_ ;
	wire _w3860_ ;
	wire _w3859_ ;
	wire _w3858_ ;
	wire _w3857_ ;
	wire _w3856_ ;
	wire _w3855_ ;
	wire _w3854_ ;
	wire _w3853_ ;
	wire _w3852_ ;
	wire _w3851_ ;
	wire _w3850_ ;
	wire _w3849_ ;
	wire _w3848_ ;
	wire _w3847_ ;
	wire _w3846_ ;
	wire _w3845_ ;
	wire _w3844_ ;
	wire _w3843_ ;
	wire _w3842_ ;
	wire _w3841_ ;
	wire _w3840_ ;
	wire _w3839_ ;
	wire _w3838_ ;
	wire _w3837_ ;
	wire _w3836_ ;
	wire _w3835_ ;
	wire _w3834_ ;
	wire _w3833_ ;
	wire _w3832_ ;
	wire _w3831_ ;
	wire _w3830_ ;
	wire _w3829_ ;
	wire _w3828_ ;
	wire _w3827_ ;
	wire _w3826_ ;
	wire _w3825_ ;
	wire _w3824_ ;
	wire _w3823_ ;
	wire _w3822_ ;
	wire _w3821_ ;
	wire _w3820_ ;
	wire _w3819_ ;
	wire _w3818_ ;
	wire _w3817_ ;
	wire _w3816_ ;
	wire _w3815_ ;
	wire _w3814_ ;
	wire _w3813_ ;
	wire _w3812_ ;
	wire _w3811_ ;
	wire _w3810_ ;
	wire _w3809_ ;
	wire _w3808_ ;
	wire _w3807_ ;
	wire _w3806_ ;
	wire _w3805_ ;
	wire _w3804_ ;
	wire _w3803_ ;
	wire _w3802_ ;
	wire _w3801_ ;
	wire _w3800_ ;
	wire _w3799_ ;
	wire _w3798_ ;
	wire _w3797_ ;
	wire _w3796_ ;
	wire _w3795_ ;
	wire _w3794_ ;
	wire _w3793_ ;
	wire _w3792_ ;
	wire _w3791_ ;
	wire _w3790_ ;
	wire _w3789_ ;
	wire _w3788_ ;
	wire _w3787_ ;
	wire _w3786_ ;
	wire _w3785_ ;
	wire _w3784_ ;
	wire _w3783_ ;
	wire _w3782_ ;
	wire _w3781_ ;
	wire _w3780_ ;
	wire _w3779_ ;
	wire _w3778_ ;
	wire _w3777_ ;
	wire _w3776_ ;
	wire _w3775_ ;
	wire _w3774_ ;
	wire _w3773_ ;
	wire _w3772_ ;
	wire _w3771_ ;
	wire _w3770_ ;
	wire _w3769_ ;
	wire _w3768_ ;
	wire _w3767_ ;
	wire _w3766_ ;
	wire _w3765_ ;
	wire _w3764_ ;
	wire _w3763_ ;
	wire _w3762_ ;
	wire _w3761_ ;
	wire _w3760_ ;
	wire _w3759_ ;
	wire _w3758_ ;
	wire _w3757_ ;
	wire _w3756_ ;
	wire _w3755_ ;
	wire _w3754_ ;
	wire _w3753_ ;
	wire _w3752_ ;
	wire _w3751_ ;
	wire _w3750_ ;
	wire _w3749_ ;
	wire _w3748_ ;
	wire _w3747_ ;
	wire _w3746_ ;
	wire _w3745_ ;
	wire _w3744_ ;
	wire _w3743_ ;
	wire _w3742_ ;
	wire _w3741_ ;
	wire _w3740_ ;
	wire _w3739_ ;
	wire _w3738_ ;
	wire _w3737_ ;
	wire _w3736_ ;
	wire _w3735_ ;
	wire _w3734_ ;
	wire _w3733_ ;
	wire _w3732_ ;
	wire _w3731_ ;
	wire _w3730_ ;
	wire _w3729_ ;
	wire _w3728_ ;
	wire _w3727_ ;
	wire _w3726_ ;
	wire _w3725_ ;
	wire _w3724_ ;
	wire _w3723_ ;
	wire _w3722_ ;
	wire _w3721_ ;
	wire _w3720_ ;
	wire _w3719_ ;
	wire _w3718_ ;
	wire _w3717_ ;
	wire _w3716_ ;
	wire _w3715_ ;
	wire _w3714_ ;
	wire _w3713_ ;
	wire _w3712_ ;
	wire _w3711_ ;
	wire _w3710_ ;
	wire _w3709_ ;
	wire _w3708_ ;
	wire _w3707_ ;
	wire _w3706_ ;
	wire _w3705_ ;
	wire _w3704_ ;
	wire _w3703_ ;
	wire _w3702_ ;
	wire _w3701_ ;
	wire _w3700_ ;
	wire _w3699_ ;
	wire _w3698_ ;
	wire _w3697_ ;
	wire _w3696_ ;
	wire _w3695_ ;
	wire _w3694_ ;
	wire _w3693_ ;
	wire _w3692_ ;
	wire _w3691_ ;
	wire _w3690_ ;
	wire _w3689_ ;
	wire _w3688_ ;
	wire _w3687_ ;
	wire _w3686_ ;
	wire _w3685_ ;
	wire _w3684_ ;
	wire _w3683_ ;
	wire _w3682_ ;
	wire _w3681_ ;
	wire _w3680_ ;
	wire _w3679_ ;
	wire _w3678_ ;
	wire _w3677_ ;
	wire _w3676_ ;
	wire _w3675_ ;
	wire _w3674_ ;
	wire _w3673_ ;
	wire _w3672_ ;
	wire _w3671_ ;
	wire _w3670_ ;
	wire _w3669_ ;
	wire _w3668_ ;
	wire _w3667_ ;
	wire _w3666_ ;
	wire _w3665_ ;
	wire _w3664_ ;
	wire _w3663_ ;
	wire _w3662_ ;
	wire _w3661_ ;
	wire _w3660_ ;
	wire _w3659_ ;
	wire _w3658_ ;
	wire _w3657_ ;
	wire _w3656_ ;
	wire _w3655_ ;
	wire _w3654_ ;
	wire _w3653_ ;
	wire _w3652_ ;
	wire _w3651_ ;
	wire _w3650_ ;
	wire _w3649_ ;
	wire _w3648_ ;
	wire _w3647_ ;
	wire _w3646_ ;
	wire _w3645_ ;
	wire _w3644_ ;
	wire _w3643_ ;
	wire _w3642_ ;
	wire _w3641_ ;
	wire _w3640_ ;
	wire _w3639_ ;
	wire _w3638_ ;
	wire _w3637_ ;
	wire _w3636_ ;
	wire _w3635_ ;
	wire _w3634_ ;
	wire _w3633_ ;
	wire _w3632_ ;
	wire _w3631_ ;
	wire _w3630_ ;
	wire _w3629_ ;
	wire _w3628_ ;
	wire _w3627_ ;
	wire _w3626_ ;
	wire _w3625_ ;
	wire _w3624_ ;
	wire _w3623_ ;
	wire _w3622_ ;
	wire _w3621_ ;
	wire _w3620_ ;
	wire _w3619_ ;
	wire _w3618_ ;
	wire _w3617_ ;
	wire _w3616_ ;
	wire _w3615_ ;
	wire _w3614_ ;
	wire _w3613_ ;
	wire _w3612_ ;
	wire _w3611_ ;
	wire _w3610_ ;
	wire _w3609_ ;
	wire _w3608_ ;
	wire _w3607_ ;
	wire _w3606_ ;
	wire _w3605_ ;
	wire _w3604_ ;
	wire _w3603_ ;
	wire _w3602_ ;
	wire _w3601_ ;
	wire _w3600_ ;
	wire _w3599_ ;
	wire _w3598_ ;
	wire _w3597_ ;
	wire _w3596_ ;
	wire _w3595_ ;
	wire _w3594_ ;
	wire _w3593_ ;
	wire _w3592_ ;
	wire _w3591_ ;
	wire _w3590_ ;
	wire _w3589_ ;
	wire _w3588_ ;
	wire _w3587_ ;
	wire _w3586_ ;
	wire _w3585_ ;
	wire _w3584_ ;
	wire _w3583_ ;
	wire _w3582_ ;
	wire _w3581_ ;
	wire _w3580_ ;
	wire _w3579_ ;
	wire _w3578_ ;
	wire _w3577_ ;
	wire _w3576_ ;
	wire _w3575_ ;
	wire _w3574_ ;
	wire _w3573_ ;
	wire _w3572_ ;
	wire _w3571_ ;
	wire _w3570_ ;
	wire _w3569_ ;
	wire _w3568_ ;
	wire _w3567_ ;
	wire _w3566_ ;
	wire _w3565_ ;
	wire _w3564_ ;
	wire _w3563_ ;
	wire _w3562_ ;
	wire _w3561_ ;
	wire _w3560_ ;
	wire _w3559_ ;
	wire _w3558_ ;
	wire _w3557_ ;
	wire _w3556_ ;
	wire _w3555_ ;
	wire _w3554_ ;
	wire _w3553_ ;
	wire _w3552_ ;
	wire _w3551_ ;
	wire _w3550_ ;
	wire _w3549_ ;
	wire _w3548_ ;
	wire _w3547_ ;
	wire _w3546_ ;
	wire _w3545_ ;
	wire _w3544_ ;
	wire _w3543_ ;
	wire _w3542_ ;
	wire _w3541_ ;
	wire _w3540_ ;
	wire _w3539_ ;
	wire _w3538_ ;
	wire _w3537_ ;
	wire _w3536_ ;
	wire _w3535_ ;
	wire _w3534_ ;
	wire _w3533_ ;
	wire _w3532_ ;
	wire _w3531_ ;
	wire _w3530_ ;
	wire _w3529_ ;
	wire _w3528_ ;
	wire _w3527_ ;
	wire _w3526_ ;
	wire _w3525_ ;
	wire _w3524_ ;
	wire _w3523_ ;
	wire _w3522_ ;
	wire _w3521_ ;
	wire _w3520_ ;
	wire _w3519_ ;
	wire _w3518_ ;
	wire _w3517_ ;
	wire _w3516_ ;
	wire _w3515_ ;
	wire _w3514_ ;
	wire _w3513_ ;
	wire _w3512_ ;
	wire _w3511_ ;
	wire _w3510_ ;
	wire _w3509_ ;
	wire _w3508_ ;
	wire _w3507_ ;
	wire _w3506_ ;
	wire _w3505_ ;
	wire _w3504_ ;
	wire _w3503_ ;
	wire _w3502_ ;
	wire _w3501_ ;
	wire _w3500_ ;
	wire _w3499_ ;
	wire _w3498_ ;
	wire _w3497_ ;
	wire _w3496_ ;
	wire _w3495_ ;
	wire _w3494_ ;
	wire _w3493_ ;
	wire _w3492_ ;
	wire _w3491_ ;
	wire _w3490_ ;
	wire _w3489_ ;
	wire _w3488_ ;
	wire _w3487_ ;
	wire _w3486_ ;
	wire _w3485_ ;
	wire _w3484_ ;
	wire _w3483_ ;
	wire _w3482_ ;
	wire _w3481_ ;
	wire _w3480_ ;
	wire _w3479_ ;
	wire _w3478_ ;
	wire _w3477_ ;
	wire _w3476_ ;
	wire _w3475_ ;
	wire _w3474_ ;
	wire _w3473_ ;
	wire _w3472_ ;
	wire _w3471_ ;
	wire _w3470_ ;
	wire _w3469_ ;
	wire _w3468_ ;
	wire _w3467_ ;
	wire _w3466_ ;
	wire _w3465_ ;
	wire _w3464_ ;
	wire _w3463_ ;
	wire _w3462_ ;
	wire _w3461_ ;
	wire _w3460_ ;
	wire _w3459_ ;
	wire _w3458_ ;
	wire _w3457_ ;
	wire _w3456_ ;
	wire _w3455_ ;
	wire _w3454_ ;
	wire _w3453_ ;
	wire _w3452_ ;
	wire _w3451_ ;
	wire _w3450_ ;
	wire _w3449_ ;
	wire _w3448_ ;
	wire _w3447_ ;
	wire _w3446_ ;
	wire _w3445_ ;
	wire _w3444_ ;
	wire _w3443_ ;
	wire _w3442_ ;
	wire _w3441_ ;
	wire _w3440_ ;
	wire _w3439_ ;
	wire _w3438_ ;
	wire _w3437_ ;
	wire _w3436_ ;
	wire _w3435_ ;
	wire _w3434_ ;
	wire _w3433_ ;
	wire _w3432_ ;
	wire _w3431_ ;
	wire _w3430_ ;
	wire _w3429_ ;
	wire _w3428_ ;
	wire _w3427_ ;
	wire _w3426_ ;
	wire _w3425_ ;
	wire _w3424_ ;
	wire _w3423_ ;
	wire _w3422_ ;
	wire _w3421_ ;
	wire _w3420_ ;
	wire _w3419_ ;
	wire _w3418_ ;
	wire _w3417_ ;
	wire _w3416_ ;
	wire _w3415_ ;
	wire _w3414_ ;
	wire _w3413_ ;
	wire _w3412_ ;
	wire _w3411_ ;
	wire _w3410_ ;
	wire _w3409_ ;
	wire _w3408_ ;
	wire _w3407_ ;
	wire _w3406_ ;
	wire _w3405_ ;
	wire _w3404_ ;
	wire _w3403_ ;
	wire _w3402_ ;
	wire _w3401_ ;
	wire _w3400_ ;
	wire _w3399_ ;
	wire _w3398_ ;
	wire _w3397_ ;
	wire _w3396_ ;
	wire _w3395_ ;
	wire _w3394_ ;
	wire _w3393_ ;
	wire _w3392_ ;
	wire _w3391_ ;
	wire _w3390_ ;
	wire _w3389_ ;
	wire _w3388_ ;
	wire _w3387_ ;
	wire _w3386_ ;
	wire _w3385_ ;
	wire _w3384_ ;
	wire _w3383_ ;
	wire _w3382_ ;
	wire _w3381_ ;
	wire _w3380_ ;
	wire _w3379_ ;
	wire _w3378_ ;
	wire _w3377_ ;
	wire _w3376_ ;
	wire _w3375_ ;
	wire _w3374_ ;
	wire _w3373_ ;
	wire _w3372_ ;
	wire _w3371_ ;
	wire _w3370_ ;
	wire _w3369_ ;
	wire _w3368_ ;
	wire _w3367_ ;
	wire _w3366_ ;
	wire _w3365_ ;
	wire _w3364_ ;
	wire _w3363_ ;
	wire _w3362_ ;
	wire _w3361_ ;
	wire _w3360_ ;
	wire _w3359_ ;
	wire _w3358_ ;
	wire _w3357_ ;
	wire _w3356_ ;
	wire _w3355_ ;
	wire _w3354_ ;
	wire _w3353_ ;
	wire _w3352_ ;
	wire _w3351_ ;
	wire _w3350_ ;
	wire _w3349_ ;
	wire _w3348_ ;
	wire _w3347_ ;
	wire _w3346_ ;
	wire _w3345_ ;
	wire _w3344_ ;
	wire _w3343_ ;
	wire _w3342_ ;
	wire _w3341_ ;
	wire _w3340_ ;
	wire _w3339_ ;
	wire _w3338_ ;
	wire _w3337_ ;
	wire _w3336_ ;
	wire _w3335_ ;
	wire _w3334_ ;
	wire _w3333_ ;
	wire _w3332_ ;
	wire _w3331_ ;
	wire _w3330_ ;
	wire _w3329_ ;
	wire _w3328_ ;
	wire _w3327_ ;
	wire _w3326_ ;
	wire _w3325_ ;
	wire _w3324_ ;
	wire _w3323_ ;
	wire _w3322_ ;
	wire _w3321_ ;
	wire _w3320_ ;
	wire _w3319_ ;
	wire _w3318_ ;
	wire _w3317_ ;
	wire _w3316_ ;
	wire _w3315_ ;
	wire _w3314_ ;
	wire _w3313_ ;
	wire _w3312_ ;
	wire _w3311_ ;
	wire _w3310_ ;
	wire _w3309_ ;
	wire _w3308_ ;
	wire _w3307_ ;
	wire _w3306_ ;
	wire _w3305_ ;
	wire _w3304_ ;
	wire _w3303_ ;
	wire _w3302_ ;
	wire _w3301_ ;
	wire _w3300_ ;
	wire _w3299_ ;
	wire _w3298_ ;
	wire _w3297_ ;
	wire _w3296_ ;
	wire _w3295_ ;
	wire _w3294_ ;
	wire _w3293_ ;
	wire _w3292_ ;
	wire _w3291_ ;
	wire _w3290_ ;
	wire _w3289_ ;
	wire _w3288_ ;
	wire _w3287_ ;
	wire _w3286_ ;
	wire _w3285_ ;
	wire _w3284_ ;
	wire _w3283_ ;
	wire _w3282_ ;
	wire _w3281_ ;
	wire _w3280_ ;
	wire _w3279_ ;
	wire _w3278_ ;
	wire _w3277_ ;
	wire _w3276_ ;
	wire _w3275_ ;
	wire _w3274_ ;
	wire _w3273_ ;
	wire _w3272_ ;
	wire _w3271_ ;
	wire _w3270_ ;
	wire _w3269_ ;
	wire _w3268_ ;
	wire _w3267_ ;
	wire _w3266_ ;
	wire _w3265_ ;
	wire _w3264_ ;
	wire _w3263_ ;
	wire _w3262_ ;
	wire _w3261_ ;
	wire _w3260_ ;
	wire _w3259_ ;
	wire _w3258_ ;
	wire _w3257_ ;
	wire _w3256_ ;
	wire _w3255_ ;
	wire _w3254_ ;
	wire _w3253_ ;
	wire _w3252_ ;
	wire _w3251_ ;
	wire _w3250_ ;
	wire _w3249_ ;
	wire _w3248_ ;
	wire _w3247_ ;
	wire _w3246_ ;
	wire _w3245_ ;
	wire _w3244_ ;
	wire _w3243_ ;
	wire _w3242_ ;
	wire _w3241_ ;
	wire _w3240_ ;
	wire _w3239_ ;
	wire _w3238_ ;
	wire _w3237_ ;
	wire _w3236_ ;
	wire _w3235_ ;
	wire _w3234_ ;
	wire _w3233_ ;
	wire _w3232_ ;
	wire _w3231_ ;
	wire _w3230_ ;
	wire _w3229_ ;
	wire _w3228_ ;
	wire _w3227_ ;
	wire _w3226_ ;
	wire _w3225_ ;
	wire _w3224_ ;
	wire _w3223_ ;
	wire _w3222_ ;
	wire _w3221_ ;
	wire _w3220_ ;
	wire _w3219_ ;
	wire _w3218_ ;
	wire _w3217_ ;
	wire _w3216_ ;
	wire _w3215_ ;
	wire _w3214_ ;
	wire _w3213_ ;
	wire _w3212_ ;
	wire _w3211_ ;
	wire _w3210_ ;
	wire _w3209_ ;
	wire _w3208_ ;
	wire _w3207_ ;
	wire _w3206_ ;
	wire _w3205_ ;
	wire _w3204_ ;
	wire _w3203_ ;
	wire _w3202_ ;
	wire _w3201_ ;
	wire _w3200_ ;
	wire _w3199_ ;
	wire _w3198_ ;
	wire _w3197_ ;
	wire _w3196_ ;
	wire _w3195_ ;
	wire _w3194_ ;
	wire _w3193_ ;
	wire _w3192_ ;
	wire _w3191_ ;
	wire _w3190_ ;
	wire _w3189_ ;
	wire _w3188_ ;
	wire _w3187_ ;
	wire _w3186_ ;
	wire _w3185_ ;
	wire _w3184_ ;
	wire _w3183_ ;
	wire _w3182_ ;
	wire _w3181_ ;
	wire _w3180_ ;
	wire _w3179_ ;
	wire _w3178_ ;
	wire _w3177_ ;
	wire _w3176_ ;
	wire _w3175_ ;
	wire _w3174_ ;
	wire _w3173_ ;
	wire _w3172_ ;
	wire _w3171_ ;
	wire _w3170_ ;
	wire _w3169_ ;
	wire _w3168_ ;
	wire _w3167_ ;
	wire _w3166_ ;
	wire _w3165_ ;
	wire _w3164_ ;
	wire _w3163_ ;
	wire _w3162_ ;
	wire _w3161_ ;
	wire _w3160_ ;
	wire _w3159_ ;
	wire _w3158_ ;
	wire _w3157_ ;
	wire _w3156_ ;
	wire _w3155_ ;
	wire _w3154_ ;
	wire _w3153_ ;
	wire _w3152_ ;
	wire _w3151_ ;
	wire _w3150_ ;
	wire _w3149_ ;
	wire _w3148_ ;
	wire _w3147_ ;
	wire _w3146_ ;
	wire _w3145_ ;
	wire _w3144_ ;
	wire _w3143_ ;
	wire _w3142_ ;
	wire _w3141_ ;
	wire _w3140_ ;
	wire _w3139_ ;
	wire _w3138_ ;
	wire _w3137_ ;
	wire _w3136_ ;
	wire _w3135_ ;
	wire _w3134_ ;
	wire _w3133_ ;
	wire _w3132_ ;
	wire _w3131_ ;
	wire _w3130_ ;
	wire _w3129_ ;
	wire _w3128_ ;
	wire _w3127_ ;
	wire _w3126_ ;
	wire _w3125_ ;
	wire _w3124_ ;
	wire _w3123_ ;
	wire _w3122_ ;
	wire _w3121_ ;
	wire _w3120_ ;
	wire _w3119_ ;
	wire _w3118_ ;
	wire _w3117_ ;
	wire _w3116_ ;
	wire _w3115_ ;
	wire _w3114_ ;
	wire _w3113_ ;
	wire _w3112_ ;
	wire _w3111_ ;
	wire _w3110_ ;
	wire _w3109_ ;
	wire _w3108_ ;
	wire _w3107_ ;
	wire _w3106_ ;
	wire _w3105_ ;
	wire _w3104_ ;
	wire _w3103_ ;
	wire _w3102_ ;
	wire _w3101_ ;
	wire _w3100_ ;
	wire _w3099_ ;
	wire _w3098_ ;
	wire _w3097_ ;
	wire _w3096_ ;
	wire _w3095_ ;
	wire _w3094_ ;
	wire _w3093_ ;
	wire _w3092_ ;
	wire _w3091_ ;
	wire _w3090_ ;
	wire _w3089_ ;
	wire _w3088_ ;
	wire _w3087_ ;
	wire _w3086_ ;
	wire _w3085_ ;
	wire _w3084_ ;
	wire _w3083_ ;
	wire _w3082_ ;
	wire _w3081_ ;
	wire _w3080_ ;
	wire _w3079_ ;
	wire _w3078_ ;
	wire _w3077_ ;
	wire _w3076_ ;
	wire _w3075_ ;
	wire _w3074_ ;
	wire _w3073_ ;
	wire _w3072_ ;
	wire _w3071_ ;
	wire _w3070_ ;
	wire _w3069_ ;
	wire _w3068_ ;
	wire _w3067_ ;
	wire _w3066_ ;
	wire _w3065_ ;
	wire _w3064_ ;
	wire _w3063_ ;
	wire _w3062_ ;
	wire _w3061_ ;
	wire _w3060_ ;
	wire _w3059_ ;
	wire _w3058_ ;
	wire _w3057_ ;
	wire _w3056_ ;
	wire _w3055_ ;
	wire _w3054_ ;
	wire _w3053_ ;
	wire _w3052_ ;
	wire _w3051_ ;
	wire _w3050_ ;
	wire _w3049_ ;
	wire _w3048_ ;
	wire _w3047_ ;
	wire _w3046_ ;
	wire _w3045_ ;
	wire _w3044_ ;
	wire _w3043_ ;
	wire _w3042_ ;
	wire _w3041_ ;
	wire _w3040_ ;
	wire _w3039_ ;
	wire _w3038_ ;
	wire _w3037_ ;
	wire _w3036_ ;
	wire _w3035_ ;
	wire _w3034_ ;
	wire _w3033_ ;
	wire _w3032_ ;
	wire _w3031_ ;
	wire _w3030_ ;
	wire _w3029_ ;
	wire _w3028_ ;
	wire _w3027_ ;
	wire _w3026_ ;
	wire _w3025_ ;
	wire _w3024_ ;
	wire _w3023_ ;
	wire _w3022_ ;
	wire _w3021_ ;
	wire _w3020_ ;
	wire _w3019_ ;
	wire _w3018_ ;
	wire _w3017_ ;
	wire _w3016_ ;
	wire _w3015_ ;
	wire _w3014_ ;
	wire _w3013_ ;
	wire _w3012_ ;
	wire _w3011_ ;
	wire _w3010_ ;
	wire _w3009_ ;
	wire _w3008_ ;
	wire _w3007_ ;
	wire _w3006_ ;
	wire _w3005_ ;
	wire _w3004_ ;
	wire _w3003_ ;
	wire _w3002_ ;
	wire _w3001_ ;
	wire _w3000_ ;
	wire _w2999_ ;
	wire _w2998_ ;
	wire _w2997_ ;
	wire _w2996_ ;
	wire _w2995_ ;
	wire _w2994_ ;
	wire _w2993_ ;
	wire _w2992_ ;
	wire _w2991_ ;
	wire _w2990_ ;
	wire _w2989_ ;
	wire _w2988_ ;
	wire _w2987_ ;
	wire _w2986_ ;
	wire _w2985_ ;
	wire _w2984_ ;
	wire _w2983_ ;
	wire _w2982_ ;
	wire _w2981_ ;
	wire _w2980_ ;
	wire _w2979_ ;
	wire _w2978_ ;
	wire _w2977_ ;
	wire _w2976_ ;
	wire _w2975_ ;
	wire _w2974_ ;
	wire _w2973_ ;
	wire _w2972_ ;
	wire _w2971_ ;
	wire _w2970_ ;
	wire _w2969_ ;
	wire _w2968_ ;
	wire _w2967_ ;
	wire _w2966_ ;
	wire _w2965_ ;
	wire _w2964_ ;
	wire _w2963_ ;
	wire _w2962_ ;
	wire _w2961_ ;
	wire _w2960_ ;
	wire _w2959_ ;
	wire _w2958_ ;
	wire _w2957_ ;
	wire _w2956_ ;
	wire _w2955_ ;
	wire _w2954_ ;
	wire _w2953_ ;
	wire _w2952_ ;
	wire _w2951_ ;
	wire _w2950_ ;
	wire _w2949_ ;
	wire _w2948_ ;
	wire _w2947_ ;
	wire _w2946_ ;
	wire _w2945_ ;
	wire _w2944_ ;
	wire _w2943_ ;
	wire _w2942_ ;
	wire _w2941_ ;
	wire _w2940_ ;
	wire _w2939_ ;
	wire _w2938_ ;
	wire _w2937_ ;
	wire _w2936_ ;
	wire _w2935_ ;
	wire _w2934_ ;
	wire _w2933_ ;
	wire _w2932_ ;
	wire _w2931_ ;
	wire _w2930_ ;
	wire _w2929_ ;
	wire _w2928_ ;
	wire _w2927_ ;
	wire _w2926_ ;
	wire _w2925_ ;
	wire _w2924_ ;
	wire _w2923_ ;
	wire _w2922_ ;
	wire _w2921_ ;
	wire _w2920_ ;
	wire _w2919_ ;
	wire _w2918_ ;
	wire _w2917_ ;
	wire _w2916_ ;
	wire _w2915_ ;
	wire _w2914_ ;
	wire _w2913_ ;
	wire _w2912_ ;
	wire _w2911_ ;
	wire _w2910_ ;
	wire _w2909_ ;
	wire _w2908_ ;
	wire _w2907_ ;
	wire _w2906_ ;
	wire _w2905_ ;
	wire _w2904_ ;
	wire _w2903_ ;
	wire _w2902_ ;
	wire _w2901_ ;
	wire _w2900_ ;
	wire _w2899_ ;
	wire _w2898_ ;
	wire _w2897_ ;
	wire _w2896_ ;
	wire _w2895_ ;
	wire _w2894_ ;
	wire _w2893_ ;
	wire _w2892_ ;
	wire _w2891_ ;
	wire _w2890_ ;
	wire _w2889_ ;
	wire _w2888_ ;
	wire _w2887_ ;
	wire _w2886_ ;
	wire _w2885_ ;
	wire _w2884_ ;
	wire _w2883_ ;
	wire _w2882_ ;
	wire _w2881_ ;
	wire _w2880_ ;
	wire _w2879_ ;
	wire _w2878_ ;
	wire _w2877_ ;
	wire _w2876_ ;
	wire _w2875_ ;
	wire _w2874_ ;
	wire _w2873_ ;
	wire _w2872_ ;
	wire _w2871_ ;
	wire _w2870_ ;
	wire _w2869_ ;
	wire _w2868_ ;
	wire _w2867_ ;
	wire _w2866_ ;
	wire _w2865_ ;
	wire _w2864_ ;
	wire _w2863_ ;
	wire _w2862_ ;
	wire _w2861_ ;
	wire _w2860_ ;
	wire _w2859_ ;
	wire _w2858_ ;
	wire _w2857_ ;
	wire _w2856_ ;
	wire _w2855_ ;
	wire _w2854_ ;
	wire _w2853_ ;
	wire _w2852_ ;
	wire _w2851_ ;
	wire _w2850_ ;
	wire _w2849_ ;
	wire _w2848_ ;
	wire _w2847_ ;
	wire _w2846_ ;
	wire _w2845_ ;
	wire _w2844_ ;
	wire _w2843_ ;
	wire _w2842_ ;
	wire _w2841_ ;
	wire _w2840_ ;
	wire _w2839_ ;
	wire _w2838_ ;
	wire _w2837_ ;
	wire _w2836_ ;
	wire _w2835_ ;
	wire _w2834_ ;
	wire _w2833_ ;
	wire _w2832_ ;
	wire _w2831_ ;
	wire _w2830_ ;
	wire _w2829_ ;
	wire _w2828_ ;
	wire _w2827_ ;
	wire _w2826_ ;
	wire _w2825_ ;
	wire _w2824_ ;
	wire _w2823_ ;
	wire _w2822_ ;
	wire _w2821_ ;
	wire _w2820_ ;
	wire _w2819_ ;
	wire _w2818_ ;
	wire _w2817_ ;
	wire _w2816_ ;
	wire _w2815_ ;
	wire _w2814_ ;
	wire _w2813_ ;
	wire _w2812_ ;
	wire _w2811_ ;
	wire _w2810_ ;
	wire _w2809_ ;
	wire _w2808_ ;
	wire _w2807_ ;
	wire _w2806_ ;
	wire _w2805_ ;
	wire _w2804_ ;
	wire _w2803_ ;
	wire _w2802_ ;
	wire _w2801_ ;
	wire _w2800_ ;
	wire _w2799_ ;
	wire _w2798_ ;
	wire _w2797_ ;
	wire _w2796_ ;
	wire _w2795_ ;
	wire _w2794_ ;
	wire _w2793_ ;
	wire _w2792_ ;
	wire _w2791_ ;
	wire _w2790_ ;
	wire _w2789_ ;
	wire _w2788_ ;
	wire _w2787_ ;
	wire _w2786_ ;
	wire _w2785_ ;
	wire _w2784_ ;
	wire _w2783_ ;
	wire _w2782_ ;
	wire _w2781_ ;
	wire _w2780_ ;
	wire _w2779_ ;
	wire _w2778_ ;
	wire _w2777_ ;
	wire _w2776_ ;
	wire _w2775_ ;
	wire _w2774_ ;
	wire _w2773_ ;
	wire _w2772_ ;
	wire _w2771_ ;
	wire _w2770_ ;
	wire _w2769_ ;
	wire _w2768_ ;
	wire _w2767_ ;
	wire _w2766_ ;
	wire _w2765_ ;
	wire _w2764_ ;
	wire _w2763_ ;
	wire _w2762_ ;
	wire _w2761_ ;
	wire _w2760_ ;
	wire _w2759_ ;
	wire _w2758_ ;
	wire _w2757_ ;
	wire _w2756_ ;
	wire _w2755_ ;
	wire _w2754_ ;
	wire _w2753_ ;
	wire _w2752_ ;
	wire _w2751_ ;
	wire _w2750_ ;
	wire _w2749_ ;
	wire _w2748_ ;
	wire _w2747_ ;
	wire _w2746_ ;
	wire _w2745_ ;
	wire _w2744_ ;
	wire _w2743_ ;
	wire _w2742_ ;
	wire _w2741_ ;
	wire _w2740_ ;
	wire _w2739_ ;
	wire _w2738_ ;
	wire _w2737_ ;
	wire _w2736_ ;
	wire _w2735_ ;
	wire _w2734_ ;
	wire _w2733_ ;
	wire _w2732_ ;
	wire _w2731_ ;
	wire _w2730_ ;
	wire _w2729_ ;
	wire _w2728_ ;
	wire _w2727_ ;
	wire _w2726_ ;
	wire _w2725_ ;
	wire _w2724_ ;
	wire _w2723_ ;
	wire _w2722_ ;
	wire _w2721_ ;
	wire _w2720_ ;
	wire _w2719_ ;
	wire _w2718_ ;
	wire _w2717_ ;
	wire _w2716_ ;
	wire _w2715_ ;
	wire _w2714_ ;
	wire _w2713_ ;
	wire _w2712_ ;
	wire _w2711_ ;
	wire _w2710_ ;
	wire _w2709_ ;
	wire _w2708_ ;
	wire _w2707_ ;
	wire _w2706_ ;
	wire _w2705_ ;
	wire _w2704_ ;
	wire _w2703_ ;
	wire _w2702_ ;
	wire _w2701_ ;
	wire _w2700_ ;
	wire _w2699_ ;
	wire _w2698_ ;
	wire _w2697_ ;
	wire _w2696_ ;
	wire _w2695_ ;
	wire _w2694_ ;
	wire _w2693_ ;
	wire _w2692_ ;
	wire _w2691_ ;
	wire _w2690_ ;
	wire _w2689_ ;
	wire _w2688_ ;
	wire _w2687_ ;
	wire _w2686_ ;
	wire _w2685_ ;
	wire _w2684_ ;
	wire _w2683_ ;
	wire _w2682_ ;
	wire _w2681_ ;
	wire _w2680_ ;
	wire _w2679_ ;
	wire _w2678_ ;
	wire _w2677_ ;
	wire _w2676_ ;
	wire _w2675_ ;
	wire _w2674_ ;
	wire _w2673_ ;
	wire _w2672_ ;
	wire _w2671_ ;
	wire _w2670_ ;
	wire _w2669_ ;
	wire _w2668_ ;
	wire _w2667_ ;
	wire _w2666_ ;
	wire _w2665_ ;
	wire _w2664_ ;
	wire _w2663_ ;
	wire _w2662_ ;
	wire _w2661_ ;
	wire _w2660_ ;
	wire _w2659_ ;
	wire _w2658_ ;
	wire _w2657_ ;
	wire _w2656_ ;
	wire _w2655_ ;
	wire _w2654_ ;
	wire _w2653_ ;
	wire _w2652_ ;
	wire _w2651_ ;
	wire _w2650_ ;
	wire _w2649_ ;
	wire _w2648_ ;
	wire _w2647_ ;
	wire _w2646_ ;
	wire _w2645_ ;
	wire _w2644_ ;
	wire _w2643_ ;
	wire _w2642_ ;
	wire _w2641_ ;
	wire _w2640_ ;
	wire _w2639_ ;
	wire _w2638_ ;
	wire _w2637_ ;
	wire _w2636_ ;
	wire _w2635_ ;
	wire _w2634_ ;
	wire _w2633_ ;
	wire _w2632_ ;
	wire _w2631_ ;
	wire _w2630_ ;
	wire _w2629_ ;
	wire _w2628_ ;
	wire _w2627_ ;
	wire _w2626_ ;
	wire _w2625_ ;
	wire _w2624_ ;
	wire _w2623_ ;
	wire _w2622_ ;
	wire _w2621_ ;
	wire _w2620_ ;
	wire _w2619_ ;
	wire _w2618_ ;
	wire _w2617_ ;
	wire _w2616_ ;
	wire _w2615_ ;
	wire _w2614_ ;
	wire _w2613_ ;
	wire _w2612_ ;
	wire _w2611_ ;
	wire _w2610_ ;
	wire _w2609_ ;
	wire _w2608_ ;
	wire _w2607_ ;
	wire _w2606_ ;
	wire _w2605_ ;
	wire _w2604_ ;
	wire _w2603_ ;
	wire _w2602_ ;
	wire _w2601_ ;
	wire _w2600_ ;
	wire _w2599_ ;
	wire _w2598_ ;
	wire _w2597_ ;
	wire _w2596_ ;
	wire _w2595_ ;
	wire _w2594_ ;
	wire _w2593_ ;
	wire _w2592_ ;
	wire _w2591_ ;
	wire _w2590_ ;
	wire _w2589_ ;
	wire _w2588_ ;
	wire _w2587_ ;
	wire _w2586_ ;
	wire _w2585_ ;
	wire _w2584_ ;
	wire _w2583_ ;
	wire _w2582_ ;
	wire _w2581_ ;
	wire _w2580_ ;
	wire _w2579_ ;
	wire _w2578_ ;
	wire _w2577_ ;
	wire _w2576_ ;
	wire _w2575_ ;
	wire _w2574_ ;
	wire _w2573_ ;
	wire _w2572_ ;
	wire _w2571_ ;
	wire _w2570_ ;
	wire _w2569_ ;
	wire _w2568_ ;
	wire _w2567_ ;
	wire _w2566_ ;
	wire _w2565_ ;
	wire _w2564_ ;
	wire _w2563_ ;
	wire _w2562_ ;
	wire _w2561_ ;
	wire _w2560_ ;
	wire _w2559_ ;
	wire _w2558_ ;
	wire _w2557_ ;
	wire _w2556_ ;
	wire _w2555_ ;
	wire _w2554_ ;
	wire _w2553_ ;
	wire _w2552_ ;
	wire _w2551_ ;
	wire _w2550_ ;
	wire _w2549_ ;
	wire _w2548_ ;
	wire _w2547_ ;
	wire _w2546_ ;
	wire _w2545_ ;
	wire _w2544_ ;
	wire _w2543_ ;
	wire _w2542_ ;
	wire _w2541_ ;
	wire _w2540_ ;
	wire _w2539_ ;
	wire _w2538_ ;
	wire _w2537_ ;
	wire _w2536_ ;
	wire _w2535_ ;
	wire _w2534_ ;
	wire _w2533_ ;
	wire _w2532_ ;
	wire _w2531_ ;
	wire _w2530_ ;
	wire _w2529_ ;
	wire _w2528_ ;
	wire _w2527_ ;
	wire _w2526_ ;
	wire _w2525_ ;
	wire _w2524_ ;
	wire _w2523_ ;
	wire _w2522_ ;
	wire _w2521_ ;
	wire _w2520_ ;
	wire _w2519_ ;
	wire _w2518_ ;
	wire _w2517_ ;
	wire _w2516_ ;
	wire _w2515_ ;
	wire _w2514_ ;
	wire _w2513_ ;
	wire _w2512_ ;
	wire _w2511_ ;
	wire _w2510_ ;
	wire _w2509_ ;
	wire _w2508_ ;
	wire _w2507_ ;
	wire _w2506_ ;
	wire _w2505_ ;
	wire _w2504_ ;
	wire _w2503_ ;
	wire _w2502_ ;
	wire _w2501_ ;
	wire _w2500_ ;
	wire _w2499_ ;
	wire _w2498_ ;
	wire _w2497_ ;
	wire _w2496_ ;
	wire _w2495_ ;
	wire _w2494_ ;
	wire _w2493_ ;
	wire _w2492_ ;
	wire _w2491_ ;
	wire _w2490_ ;
	wire _w2489_ ;
	wire _w2488_ ;
	wire _w2487_ ;
	wire _w2486_ ;
	wire _w2485_ ;
	wire _w2484_ ;
	wire _w2483_ ;
	wire _w2482_ ;
	wire _w2481_ ;
	wire _w2480_ ;
	wire _w2479_ ;
	wire _w2478_ ;
	wire _w2477_ ;
	wire _w2476_ ;
	wire _w2475_ ;
	wire _w2474_ ;
	wire _w2473_ ;
	wire _w2472_ ;
	wire _w2471_ ;
	wire _w2470_ ;
	wire _w2469_ ;
	wire _w2468_ ;
	wire _w2467_ ;
	wire _w2466_ ;
	wire _w2465_ ;
	wire _w2464_ ;
	wire _w2463_ ;
	wire _w2462_ ;
	wire _w2461_ ;
	wire _w2460_ ;
	wire _w2459_ ;
	wire _w2458_ ;
	wire _w2457_ ;
	wire _w2456_ ;
	wire _w2455_ ;
	wire _w2454_ ;
	wire _w2453_ ;
	wire _w2452_ ;
	wire _w2451_ ;
	wire _w2450_ ;
	wire _w2449_ ;
	wire _w2448_ ;
	wire _w2447_ ;
	wire _w2446_ ;
	wire _w2445_ ;
	wire _w2444_ ;
	wire _w2443_ ;
	wire _w2442_ ;
	wire _w2441_ ;
	wire _w2440_ ;
	wire _w2439_ ;
	wire _w2438_ ;
	wire _w2437_ ;
	wire _w2436_ ;
	wire _w2435_ ;
	wire _w2434_ ;
	wire _w2433_ ;
	wire _w2432_ ;
	wire _w2431_ ;
	wire _w2430_ ;
	wire _w2429_ ;
	wire _w2428_ ;
	wire _w2427_ ;
	wire _w2426_ ;
	wire _w2425_ ;
	wire _w2424_ ;
	wire _w2423_ ;
	wire _w2422_ ;
	wire _w2421_ ;
	wire _w2420_ ;
	wire _w2419_ ;
	wire _w2418_ ;
	wire _w2417_ ;
	wire _w2416_ ;
	wire _w2415_ ;
	wire _w2414_ ;
	wire _w2413_ ;
	wire _w2412_ ;
	wire _w2411_ ;
	wire _w2410_ ;
	wire _w2409_ ;
	wire _w2408_ ;
	wire _w2407_ ;
	wire _w2406_ ;
	wire _w2405_ ;
	wire _w2404_ ;
	wire _w2403_ ;
	wire _w2402_ ;
	wire _w2401_ ;
	wire _w2400_ ;
	wire _w2399_ ;
	wire _w2398_ ;
	wire _w2397_ ;
	wire _w2396_ ;
	wire _w2395_ ;
	wire _w2394_ ;
	wire _w2393_ ;
	wire _w2392_ ;
	wire _w2391_ ;
	wire _w1142_ ;
	wire _w1141_ ;
	wire _w1140_ ;
	wire _w1139_ ;
	wire _w1138_ ;
	wire _w1137_ ;
	wire _w1136_ ;
	wire _w1135_ ;
	wire _w1134_ ;
	wire _w1133_ ;
	wire _w1132_ ;
	wire _w1131_ ;
	wire _w1130_ ;
	wire _w1129_ ;
	wire _w1128_ ;
	wire _w1127_ ;
	wire _w1126_ ;
	wire _w1125_ ;
	wire _w1124_ ;
	wire _w1123_ ;
	wire _w1122_ ;
	wire _w1121_ ;
	wire _w1120_ ;
	wire _w1119_ ;
	wire _w1118_ ;
	wire _w1117_ ;
	wire _w1116_ ;
	wire _w1115_ ;
	wire _w1114_ ;
	wire _w1113_ ;
	wire _w1112_ ;
	wire _w1111_ ;
	wire _w1110_ ;
	wire _w1109_ ;
	wire _w1108_ ;
	wire _w1107_ ;
	wire _w1106_ ;
	wire _w1105_ ;
	wire _w1104_ ;
	wire _w1103_ ;
	wire _w1102_ ;
	wire _w1101_ ;
	wire _w1100_ ;
	wire _w1099_ ;
	wire _w1098_ ;
	wire _w1097_ ;
	wire _w1096_ ;
	wire _w1095_ ;
	wire _w1094_ ;
	wire _w1093_ ;
	wire _w1092_ ;
	wire _w1091_ ;
	wire _w1090_ ;
	wire _w1089_ ;
	wire _w1088_ ;
	wire _w1087_ ;
	wire _w1086_ ;
	wire _w1085_ ;
	wire _w1084_ ;
	wire _w1083_ ;
	wire _w1082_ ;
	wire _w1081_ ;
	wire _w1080_ ;
	wire _w1079_ ;
	wire _w1078_ ;
	wire _w1077_ ;
	wire _w1076_ ;
	wire _w1075_ ;
	wire _w1074_ ;
	wire _w1073_ ;
	wire _w1072_ ;
	wire _w1071_ ;
	wire _w1070_ ;
	wire _w1069_ ;
	wire _w1068_ ;
	wire _w1067_ ;
	wire _w1066_ ;
	wire _w1065_ ;
	wire _w1064_ ;
	wire _w1063_ ;
	wire _w1062_ ;
	wire _w1061_ ;
	wire _w1060_ ;
	wire _w1059_ ;
	wire _w1058_ ;
	wire _w1057_ ;
	wire _w1056_ ;
	wire _w1055_ ;
	wire _w1054_ ;
	wire _w1053_ ;
	wire _w1052_ ;
	wire _w1051_ ;
	wire _w1050_ ;
	wire _w1049_ ;
	wire _w1048_ ;
	wire _w1047_ ;
	wire _w1046_ ;
	wire _w1045_ ;
	wire _w1044_ ;
	wire _w1043_ ;
	wire _w1042_ ;
	wire _w1041_ ;
	wire _w1040_ ;
	wire _w1039_ ;
	wire _w1038_ ;
	wire _w1037_ ;
	wire _w1036_ ;
	wire _w1035_ ;
	wire _w1034_ ;
	wire _w1033_ ;
	wire _w1032_ ;
	wire _w1031_ ;
	wire _w1030_ ;
	wire _w1029_ ;
	wire _w1028_ ;
	wire _w1027_ ;
	wire _w1026_ ;
	wire _w1025_ ;
	wire _w1024_ ;
	wire _w1023_ ;
	wire _w1022_ ;
	wire _w1021_ ;
	wire _w1020_ ;
	wire _w1019_ ;
	wire _w1018_ ;
	wire _w1017_ ;
	wire _w1016_ ;
	wire _w1015_ ;
	wire _w1014_ ;
	wire _w1013_ ;
	wire _w1012_ ;
	wire _w1011_ ;
	wire _w1010_ ;
	wire _w1009_ ;
	wire _w1008_ ;
	wire _w1007_ ;
	wire _w1006_ ;
	wire _w1005_ ;
	wire _w1004_ ;
	wire _w1003_ ;
	wire _w1002_ ;
	wire _w1001_ ;
	wire _w1000_ ;
	wire _w999_ ;
	wire _w998_ ;
	wire _w997_ ;
	wire _w996_ ;
	wire _w995_ ;
	wire _w994_ ;
	wire _w993_ ;
	wire _w992_ ;
	wire _w991_ ;
	wire _w990_ ;
	wire _w989_ ;
	wire _w988_ ;
	wire _w987_ ;
	wire _w986_ ;
	wire _w985_ ;
	wire _w984_ ;
	wire _w983_ ;
	wire _w982_ ;
	wire _w981_ ;
	wire _w980_ ;
	wire _w979_ ;
	wire _w978_ ;
	wire _w977_ ;
	wire _w976_ ;
	wire _w975_ ;
	wire _w974_ ;
	wire _w973_ ;
	wire _w972_ ;
	wire _w971_ ;
	wire _w970_ ;
	wire _w969_ ;
	wire _w968_ ;
	wire _w967_ ;
	wire _w966_ ;
	wire _w965_ ;
	wire _w964_ ;
	wire _w963_ ;
	wire _w962_ ;
	wire _w961_ ;
	wire _w960_ ;
	wire _w959_ ;
	wire _w958_ ;
	wire _w957_ ;
	wire _w956_ ;
	wire _w955_ ;
	wire _w954_ ;
	wire _w953_ ;
	wire _w952_ ;
	wire _w951_ ;
	wire _w950_ ;
	wire _w949_ ;
	wire _w948_ ;
	wire _w947_ ;
	wire _w946_ ;
	wire _w945_ ;
	wire _w944_ ;
	wire _w943_ ;
	wire _w942_ ;
	wire _w941_ ;
	wire _w940_ ;
	wire _w939_ ;
	wire _w938_ ;
	wire _w937_ ;
	wire _w936_ ;
	wire _w935_ ;
	wire _w934_ ;
	wire _w933_ ;
	wire _w932_ ;
	wire _w931_ ;
	wire _w930_ ;
	wire _w929_ ;
	wire _w928_ ;
	wire _w927_ ;
	wire _w926_ ;
	wire _w925_ ;
	wire _w924_ ;
	wire _w923_ ;
	wire _w922_ ;
	wire _w921_ ;
	wire _w920_ ;
	wire _w919_ ;
	wire _w918_ ;
	wire _w917_ ;
	wire _w916_ ;
	wire _w915_ ;
	wire _w914_ ;
	wire _w913_ ;
	wire _w912_ ;
	wire _w911_ ;
	wire _w910_ ;
	wire _w909_ ;
	wire _w908_ ;
	wire _w907_ ;
	wire _w906_ ;
	wire _w905_ ;
	wire _w904_ ;
	wire _w903_ ;
	wire _w902_ ;
	wire _w901_ ;
	wire _w900_ ;
	wire _w899_ ;
	wire _w898_ ;
	wire _w897_ ;
	wire _w896_ ;
	wire _w895_ ;
	wire _w894_ ;
	wire _w893_ ;
	wire _w892_ ;
	wire _w891_ ;
	wire _w890_ ;
	wire _w889_ ;
	wire _w888_ ;
	wire _w887_ ;
	wire _w886_ ;
	wire _w885_ ;
	wire _w884_ ;
	wire _w883_ ;
	wire _w882_ ;
	wire _w881_ ;
	wire _w880_ ;
	wire _w879_ ;
	wire _w878_ ;
	wire _w877_ ;
	wire _w876_ ;
	wire _w875_ ;
	wire _w874_ ;
	wire _w873_ ;
	wire _w872_ ;
	wire _w871_ ;
	wire _w870_ ;
	wire _w869_ ;
	wire _w868_ ;
	wire _w867_ ;
	wire _w866_ ;
	wire _w865_ ;
	wire _w864_ ;
	wire _w863_ ;
	wire _w862_ ;
	wire _w861_ ;
	wire _w860_ ;
	wire _w859_ ;
	wire _w858_ ;
	wire _w857_ ;
	wire _w856_ ;
	wire _w855_ ;
	wire _w854_ ;
	wire _w853_ ;
	wire _w852_ ;
	wire _w851_ ;
	wire _w850_ ;
	wire _w849_ ;
	wire _w848_ ;
	wire _w847_ ;
	wire _w846_ ;
	wire _w845_ ;
	wire _w844_ ;
	wire _w843_ ;
	wire _w842_ ;
	wire _w841_ ;
	wire _w840_ ;
	wire _w839_ ;
	wire _w838_ ;
	wire _w837_ ;
	wire _w836_ ;
	wire _w835_ ;
	wire _w834_ ;
	wire _w833_ ;
	wire _w832_ ;
	wire _w831_ ;
	wire _w830_ ;
	wire _w829_ ;
	wire _w828_ ;
	wire _w827_ ;
	wire _w826_ ;
	wire _w825_ ;
	wire _w824_ ;
	wire _w823_ ;
	wire _w822_ ;
	wire _w821_ ;
	wire _w820_ ;
	wire _w819_ ;
	wire _w818_ ;
	wire _w817_ ;
	wire _w816_ ;
	wire _w815_ ;
	wire _w814_ ;
	wire _w813_ ;
	wire _w812_ ;
	wire _w811_ ;
	wire _w810_ ;
	wire _w809_ ;
	wire _w808_ ;
	wire _w807_ ;
	wire _w806_ ;
	wire _w805_ ;
	wire _w804_ ;
	wire _w803_ ;
	wire _w802_ ;
	wire _w801_ ;
	wire _w800_ ;
	wire _w799_ ;
	wire _w798_ ;
	wire _w797_ ;
	wire _w796_ ;
	wire _w795_ ;
	wire _w794_ ;
	wire _w793_ ;
	wire _w792_ ;
	wire _w791_ ;
	wire _w790_ ;
	wire _w789_ ;
	wire _w788_ ;
	wire _w787_ ;
	wire _w786_ ;
	wire _w785_ ;
	wire _w784_ ;
	wire _w783_ ;
	wire _w782_ ;
	wire _w781_ ;
	wire _w780_ ;
	wire _w779_ ;
	wire _w778_ ;
	wire _w777_ ;
	wire _w776_ ;
	wire _w775_ ;
	wire _w774_ ;
	wire _w773_ ;
	wire _w772_ ;
	wire _w771_ ;
	wire _w770_ ;
	wire _w769_ ;
	wire _w768_ ;
	wire _w767_ ;
	wire _w766_ ;
	wire _w765_ ;
	wire _w764_ ;
	wire _w763_ ;
	wire _w762_ ;
	wire _w761_ ;
	wire _w760_ ;
	wire _w759_ ;
	wire _w758_ ;
	wire _w757_ ;
	wire _w756_ ;
	wire _w755_ ;
	wire _w754_ ;
	wire _w753_ ;
	wire _w752_ ;
	wire _w751_ ;
	wire _w750_ ;
	wire _w749_ ;
	wire _w748_ ;
	wire _w747_ ;
	wire _w746_ ;
	wire _w745_ ;
	wire _w744_ ;
	wire _w743_ ;
	wire _w742_ ;
	wire _w741_ ;
	wire _w740_ ;
	wire _w739_ ;
	wire _w738_ ;
	wire _w737_ ;
	wire _w736_ ;
	wire _w735_ ;
	wire _w734_ ;
	wire _w733_ ;
	wire _w732_ ;
	wire _w731_ ;
	wire _w730_ ;
	wire _w729_ ;
	wire _w728_ ;
	wire _w727_ ;
	wire _w726_ ;
	wire _w725_ ;
	wire _w724_ ;
	wire _w723_ ;
	wire _w722_ ;
	wire _w721_ ;
	wire _w720_ ;
	wire _w719_ ;
	wire _w718_ ;
	wire _w717_ ;
	wire _w716_ ;
	wire _w715_ ;
	wire _w714_ ;
	wire _w713_ ;
	wire _w712_ ;
	wire _w711_ ;
	wire _w710_ ;
	wire _w709_ ;
	wire _w708_ ;
	wire _w707_ ;
	wire _w706_ ;
	wire _w705_ ;
	wire _w704_ ;
	wire _w703_ ;
	wire _w702_ ;
	wire _w701_ ;
	wire _w700_ ;
	wire _w699_ ;
	wire _w698_ ;
	wire _w697_ ;
	wire _w696_ ;
	wire _w695_ ;
	wire _w694_ ;
	wire _w693_ ;
	wire _w692_ ;
	wire _w691_ ;
	wire _w690_ ;
	wire _w689_ ;
	wire _w688_ ;
	wire _w687_ ;
	wire _w686_ ;
	wire _w685_ ;
	wire _w684_ ;
	wire _w683_ ;
	wire _w682_ ;
	wire _w681_ ;
	wire _w680_ ;
	wire _w679_ ;
	wire _w678_ ;
	wire _w677_ ;
	wire _w676_ ;
	wire _w675_ ;
	wire _w674_ ;
	wire _w673_ ;
	wire _w672_ ;
	wire _w671_ ;
	wire _w670_ ;
	wire _w669_ ;
	wire _w668_ ;
	wire _w667_ ;
	wire _w666_ ;
	wire _w665_ ;
	wire _w664_ ;
	wire _w663_ ;
	wire _w662_ ;
	wire _w661_ ;
	wire _w660_ ;
	wire _w659_ ;
	wire _w658_ ;
	wire _w657_ ;
	wire _w656_ ;
	wire _w655_ ;
	wire _w654_ ;
	wire _w653_ ;
	wire _w652_ ;
	wire _w651_ ;
	wire _w650_ ;
	wire _w649_ ;
	wire _w648_ ;
	wire _w647_ ;
	wire _w646_ ;
	wire _w645_ ;
	wire _w644_ ;
	wire _w643_ ;
	wire _w642_ ;
	wire _w641_ ;
	wire _w640_ ;
	wire _w639_ ;
	wire _w638_ ;
	wire _w637_ ;
	wire _w636_ ;
	wire _w635_ ;
	wire _w634_ ;
	wire _w633_ ;
	wire _w632_ ;
	wire _w631_ ;
	wire _w630_ ;
	wire _w629_ ;
	wire _w628_ ;
	wire _w627_ ;
	wire _w626_ ;
	wire _w625_ ;
	wire _w624_ ;
	wire _w623_ ;
	wire _w622_ ;
	wire _w621_ ;
	wire _w620_ ;
	wire _w619_ ;
	wire _w618_ ;
	wire _w617_ ;
	wire _w616_ ;
	wire _w615_ ;
	wire _w614_ ;
	wire _w613_ ;
	wire _w612_ ;
	wire _w611_ ;
	wire _w610_ ;
	wire _w609_ ;
	wire _w608_ ;
	wire _w607_ ;
	wire _w606_ ;
	wire _w605_ ;
	wire _w604_ ;
	wire _w603_ ;
	wire _w602_ ;
	wire _w601_ ;
	wire _w600_ ;
	wire _w599_ ;
	wire _w598_ ;
	wire _w597_ ;
	wire _w596_ ;
	wire _w595_ ;
	wire _w594_ ;
	wire _w593_ ;
	wire _w592_ ;
	wire _w591_ ;
	wire _w590_ ;
	wire _w589_ ;
	wire _w588_ ;
	wire _w587_ ;
	wire _w586_ ;
	wire _w585_ ;
	wire _w584_ ;
	wire _w583_ ;
	wire _w582_ ;
	wire _w581_ ;
	wire _w580_ ;
	wire _w579_ ;
	wire _w578_ ;
	wire _w577_ ;
	wire _w576_ ;
	wire _w575_ ;
	wire _w290_ ;
	wire _w289_ ;
	wire _w288_ ;
	wire _w287_ ;
	wire _w286_ ;
	wire _w285_ ;
	wire _w284_ ;
	wire _w283_ ;
	wire _w282_ ;
	wire _w281_ ;
	wire _w280_ ;
	wire _w279_ ;
	wire _w278_ ;
	wire _w277_ ;
	wire _w276_ ;
	wire _w275_ ;
	wire _w274_ ;
	wire _w273_ ;
	wire _w272_ ;
	wire _w271_ ;
	wire _w270_ ;
	wire _w269_ ;
	wire _w268_ ;
	wire _w267_ ;
	wire _w266_ ;
	wire _w265_ ;
	wire _w264_ ;
	wire _w263_ ;
	wire _w262_ ;
	wire _w261_ ;
	wire _w260_ ;
	wire _w259_ ;
	wire _w258_ ;
	wire _w257_ ;
	wire _w256_ ;
	wire _w255_ ;
	wire _w254_ ;
	wire _w253_ ;
	wire _w252_ ;
	wire _w251_ ;
	wire _w250_ ;
	wire _w249_ ;
	wire _w248_ ;
	wire _w247_ ;
	wire _w246_ ;
	wire _w245_ ;
	wire _w244_ ;
	wire _w243_ ;
	wire _w242_ ;
	wire _w241_ ;
	wire _w240_ ;
	wire _w239_ ;
	wire _w238_ ;
	wire _w237_ ;
	wire _w236_ ;
	wire _w235_ ;
	wire _w234_ ;
	wire _w233_ ;
	wire _w232_ ;
	wire _w231_ ;
	wire _w230_ ;
	wire _w229_ ;
	wire _w228_ ;
	wire _w227_ ;
	wire _w226_ ;
	wire _w225_ ;
	wire _w224_ ;
	wire _w223_ ;
	wire _w222_ ;
	wire _w221_ ;
	wire _w220_ ;
	wire _w219_ ;
	wire _w218_ ;
	wire _w217_ ;
	wire _w216_ ;
	wire _w215_ ;
	wire _w214_ ;
	wire _w213_ ;
	wire _w212_ ;
	wire _w211_ ;
	wire _w210_ ;
	wire _w209_ ;
	wire _w208_ ;
	wire _w207_ ;
	wire _w206_ ;
	wire _w205_ ;
	wire _w204_ ;
	wire _w203_ ;
	wire _w202_ ;
	wire _w201_ ;
	wire _w200_ ;
	wire _w199_ ;
	wire _w198_ ;
	wire _w197_ ;
	wire _w196_ ;
	wire _w195_ ;
	wire _w194_ ;
	wire _w193_ ;
	wire _w192_ ;
	wire _w191_ ;
	wire _w190_ ;
	wire _w189_ ;
	wire _w188_ ;
	wire _w187_ ;
	wire _w186_ ;
	wire _w185_ ;
	wire _w184_ ;
	wire _w183_ ;
	wire _w182_ ;
	wire _w181_ ;
	wire _w180_ ;
	wire _w179_ ;
	wire _w178_ ;
	wire _w177_ ;
	wire _w176_ ;
	wire _w175_ ;
	wire _w174_ ;
	wire _w173_ ;
	wire _w172_ ;
	wire _w171_ ;
	wire _w170_ ;
	wire _w169_ ;
	wire _w168_ ;
	wire _w167_ ;
	wire _w166_ ;
	wire _w165_ ;
	wire _w164_ ;
	wire _w163_ ;
	wire _w162_ ;
	wire _w161_ ;
	wire _w92_ ;
	wire _w91_ ;
	wire _w90_ ;
	wire _w89_ ;
	wire _w88_ ;
	wire _w87_ ;
	wire _w86_ ;
	wire _w85_ ;
	wire _w84_ ;
	wire _w83_ ;
	wire _w82_ ;
	wire _w81_ ;
	wire _w80_ ;
	wire _w79_ ;
	wire _w78_ ;
	wire _w77_ ;
	wire _w76_ ;
	wire _w75_ ;
	wire _w74_ ;
	wire _w73_ ;
	wire _w72_ ;
	wire _w71_ ;
	wire _w70_ ;
	wire _w69_ ;
	wire _w68_ ;
	wire _w67_ ;
	wire _w66_ ;
	wire _w65_ ;
	wire _w64_ ;
	wire _w63_ ;
	wire _w46_ ;
	wire _w45_ ;
	wire _w44_ ;
	wire _w43_ ;
	wire _w42_ ;
	wire _w41_ ;
	wire _w40_ ;
	wire _w39_ ;
	wire _w38_ ;
	wire _w37_ ;
	wire _w36_ ;
	wire _w35_ ;
	wire _w34_ ;
	wire _w47_ ;
	wire _w48_ ;
	wire _w49_ ;
	wire _w50_ ;
	wire _w51_ ;
	wire _w52_ ;
	wire _w53_ ;
	wire _w54_ ;
	wire _w55_ ;
	wire _w56_ ;
	wire _w57_ ;
	wire _w58_ ;
	wire _w59_ ;
	wire _w60_ ;
	wire _w61_ ;
	wire _w62_ ;
	wire _w93_ ;
	wire _w94_ ;
	wire _w95_ ;
	wire _w96_ ;
	wire _w97_ ;
	wire _w98_ ;
	wire _w99_ ;
	wire _w100_ ;
	wire _w101_ ;
	wire _w102_ ;
	wire _w103_ ;
	wire _w104_ ;
	wire _w105_ ;
	wire _w106_ ;
	wire _w107_ ;
	wire _w108_ ;
	wire _w109_ ;
	wire _w110_ ;
	wire _w111_ ;
	wire _w112_ ;
	wire _w113_ ;
	wire _w114_ ;
	wire _w115_ ;
	wire _w116_ ;
	wire _w117_ ;
	wire _w118_ ;
	wire _w119_ ;
	wire _w120_ ;
	wire _w121_ ;
	wire _w122_ ;
	wire _w123_ ;
	wire _w124_ ;
	wire _w125_ ;
	wire _w126_ ;
	wire _w127_ ;
	wire _w128_ ;
	wire _w129_ ;
	wire _w130_ ;
	wire _w131_ ;
	wire _w132_ ;
	wire _w133_ ;
	wire _w134_ ;
	wire _w135_ ;
	wire _w136_ ;
	wire _w137_ ;
	wire _w138_ ;
	wire _w139_ ;
	wire _w140_ ;
	wire _w141_ ;
	wire _w142_ ;
	wire _w143_ ;
	wire _w144_ ;
	wire _w145_ ;
	wire _w146_ ;
	wire _w147_ ;
	wire _w148_ ;
	wire _w149_ ;
	wire _w150_ ;
	wire _w151_ ;
	wire _w152_ ;
	wire _w153_ ;
	wire _w154_ ;
	wire _w155_ ;
	wire _w156_ ;
	wire _w157_ ;
	wire _w158_ ;
	wire _w159_ ;
	wire _w160_ ;
	wire _w291_ ;
	wire _w292_ ;
	wire _w293_ ;
	wire _w294_ ;
	wire _w295_ ;
	wire _w296_ ;
	wire _w297_ ;
	wire _w298_ ;
	wire _w299_ ;
	wire _w300_ ;
	wire _w301_ ;
	wire _w302_ ;
	wire _w303_ ;
	wire _w304_ ;
	wire _w305_ ;
	wire _w306_ ;
	wire _w307_ ;
	wire _w308_ ;
	wire _w309_ ;
	wire _w310_ ;
	wire _w311_ ;
	wire _w312_ ;
	wire _w313_ ;
	wire _w314_ ;
	wire _w315_ ;
	wire _w316_ ;
	wire _w317_ ;
	wire _w318_ ;
	wire _w319_ ;
	wire _w320_ ;
	wire _w321_ ;
	wire _w322_ ;
	wire _w323_ ;
	wire _w324_ ;
	wire _w325_ ;
	wire _w326_ ;
	wire _w327_ ;
	wire _w328_ ;
	wire _w329_ ;
	wire _w330_ ;
	wire _w331_ ;
	wire _w332_ ;
	wire _w333_ ;
	wire _w334_ ;
	wire _w335_ ;
	wire _w336_ ;
	wire _w337_ ;
	wire _w338_ ;
	wire _w339_ ;
	wire _w340_ ;
	wire _w341_ ;
	wire _w342_ ;
	wire _w343_ ;
	wire _w344_ ;
	wire _w345_ ;
	wire _w346_ ;
	wire _w347_ ;
	wire _w348_ ;
	wire _w349_ ;
	wire _w350_ ;
	wire _w351_ ;
	wire _w352_ ;
	wire _w353_ ;
	wire _w354_ ;
	wire _w355_ ;
	wire _w356_ ;
	wire _w357_ ;
	wire _w358_ ;
	wire _w359_ ;
	wire _w360_ ;
	wire _w361_ ;
	wire _w362_ ;
	wire _w363_ ;
	wire _w364_ ;
	wire _w365_ ;
	wire _w366_ ;
	wire _w367_ ;
	wire _w368_ ;
	wire _w369_ ;
	wire _w370_ ;
	wire _w371_ ;
	wire _w372_ ;
	wire _w373_ ;
	wire _w374_ ;
	wire _w375_ ;
	wire _w376_ ;
	wire _w377_ ;
	wire _w378_ ;
	wire _w379_ ;
	wire _w380_ ;
	wire _w381_ ;
	wire _w382_ ;
	wire _w383_ ;
	wire _w384_ ;
	wire _w385_ ;
	wire _w386_ ;
	wire _w387_ ;
	wire _w388_ ;
	wire _w389_ ;
	wire _w390_ ;
	wire _w391_ ;
	wire _w392_ ;
	wire _w393_ ;
	wire _w394_ ;
	wire _w395_ ;
	wire _w396_ ;
	wire _w397_ ;
	wire _w398_ ;
	wire _w399_ ;
	wire _w400_ ;
	wire _w401_ ;
	wire _w402_ ;
	wire _w403_ ;
	wire _w404_ ;
	wire _w405_ ;
	wire _w406_ ;
	wire _w407_ ;
	wire _w408_ ;
	wire _w409_ ;
	wire _w410_ ;
	wire _w411_ ;
	wire _w412_ ;
	wire _w413_ ;
	wire _w414_ ;
	wire _w415_ ;
	wire _w416_ ;
	wire _w417_ ;
	wire _w418_ ;
	wire _w419_ ;
	wire _w420_ ;
	wire _w421_ ;
	wire _w422_ ;
	wire _w423_ ;
	wire _w424_ ;
	wire _w425_ ;
	wire _w426_ ;
	wire _w427_ ;
	wire _w428_ ;
	wire _w429_ ;
	wire _w430_ ;
	wire _w431_ ;
	wire _w432_ ;
	wire _w433_ ;
	wire _w434_ ;
	wire _w435_ ;
	wire _w436_ ;
	wire _w437_ ;
	wire _w438_ ;
	wire _w439_ ;
	wire _w440_ ;
	wire _w441_ ;
	wire _w442_ ;
	wire _w443_ ;
	wire _w444_ ;
	wire _w445_ ;
	wire _w446_ ;
	wire _w447_ ;
	wire _w448_ ;
	wire _w449_ ;
	wire _w450_ ;
	wire _w451_ ;
	wire _w452_ ;
	wire _w453_ ;
	wire _w454_ ;
	wire _w455_ ;
	wire _w456_ ;
	wire _w457_ ;
	wire _w458_ ;
	wire _w459_ ;
	wire _w460_ ;
	wire _w461_ ;
	wire _w462_ ;
	wire _w463_ ;
	wire _w464_ ;
	wire _w465_ ;
	wire _w466_ ;
	wire _w467_ ;
	wire _w468_ ;
	wire _w469_ ;
	wire _w470_ ;
	wire _w471_ ;
	wire _w472_ ;
	wire _w473_ ;
	wire _w474_ ;
	wire _w475_ ;
	wire _w476_ ;
	wire _w477_ ;
	wire _w478_ ;
	wire _w479_ ;
	wire _w480_ ;
	wire _w481_ ;
	wire _w482_ ;
	wire _w483_ ;
	wire _w484_ ;
	wire _w485_ ;
	wire _w486_ ;
	wire _w487_ ;
	wire _w488_ ;
	wire _w489_ ;
	wire _w490_ ;
	wire _w491_ ;
	wire _w492_ ;
	wire _w493_ ;
	wire _w494_ ;
	wire _w495_ ;
	wire _w496_ ;
	wire _w497_ ;
	wire _w498_ ;
	wire _w499_ ;
	wire _w500_ ;
	wire _w501_ ;
	wire _w502_ ;
	wire _w503_ ;
	wire _w504_ ;
	wire _w505_ ;
	wire _w506_ ;
	wire _w507_ ;
	wire _w508_ ;
	wire _w509_ ;
	wire _w510_ ;
	wire _w511_ ;
	wire _w512_ ;
	wire _w513_ ;
	wire _w514_ ;
	wire _w515_ ;
	wire _w516_ ;
	wire _w517_ ;
	wire _w518_ ;
	wire _w519_ ;
	wire _w520_ ;
	wire _w521_ ;
	wire _w522_ ;
	wire _w523_ ;
	wire _w524_ ;
	wire _w525_ ;
	wire _w526_ ;
	wire _w527_ ;
	wire _w528_ ;
	wire _w529_ ;
	wire _w530_ ;
	wire _w531_ ;
	wire _w532_ ;
	wire _w533_ ;
	wire _w534_ ;
	wire _w535_ ;
	wire _w536_ ;
	wire _w537_ ;
	wire _w538_ ;
	wire _w539_ ;
	wire _w540_ ;
	wire _w541_ ;
	wire _w542_ ;
	wire _w543_ ;
	wire _w544_ ;
	wire _w545_ ;
	wire _w546_ ;
	wire _w547_ ;
	wire _w548_ ;
	wire _w549_ ;
	wire _w550_ ;
	wire _w551_ ;
	wire _w552_ ;
	wire _w553_ ;
	wire _w554_ ;
	wire _w555_ ;
	wire _w556_ ;
	wire _w557_ ;
	wire _w558_ ;
	wire _w559_ ;
	wire _w560_ ;
	wire _w561_ ;
	wire _w562_ ;
	wire _w563_ ;
	wire _w564_ ;
	wire _w565_ ;
	wire _w566_ ;
	wire _w567_ ;
	wire _w568_ ;
	wire _w569_ ;
	wire _w570_ ;
	wire _w571_ ;
	wire _w572_ ;
	wire _w573_ ;
	wire _w574_ ;
	wire _w1143_ ;
	wire _w1144_ ;
	wire _w1145_ ;
	wire _w1146_ ;
	wire _w1147_ ;
	wire _w1148_ ;
	wire _w1149_ ;
	wire _w1150_ ;
	wire _w1151_ ;
	wire _w1152_ ;
	wire _w1153_ ;
	wire _w1154_ ;
	wire _w1155_ ;
	wire _w1156_ ;
	wire _w1157_ ;
	wire _w1158_ ;
	wire _w1159_ ;
	wire _w1160_ ;
	wire _w1161_ ;
	wire _w1162_ ;
	wire _w1163_ ;
	wire _w1164_ ;
	wire _w1165_ ;
	wire _w1166_ ;
	wire _w1167_ ;
	wire _w1168_ ;
	wire _w1169_ ;
	wire _w1170_ ;
	wire _w1171_ ;
	wire _w1172_ ;
	wire _w1173_ ;
	wire _w1174_ ;
	wire _w1175_ ;
	wire _w1176_ ;
	wire _w1177_ ;
	wire _w1178_ ;
	wire _w1179_ ;
	wire _w1180_ ;
	wire _w1181_ ;
	wire _w1182_ ;
	wire _w1183_ ;
	wire _w1184_ ;
	wire _w1185_ ;
	wire _w1186_ ;
	wire _w1187_ ;
	wire _w1188_ ;
	wire _w1189_ ;
	wire _w1190_ ;
	wire _w1191_ ;
	wire _w1192_ ;
	wire _w1193_ ;
	wire _w1194_ ;
	wire _w1195_ ;
	wire _w1196_ ;
	wire _w1197_ ;
	wire _w1198_ ;
	wire _w1199_ ;
	wire _w1200_ ;
	wire _w1201_ ;
	wire _w1202_ ;
	wire _w1203_ ;
	wire _w1204_ ;
	wire _w1205_ ;
	wire _w1206_ ;
	wire _w1207_ ;
	wire _w1208_ ;
	wire _w1209_ ;
	wire _w1210_ ;
	wire _w1211_ ;
	wire _w1212_ ;
	wire _w1213_ ;
	wire _w1214_ ;
	wire _w1215_ ;
	wire _w1216_ ;
	wire _w1217_ ;
	wire _w1218_ ;
	wire _w1219_ ;
	wire _w1220_ ;
	wire _w1221_ ;
	wire _w1222_ ;
	wire _w1223_ ;
	wire _w1224_ ;
	wire _w1225_ ;
	wire _w1226_ ;
	wire _w1227_ ;
	wire _w1228_ ;
	wire _w1229_ ;
	wire _w1230_ ;
	wire _w1231_ ;
	wire _w1232_ ;
	wire _w1233_ ;
	wire _w1234_ ;
	wire _w1235_ ;
	wire _w1236_ ;
	wire _w1237_ ;
	wire _w1238_ ;
	wire _w1239_ ;
	wire _w1240_ ;
	wire _w1241_ ;
	wire _w1242_ ;
	wire _w1243_ ;
	wire _w1244_ ;
	wire _w1245_ ;
	wire _w1246_ ;
	wire _w1247_ ;
	wire _w1248_ ;
	wire _w1249_ ;
	wire _w1250_ ;
	wire _w1251_ ;
	wire _w1252_ ;
	wire _w1253_ ;
	wire _w1254_ ;
	wire _w1255_ ;
	wire _w1256_ ;
	wire _w1257_ ;
	wire _w1258_ ;
	wire _w1259_ ;
	wire _w1260_ ;
	wire _w1261_ ;
	wire _w1262_ ;
	wire _w1263_ ;
	wire _w1264_ ;
	wire _w1265_ ;
	wire _w1266_ ;
	wire _w1267_ ;
	wire _w1268_ ;
	wire _w1269_ ;
	wire _w1270_ ;
	wire _w1271_ ;
	wire _w1272_ ;
	wire _w1273_ ;
	wire _w1274_ ;
	wire _w1275_ ;
	wire _w1276_ ;
	wire _w1277_ ;
	wire _w1278_ ;
	wire _w1279_ ;
	wire _w1280_ ;
	wire _w1281_ ;
	wire _w1282_ ;
	wire _w1283_ ;
	wire _w1284_ ;
	wire _w1285_ ;
	wire _w1286_ ;
	wire _w1287_ ;
	wire _w1288_ ;
	wire _w1289_ ;
	wire _w1290_ ;
	wire _w1291_ ;
	wire _w1292_ ;
	wire _w1293_ ;
	wire _w1294_ ;
	wire _w1295_ ;
	wire _w1296_ ;
	wire _w1297_ ;
	wire _w1298_ ;
	wire _w1299_ ;
	wire _w1300_ ;
	wire _w1301_ ;
	wire _w1302_ ;
	wire _w1303_ ;
	wire _w1304_ ;
	wire _w1305_ ;
	wire _w1306_ ;
	wire _w1307_ ;
	wire _w1308_ ;
	wire _w1309_ ;
	wire _w1310_ ;
	wire _w1311_ ;
	wire _w1312_ ;
	wire _w1313_ ;
	wire _w1314_ ;
	wire _w1315_ ;
	wire _w1316_ ;
	wire _w1317_ ;
	wire _w1318_ ;
	wire _w1319_ ;
	wire _w1320_ ;
	wire _w1321_ ;
	wire _w1322_ ;
	wire _w1323_ ;
	wire _w1324_ ;
	wire _w1325_ ;
	wire _w1326_ ;
	wire _w1327_ ;
	wire _w1328_ ;
	wire _w1329_ ;
	wire _w1330_ ;
	wire _w1331_ ;
	wire _w1332_ ;
	wire _w1333_ ;
	wire _w1334_ ;
	wire _w1335_ ;
	wire _w1336_ ;
	wire _w1337_ ;
	wire _w1338_ ;
	wire _w1339_ ;
	wire _w1340_ ;
	wire _w1341_ ;
	wire _w1342_ ;
	wire _w1343_ ;
	wire _w1344_ ;
	wire _w1345_ ;
	wire _w1346_ ;
	wire _w1347_ ;
	wire _w1348_ ;
	wire _w1349_ ;
	wire _w1350_ ;
	wire _w1351_ ;
	wire _w1352_ ;
	wire _w1353_ ;
	wire _w1354_ ;
	wire _w1355_ ;
	wire _w1356_ ;
	wire _w1357_ ;
	wire _w1358_ ;
	wire _w1359_ ;
	wire _w1360_ ;
	wire _w1361_ ;
	wire _w1362_ ;
	wire _w1363_ ;
	wire _w1364_ ;
	wire _w1365_ ;
	wire _w1366_ ;
	wire _w1367_ ;
	wire _w1368_ ;
	wire _w1369_ ;
	wire _w1370_ ;
	wire _w1371_ ;
	wire _w1372_ ;
	wire _w1373_ ;
	wire _w1374_ ;
	wire _w1375_ ;
	wire _w1376_ ;
	wire _w1377_ ;
	wire _w1378_ ;
	wire _w1379_ ;
	wire _w1380_ ;
	wire _w1381_ ;
	wire _w1382_ ;
	wire _w1383_ ;
	wire _w1384_ ;
	wire _w1385_ ;
	wire _w1386_ ;
	wire _w1387_ ;
	wire _w1388_ ;
	wire _w1389_ ;
	wire _w1390_ ;
	wire _w1391_ ;
	wire _w1392_ ;
	wire _w1393_ ;
	wire _w1394_ ;
	wire _w1395_ ;
	wire _w1396_ ;
	wire _w1397_ ;
	wire _w1398_ ;
	wire _w1399_ ;
	wire _w1400_ ;
	wire _w1401_ ;
	wire _w1402_ ;
	wire _w1403_ ;
	wire _w1404_ ;
	wire _w1405_ ;
	wire _w1406_ ;
	wire _w1407_ ;
	wire _w1408_ ;
	wire _w1409_ ;
	wire _w1410_ ;
	wire _w1411_ ;
	wire _w1412_ ;
	wire _w1413_ ;
	wire _w1414_ ;
	wire _w1415_ ;
	wire _w1416_ ;
	wire _w1417_ ;
	wire _w1418_ ;
	wire _w1419_ ;
	wire _w1420_ ;
	wire _w1421_ ;
	wire _w1422_ ;
	wire _w1423_ ;
	wire _w1424_ ;
	wire _w1425_ ;
	wire _w1426_ ;
	wire _w1427_ ;
	wire _w1428_ ;
	wire _w1429_ ;
	wire _w1430_ ;
	wire _w1431_ ;
	wire _w1432_ ;
	wire _w1433_ ;
	wire _w1434_ ;
	wire _w1435_ ;
	wire _w1436_ ;
	wire _w1437_ ;
	wire _w1438_ ;
	wire _w1439_ ;
	wire _w1440_ ;
	wire _w1441_ ;
	wire _w1442_ ;
	wire _w1443_ ;
	wire _w1444_ ;
	wire _w1445_ ;
	wire _w1446_ ;
	wire _w1447_ ;
	wire _w1448_ ;
	wire _w1449_ ;
	wire _w1450_ ;
	wire _w1451_ ;
	wire _w1452_ ;
	wire _w1453_ ;
	wire _w1454_ ;
	wire _w1455_ ;
	wire _w1456_ ;
	wire _w1457_ ;
	wire _w1458_ ;
	wire _w1459_ ;
	wire _w1460_ ;
	wire _w1461_ ;
	wire _w1462_ ;
	wire _w1463_ ;
	wire _w1464_ ;
	wire _w1465_ ;
	wire _w1466_ ;
	wire _w1467_ ;
	wire _w1468_ ;
	wire _w1469_ ;
	wire _w1470_ ;
	wire _w1471_ ;
	wire _w1472_ ;
	wire _w1473_ ;
	wire _w1474_ ;
	wire _w1475_ ;
	wire _w1476_ ;
	wire _w1477_ ;
	wire _w1478_ ;
	wire _w1479_ ;
	wire _w1480_ ;
	wire _w1481_ ;
	wire _w1482_ ;
	wire _w1483_ ;
	wire _w1484_ ;
	wire _w1485_ ;
	wire _w1486_ ;
	wire _w1487_ ;
	wire _w1488_ ;
	wire _w1489_ ;
	wire _w1490_ ;
	wire _w1491_ ;
	wire _w1492_ ;
	wire _w1493_ ;
	wire _w1494_ ;
	wire _w1495_ ;
	wire _w1496_ ;
	wire _w1497_ ;
	wire _w1498_ ;
	wire _w1499_ ;
	wire _w1500_ ;
	wire _w1501_ ;
	wire _w1502_ ;
	wire _w1503_ ;
	wire _w1504_ ;
	wire _w1505_ ;
	wire _w1506_ ;
	wire _w1507_ ;
	wire _w1508_ ;
	wire _w1509_ ;
	wire _w1510_ ;
	wire _w1511_ ;
	wire _w1512_ ;
	wire _w1513_ ;
	wire _w1514_ ;
	wire _w1515_ ;
	wire _w1516_ ;
	wire _w1517_ ;
	wire _w1518_ ;
	wire _w1519_ ;
	wire _w1520_ ;
	wire _w1521_ ;
	wire _w1522_ ;
	wire _w1523_ ;
	wire _w1524_ ;
	wire _w1525_ ;
	wire _w1526_ ;
	wire _w1527_ ;
	wire _w1528_ ;
	wire _w1529_ ;
	wire _w1530_ ;
	wire _w1531_ ;
	wire _w1532_ ;
	wire _w1533_ ;
	wire _w1534_ ;
	wire _w1535_ ;
	wire _w1536_ ;
	wire _w1537_ ;
	wire _w1538_ ;
	wire _w1539_ ;
	wire _w1540_ ;
	wire _w1541_ ;
	wire _w1542_ ;
	wire _w1543_ ;
	wire _w1544_ ;
	wire _w1545_ ;
	wire _w1546_ ;
	wire _w1547_ ;
	wire _w1548_ ;
	wire _w1549_ ;
	wire _w1550_ ;
	wire _w1551_ ;
	wire _w1552_ ;
	wire _w1553_ ;
	wire _w1554_ ;
	wire _w1555_ ;
	wire _w1556_ ;
	wire _w1557_ ;
	wire _w1558_ ;
	wire _w1559_ ;
	wire _w1560_ ;
	wire _w1561_ ;
	wire _w1562_ ;
	wire _w1563_ ;
	wire _w1564_ ;
	wire _w1565_ ;
	wire _w1566_ ;
	wire _w1567_ ;
	wire _w1568_ ;
	wire _w1569_ ;
	wire _w1570_ ;
	wire _w1571_ ;
	wire _w1572_ ;
	wire _w1573_ ;
	wire _w1574_ ;
	wire _w1575_ ;
	wire _w1576_ ;
	wire _w1577_ ;
	wire _w1578_ ;
	wire _w1579_ ;
	wire _w1580_ ;
	wire _w1581_ ;
	wire _w1582_ ;
	wire _w1583_ ;
	wire _w1584_ ;
	wire _w1585_ ;
	wire _w1586_ ;
	wire _w1587_ ;
	wire _w1588_ ;
	wire _w1589_ ;
	wire _w1590_ ;
	wire _w1591_ ;
	wire _w1592_ ;
	wire _w1593_ ;
	wire _w1594_ ;
	wire _w1595_ ;
	wire _w1596_ ;
	wire _w1597_ ;
	wire _w1598_ ;
	wire _w1599_ ;
	wire _w1600_ ;
	wire _w1601_ ;
	wire _w1602_ ;
	wire _w1603_ ;
	wire _w1604_ ;
	wire _w1605_ ;
	wire _w1606_ ;
	wire _w1607_ ;
	wire _w1608_ ;
	wire _w1609_ ;
	wire _w1610_ ;
	wire _w1611_ ;
	wire _w1612_ ;
	wire _w1613_ ;
	wire _w1614_ ;
	wire _w1615_ ;
	wire _w1616_ ;
	wire _w1617_ ;
	wire _w1618_ ;
	wire _w1619_ ;
	wire _w1620_ ;
	wire _w1621_ ;
	wire _w1622_ ;
	wire _w1623_ ;
	wire _w1624_ ;
	wire _w1625_ ;
	wire _w1626_ ;
	wire _w1627_ ;
	wire _w1628_ ;
	wire _w1629_ ;
	wire _w1630_ ;
	wire _w1631_ ;
	wire _w1632_ ;
	wire _w1633_ ;
	wire _w1634_ ;
	wire _w1635_ ;
	wire _w1636_ ;
	wire _w1637_ ;
	wire _w1638_ ;
	wire _w1639_ ;
	wire _w1640_ ;
	wire _w1641_ ;
	wire _w1642_ ;
	wire _w1643_ ;
	wire _w1644_ ;
	wire _w1645_ ;
	wire _w1646_ ;
	wire _w1647_ ;
	wire _w1648_ ;
	wire _w1649_ ;
	wire _w1650_ ;
	wire _w1651_ ;
	wire _w1652_ ;
	wire _w1653_ ;
	wire _w1654_ ;
	wire _w1655_ ;
	wire _w1656_ ;
	wire _w1657_ ;
	wire _w1658_ ;
	wire _w1659_ ;
	wire _w1660_ ;
	wire _w1661_ ;
	wire _w1662_ ;
	wire _w1663_ ;
	wire _w1664_ ;
	wire _w1665_ ;
	wire _w1666_ ;
	wire _w1667_ ;
	wire _w1668_ ;
	wire _w1669_ ;
	wire _w1670_ ;
	wire _w1671_ ;
	wire _w1672_ ;
	wire _w1673_ ;
	wire _w1674_ ;
	wire _w1675_ ;
	wire _w1676_ ;
	wire _w1677_ ;
	wire _w1678_ ;
	wire _w1679_ ;
	wire _w1680_ ;
	wire _w1681_ ;
	wire _w1682_ ;
	wire _w1683_ ;
	wire _w1684_ ;
	wire _w1685_ ;
	wire _w1686_ ;
	wire _w1687_ ;
	wire _w1688_ ;
	wire _w1689_ ;
	wire _w1690_ ;
	wire _w1691_ ;
	wire _w1692_ ;
	wire _w1693_ ;
	wire _w1694_ ;
	wire _w1695_ ;
	wire _w1696_ ;
	wire _w1697_ ;
	wire _w1698_ ;
	wire _w1699_ ;
	wire _w1700_ ;
	wire _w1701_ ;
	wire _w1702_ ;
	wire _w1703_ ;
	wire _w1704_ ;
	wire _w1705_ ;
	wire _w1706_ ;
	wire _w1707_ ;
	wire _w1708_ ;
	wire _w1709_ ;
	wire _w1710_ ;
	wire _w1711_ ;
	wire _w1712_ ;
	wire _w1713_ ;
	wire _w1714_ ;
	wire _w1715_ ;
	wire _w1716_ ;
	wire _w1717_ ;
	wire _w1718_ ;
	wire _w1719_ ;
	wire _w1720_ ;
	wire _w1721_ ;
	wire _w1722_ ;
	wire _w1723_ ;
	wire _w1724_ ;
	wire _w1725_ ;
	wire _w1726_ ;
	wire _w1727_ ;
	wire _w1728_ ;
	wire _w1729_ ;
	wire _w1730_ ;
	wire _w1731_ ;
	wire _w1732_ ;
	wire _w1733_ ;
	wire _w1734_ ;
	wire _w1735_ ;
	wire _w1736_ ;
	wire _w1737_ ;
	wire _w1738_ ;
	wire _w1739_ ;
	wire _w1740_ ;
	wire _w1741_ ;
	wire _w1742_ ;
	wire _w1743_ ;
	wire _w1744_ ;
	wire _w1745_ ;
	wire _w1746_ ;
	wire _w1747_ ;
	wire _w1748_ ;
	wire _w1749_ ;
	wire _w1750_ ;
	wire _w1751_ ;
	wire _w1752_ ;
	wire _w1753_ ;
	wire _w1754_ ;
	wire _w1755_ ;
	wire _w1756_ ;
	wire _w1757_ ;
	wire _w1758_ ;
	wire _w1759_ ;
	wire _w1760_ ;
	wire _w1761_ ;
	wire _w1762_ ;
	wire _w1763_ ;
	wire _w1764_ ;
	wire _w1765_ ;
	wire _w1766_ ;
	wire _w1767_ ;
	wire _w1768_ ;
	wire _w1769_ ;
	wire _w1770_ ;
	wire _w1771_ ;
	wire _w1772_ ;
	wire _w1773_ ;
	wire _w1774_ ;
	wire _w1775_ ;
	wire _w1776_ ;
	wire _w1777_ ;
	wire _w1778_ ;
	wire _w1779_ ;
	wire _w1780_ ;
	wire _w1781_ ;
	wire _w1782_ ;
	wire _w1783_ ;
	wire _w1784_ ;
	wire _w1785_ ;
	wire _w1786_ ;
	wire _w1787_ ;
	wire _w1788_ ;
	wire _w1789_ ;
	wire _w1790_ ;
	wire _w1791_ ;
	wire _w1792_ ;
	wire _w1793_ ;
	wire _w1794_ ;
	wire _w1795_ ;
	wire _w1796_ ;
	wire _w1797_ ;
	wire _w1798_ ;
	wire _w1799_ ;
	wire _w1800_ ;
	wire _w1801_ ;
	wire _w1802_ ;
	wire _w1803_ ;
	wire _w1804_ ;
	wire _w1805_ ;
	wire _w1806_ ;
	wire _w1807_ ;
	wire _w1808_ ;
	wire _w1809_ ;
	wire _w1810_ ;
	wire _w1811_ ;
	wire _w1812_ ;
	wire _w1813_ ;
	wire _w1814_ ;
	wire _w1815_ ;
	wire _w1816_ ;
	wire _w1817_ ;
	wire _w1818_ ;
	wire _w1819_ ;
	wire _w1820_ ;
	wire _w1821_ ;
	wire _w1822_ ;
	wire _w1823_ ;
	wire _w1824_ ;
	wire _w1825_ ;
	wire _w1826_ ;
	wire _w1827_ ;
	wire _w1828_ ;
	wire _w1829_ ;
	wire _w1830_ ;
	wire _w1831_ ;
	wire _w1832_ ;
	wire _w1833_ ;
	wire _w1834_ ;
	wire _w1835_ ;
	wire _w1836_ ;
	wire _w1837_ ;
	wire _w1838_ ;
	wire _w1839_ ;
	wire _w1840_ ;
	wire _w1841_ ;
	wire _w1842_ ;
	wire _w1843_ ;
	wire _w1844_ ;
	wire _w1845_ ;
	wire _w1846_ ;
	wire _w1847_ ;
	wire _w1848_ ;
	wire _w1849_ ;
	wire _w1850_ ;
	wire _w1851_ ;
	wire _w1852_ ;
	wire _w1853_ ;
	wire _w1854_ ;
	wire _w1855_ ;
	wire _w1856_ ;
	wire _w1857_ ;
	wire _w1858_ ;
	wire _w1859_ ;
	wire _w1860_ ;
	wire _w1861_ ;
	wire _w1862_ ;
	wire _w1863_ ;
	wire _w1864_ ;
	wire _w1865_ ;
	wire _w1866_ ;
	wire _w1867_ ;
	wire _w1868_ ;
	wire _w1869_ ;
	wire _w1870_ ;
	wire _w1871_ ;
	wire _w1872_ ;
	wire _w1873_ ;
	wire _w1874_ ;
	wire _w1875_ ;
	wire _w1876_ ;
	wire _w1877_ ;
	wire _w1878_ ;
	wire _w1879_ ;
	wire _w1880_ ;
	wire _w1881_ ;
	wire _w1882_ ;
	wire _w1883_ ;
	wire _w1884_ ;
	wire _w1885_ ;
	wire _w1886_ ;
	wire _w1887_ ;
	wire _w1888_ ;
	wire _w1889_ ;
	wire _w1890_ ;
	wire _w1891_ ;
	wire _w1892_ ;
	wire _w1893_ ;
	wire _w1894_ ;
	wire _w1895_ ;
	wire _w1896_ ;
	wire _w1897_ ;
	wire _w1898_ ;
	wire _w1899_ ;
	wire _w1900_ ;
	wire _w1901_ ;
	wire _w1902_ ;
	wire _w1903_ ;
	wire _w1904_ ;
	wire _w1905_ ;
	wire _w1906_ ;
	wire _w1907_ ;
	wire _w1908_ ;
	wire _w1909_ ;
	wire _w1910_ ;
	wire _w1911_ ;
	wire _w1912_ ;
	wire _w1913_ ;
	wire _w1914_ ;
	wire _w1915_ ;
	wire _w1916_ ;
	wire _w1917_ ;
	wire _w1918_ ;
	wire _w1919_ ;
	wire _w1920_ ;
	wire _w1921_ ;
	wire _w1922_ ;
	wire _w1923_ ;
	wire _w1924_ ;
	wire _w1925_ ;
	wire _w1926_ ;
	wire _w1927_ ;
	wire _w1928_ ;
	wire _w1929_ ;
	wire _w1930_ ;
	wire _w1931_ ;
	wire _w1932_ ;
	wire _w1933_ ;
	wire _w1934_ ;
	wire _w1935_ ;
	wire _w1936_ ;
	wire _w1937_ ;
	wire _w1938_ ;
	wire _w1939_ ;
	wire _w1940_ ;
	wire _w1941_ ;
	wire _w1942_ ;
	wire _w1943_ ;
	wire _w1944_ ;
	wire _w1945_ ;
	wire _w1946_ ;
	wire _w1947_ ;
	wire _w1948_ ;
	wire _w1949_ ;
	wire _w1950_ ;
	wire _w1951_ ;
	wire _w1952_ ;
	wire _w1953_ ;
	wire _w1954_ ;
	wire _w1955_ ;
	wire _w1956_ ;
	wire _w1957_ ;
	wire _w1958_ ;
	wire _w1959_ ;
	wire _w1960_ ;
	wire _w1961_ ;
	wire _w1962_ ;
	wire _w1963_ ;
	wire _w1964_ ;
	wire _w1965_ ;
	wire _w1966_ ;
	wire _w1967_ ;
	wire _w1968_ ;
	wire _w1969_ ;
	wire _w1970_ ;
	wire _w1971_ ;
	wire _w1972_ ;
	wire _w1973_ ;
	wire _w1974_ ;
	wire _w1975_ ;
	wire _w1976_ ;
	wire _w1977_ ;
	wire _w1978_ ;
	wire _w1979_ ;
	wire _w1980_ ;
	wire _w1981_ ;
	wire _w1982_ ;
	wire _w1983_ ;
	wire _w1984_ ;
	wire _w1985_ ;
	wire _w1986_ ;
	wire _w1987_ ;
	wire _w1988_ ;
	wire _w1989_ ;
	wire _w1990_ ;
	wire _w1991_ ;
	wire _w1992_ ;
	wire _w1993_ ;
	wire _w1994_ ;
	wire _w1995_ ;
	wire _w1996_ ;
	wire _w1997_ ;
	wire _w1998_ ;
	wire _w1999_ ;
	wire _w2000_ ;
	wire _w2001_ ;
	wire _w2002_ ;
	wire _w2003_ ;
	wire _w2004_ ;
	wire _w2005_ ;
	wire _w2006_ ;
	wire _w2007_ ;
	wire _w2008_ ;
	wire _w2009_ ;
	wire _w2010_ ;
	wire _w2011_ ;
	wire _w2012_ ;
	wire _w2013_ ;
	wire _w2014_ ;
	wire _w2015_ ;
	wire _w2016_ ;
	wire _w2017_ ;
	wire _w2018_ ;
	wire _w2019_ ;
	wire _w2020_ ;
	wire _w2021_ ;
	wire _w2022_ ;
	wire _w2023_ ;
	wire _w2024_ ;
	wire _w2025_ ;
	wire _w2026_ ;
	wire _w2027_ ;
	wire _w2028_ ;
	wire _w2029_ ;
	wire _w2030_ ;
	wire _w2031_ ;
	wire _w2032_ ;
	wire _w2033_ ;
	wire _w2034_ ;
	wire _w2035_ ;
	wire _w2036_ ;
	wire _w2037_ ;
	wire _w2038_ ;
	wire _w2039_ ;
	wire _w2040_ ;
	wire _w2041_ ;
	wire _w2042_ ;
	wire _w2043_ ;
	wire _w2044_ ;
	wire _w2045_ ;
	wire _w2046_ ;
	wire _w2047_ ;
	wire _w2048_ ;
	wire _w2049_ ;
	wire _w2050_ ;
	wire _w2051_ ;
	wire _w2052_ ;
	wire _w2053_ ;
	wire _w2054_ ;
	wire _w2055_ ;
	wire _w2056_ ;
	wire _w2057_ ;
	wire _w2058_ ;
	wire _w2059_ ;
	wire _w2060_ ;
	wire _w2061_ ;
	wire _w2062_ ;
	wire _w2063_ ;
	wire _w2064_ ;
	wire _w2065_ ;
	wire _w2066_ ;
	wire _w2067_ ;
	wire _w2068_ ;
	wire _w2069_ ;
	wire _w2070_ ;
	wire _w2071_ ;
	wire _w2072_ ;
	wire _w2073_ ;
	wire _w2074_ ;
	wire _w2075_ ;
	wire _w2076_ ;
	wire _w2077_ ;
	wire _w2078_ ;
	wire _w2079_ ;
	wire _w2080_ ;
	wire _w2081_ ;
	wire _w2082_ ;
	wire _w2083_ ;
	wire _w2084_ ;
	wire _w2085_ ;
	wire _w2086_ ;
	wire _w2087_ ;
	wire _w2088_ ;
	wire _w2089_ ;
	wire _w2090_ ;
	wire _w2091_ ;
	wire _w2092_ ;
	wire _w2093_ ;
	wire _w2094_ ;
	wire _w2095_ ;
	wire _w2096_ ;
	wire _w2097_ ;
	wire _w2098_ ;
	wire _w2099_ ;
	wire _w2100_ ;
	wire _w2101_ ;
	wire _w2102_ ;
	wire _w2103_ ;
	wire _w2104_ ;
	wire _w2105_ ;
	wire _w2106_ ;
	wire _w2107_ ;
	wire _w2108_ ;
	wire _w2109_ ;
	wire _w2110_ ;
	wire _w2111_ ;
	wire _w2112_ ;
	wire _w2113_ ;
	wire _w2114_ ;
	wire _w2115_ ;
	wire _w2116_ ;
	wire _w2117_ ;
	wire _w2118_ ;
	wire _w2119_ ;
	wire _w2120_ ;
	wire _w2121_ ;
	wire _w2122_ ;
	wire _w2123_ ;
	wire _w2124_ ;
	wire _w2125_ ;
	wire _w2126_ ;
	wire _w2127_ ;
	wire _w2128_ ;
	wire _w2129_ ;
	wire _w2130_ ;
	wire _w2131_ ;
	wire _w2132_ ;
	wire _w2133_ ;
	wire _w2134_ ;
	wire _w2135_ ;
	wire _w2136_ ;
	wire _w2137_ ;
	wire _w2138_ ;
	wire _w2139_ ;
	wire _w2140_ ;
	wire _w2141_ ;
	wire _w2142_ ;
	wire _w2143_ ;
	wire _w2144_ ;
	wire _w2145_ ;
	wire _w2146_ ;
	wire _w2147_ ;
	wire _w2148_ ;
	wire _w2149_ ;
	wire _w2150_ ;
	wire _w2151_ ;
	wire _w2152_ ;
	wire _w2153_ ;
	wire _w2154_ ;
	wire _w2155_ ;
	wire _w2156_ ;
	wire _w2157_ ;
	wire _w2158_ ;
	wire _w2159_ ;
	wire _w2160_ ;
	wire _w2161_ ;
	wire _w2162_ ;
	wire _w2163_ ;
	wire _w2164_ ;
	wire _w2165_ ;
	wire _w2166_ ;
	wire _w2167_ ;
	wire _w2168_ ;
	wire _w2169_ ;
	wire _w2170_ ;
	wire _w2171_ ;
	wire _w2172_ ;
	wire _w2173_ ;
	wire _w2174_ ;
	wire _w2175_ ;
	wire _w2176_ ;
	wire _w2177_ ;
	wire _w2178_ ;
	wire _w2179_ ;
	wire _w2180_ ;
	wire _w2181_ ;
	wire _w2182_ ;
	wire _w2183_ ;
	wire _w2184_ ;
	wire _w2185_ ;
	wire _w2186_ ;
	wire _w2187_ ;
	wire _w2188_ ;
	wire _w2189_ ;
	wire _w2190_ ;
	wire _w2191_ ;
	wire _w2192_ ;
	wire _w2193_ ;
	wire _w2194_ ;
	wire _w2195_ ;
	wire _w2196_ ;
	wire _w2197_ ;
	wire _w2198_ ;
	wire _w2199_ ;
	wire _w2200_ ;
	wire _w2201_ ;
	wire _w2202_ ;
	wire _w2203_ ;
	wire _w2204_ ;
	wire _w2205_ ;
	wire _w2206_ ;
	wire _w2207_ ;
	wire _w2208_ ;
	wire _w2209_ ;
	wire _w2210_ ;
	wire _w2211_ ;
	wire _w2212_ ;
	wire _w2213_ ;
	wire _w2214_ ;
	wire _w2215_ ;
	wire _w2216_ ;
	wire _w2217_ ;
	wire _w2218_ ;
	wire _w2219_ ;
	wire _w2220_ ;
	wire _w2221_ ;
	wire _w2222_ ;
	wire _w2223_ ;
	wire _w2224_ ;
	wire _w2225_ ;
	wire _w2226_ ;
	wire _w2227_ ;
	wire _w2228_ ;
	wire _w2229_ ;
	wire _w2230_ ;
	wire _w2231_ ;
	wire _w2232_ ;
	wire _w2233_ ;
	wire _w2234_ ;
	wire _w2235_ ;
	wire _w2236_ ;
	wire _w2237_ ;
	wire _w2238_ ;
	wire _w2239_ ;
	wire _w2240_ ;
	wire _w2241_ ;
	wire _w2242_ ;
	wire _w2243_ ;
	wire _w2244_ ;
	wire _w2245_ ;
	wire _w2246_ ;
	wire _w2247_ ;
	wire _w2248_ ;
	wire _w2249_ ;
	wire _w2250_ ;
	wire _w2251_ ;
	wire _w2252_ ;
	wire _w2253_ ;
	wire _w2254_ ;
	wire _w2255_ ;
	wire _w2256_ ;
	wire _w2257_ ;
	wire _w2258_ ;
	wire _w2259_ ;
	wire _w2260_ ;
	wire _w2261_ ;
	wire _w2262_ ;
	wire _w2263_ ;
	wire _w2264_ ;
	wire _w2265_ ;
	wire _w2266_ ;
	wire _w2267_ ;
	wire _w2268_ ;
	wire _w2269_ ;
	wire _w2270_ ;
	wire _w2271_ ;
	wire _w2272_ ;
	wire _w2273_ ;
	wire _w2274_ ;
	wire _w2275_ ;
	wire _w2276_ ;
	wire _w2277_ ;
	wire _w2278_ ;
	wire _w2279_ ;
	wire _w2280_ ;
	wire _w2281_ ;
	wire _w2282_ ;
	wire _w2283_ ;
	wire _w2284_ ;
	wire _w2285_ ;
	wire _w2286_ ;
	wire _w2287_ ;
	wire _w2288_ ;
	wire _w2289_ ;
	wire _w2290_ ;
	wire _w2291_ ;
	wire _w2292_ ;
	wire _w2293_ ;
	wire _w2294_ ;
	wire _w2295_ ;
	wire _w2296_ ;
	wire _w2297_ ;
	wire _w2298_ ;
	wire _w2299_ ;
	wire _w2300_ ;
	wire _w2301_ ;
	wire _w2302_ ;
	wire _w2303_ ;
	wire _w2304_ ;
	wire _w2305_ ;
	wire _w2306_ ;
	wire _w2307_ ;
	wire _w2308_ ;
	wire _w2309_ ;
	wire _w2310_ ;
	wire _w2311_ ;
	wire _w2312_ ;
	wire _w2313_ ;
	wire _w2314_ ;
	wire _w2315_ ;
	wire _w2316_ ;
	wire _w2317_ ;
	wire _w2318_ ;
	wire _w2319_ ;
	wire _w2320_ ;
	wire _w2321_ ;
	wire _w2322_ ;
	wire _w2323_ ;
	wire _w2324_ ;
	wire _w2325_ ;
	wire _w2326_ ;
	wire _w2327_ ;
	wire _w2328_ ;
	wire _w2329_ ;
	wire _w2330_ ;
	wire _w2331_ ;
	wire _w2332_ ;
	wire _w2333_ ;
	wire _w2334_ ;
	wire _w2335_ ;
	wire _w2336_ ;
	wire _w2337_ ;
	wire _w2338_ ;
	wire _w2339_ ;
	wire _w2340_ ;
	wire _w2341_ ;
	wire _w2342_ ;
	wire _w2343_ ;
	wire _w2344_ ;
	wire _w2345_ ;
	wire _w2346_ ;
	wire _w2347_ ;
	wire _w2348_ ;
	wire _w2349_ ;
	wire _w2350_ ;
	wire _w2351_ ;
	wire _w2352_ ;
	wire _w2353_ ;
	wire _w2354_ ;
	wire _w2355_ ;
	wire _w2356_ ;
	wire _w2357_ ;
	wire _w2358_ ;
	wire _w2359_ ;
	wire _w2360_ ;
	wire _w2361_ ;
	wire _w2362_ ;
	wire _w2363_ ;
	wire _w2364_ ;
	wire _w2365_ ;
	wire _w2366_ ;
	wire _w2367_ ;
	wire _w2368_ ;
	wire _w2369_ ;
	wire _w2370_ ;
	wire _w2371_ ;
	wire _w2372_ ;
	wire _w2373_ ;
	wire _w2374_ ;
	wire _w2375_ ;
	wire _w2376_ ;
	wire _w2377_ ;
	wire _w2378_ ;
	wire _w2379_ ;
	wire _w2380_ ;
	wire _w2381_ ;
	wire _w2382_ ;
	wire _w2383_ ;
	wire _w2384_ ;
	wire _w2385_ ;
	wire _w2386_ ;
	wire _w2387_ ;
	wire _w2388_ ;
	wire _w2389_ ;
	wire _w2390_ ;
	wire _w5121_ ;
	wire _w5122_ ;
	wire _w5123_ ;
	wire _w5124_ ;
	wire _w5125_ ;
	wire _w5126_ ;
	wire _w5127_ ;
	wire _w5128_ ;
	wire _w5129_ ;
	wire _w5130_ ;
	wire _w5131_ ;
	wire _w5132_ ;
	wire _w5133_ ;
	wire _w5134_ ;
	wire _w5135_ ;
	wire _w5136_ ;
	wire _w5137_ ;
	wire _w5138_ ;
	wire _w5139_ ;
	wire _w5140_ ;
	wire _w5141_ ;
	wire _w5142_ ;
	wire _w5143_ ;
	wire _w5144_ ;
	wire _w5145_ ;
	wire _w5146_ ;
	wire _w5147_ ;
	wire _w5148_ ;
	wire _w5149_ ;
	wire _w5150_ ;
	wire _w5151_ ;
	wire _w5152_ ;
	wire _w5153_ ;
	wire _w5154_ ;
	wire _w5155_ ;
	wire _w5156_ ;
	wire _w5157_ ;
	wire _w5158_ ;
	wire _w5159_ ;
	wire _w5160_ ;
	wire _w5161_ ;
	wire _w5162_ ;
	wire _w5163_ ;
	wire _w5164_ ;
	wire _w5165_ ;
	wire _w5166_ ;
	wire _w5167_ ;
	wire _w5168_ ;
	wire _w5169_ ;
	wire _w5170_ ;
	wire _w5171_ ;
	wire _w5172_ ;
	wire _w5173_ ;
	wire _w5174_ ;
	wire _w5175_ ;
	wire _w5176_ ;
	wire _w5177_ ;
	wire _w5178_ ;
	wire _w5179_ ;
	wire _w5180_ ;
	wire _w5181_ ;
	wire _w5182_ ;
	wire _w5183_ ;
	wire _w5184_ ;
	wire _w5185_ ;
	wire _w5186_ ;
	wire _w5187_ ;
	wire _w5188_ ;
	wire _w5189_ ;
	wire _w5190_ ;
	wire _w5191_ ;
	wire _w5192_ ;
	wire _w5193_ ;
	wire _w5194_ ;
	wire _w5195_ ;
	wire _w5196_ ;
	wire _w5197_ ;
	wire _w5198_ ;
	wire _w5199_ ;
	wire _w5200_ ;
	wire _w5201_ ;
	wire _w5202_ ;
	wire _w5203_ ;
	wire _w5204_ ;
	wire _w5205_ ;
	wire _w5206_ ;
	wire _w5207_ ;
	wire _w5208_ ;
	wire _w5209_ ;
	wire _w5210_ ;
	wire _w5211_ ;
	wire _w5212_ ;
	wire _w5213_ ;
	wire _w5214_ ;
	wire _w5215_ ;
	wire _w5216_ ;
	wire _w5217_ ;
	wire _w5218_ ;
	wire _w5219_ ;
	wire _w5220_ ;
	wire _w5221_ ;
	wire _w5222_ ;
	wire _w5223_ ;
	wire _w5224_ ;
	wire _w5225_ ;
	wire _w5226_ ;
	wire _w5227_ ;
	wire _w5228_ ;
	wire _w5229_ ;
	wire _w5230_ ;
	wire _w5231_ ;
	wire _w5232_ ;
	wire _w5233_ ;
	wire _w5234_ ;
	wire _w5235_ ;
	wire _w5236_ ;
	wire _w5237_ ;
	wire _w5238_ ;
	wire _w5239_ ;
	wire _w5240_ ;
	wire _w5241_ ;
	wire _w5242_ ;
	wire _w5243_ ;
	wire _w5244_ ;
	wire _w5245_ ;
	wire _w5246_ ;
	wire _w5247_ ;
	wire _w5248_ ;
	wire _w5249_ ;
	wire _w5250_ ;
	wire _w5251_ ;
	wire _w5252_ ;
	wire _w5253_ ;
	wire _w5254_ ;
	wire _w5255_ ;
	wire _w5256_ ;
	wire _w5257_ ;
	wire _w5258_ ;
	wire _w5259_ ;
	wire _w5260_ ;
	wire _w5261_ ;
	wire _w5262_ ;
	wire _w5263_ ;
	wire _w5264_ ;
	wire _w5265_ ;
	wire _w5266_ ;
	wire _w5267_ ;
	wire _w5268_ ;
	wire _w5269_ ;
	wire _w5270_ ;
	wire _w5271_ ;
	wire _w5272_ ;
	wire _w5273_ ;
	wire _w5274_ ;
	wire _w5275_ ;
	wire _w5276_ ;
	wire _w5277_ ;
	wire _w5278_ ;
	wire _w5279_ ;
	wire _w5280_ ;
	wire _w5281_ ;
	wire _w5282_ ;
	wire _w5283_ ;
	wire _w5284_ ;
	wire _w5285_ ;
	wire _w5286_ ;
	wire _w5287_ ;
	wire _w5288_ ;
	wire _w5289_ ;
	wire _w5290_ ;
	wire _w5291_ ;
	wire _w5292_ ;
	wire _w5293_ ;
	wire _w5294_ ;
	wire _w5295_ ;
	wire _w5296_ ;
	wire _w5297_ ;
	wire _w5298_ ;
	wire _w5299_ ;
	wire _w5300_ ;
	wire _w5301_ ;
	wire _w5302_ ;
	wire _w5303_ ;
	wire _w5304_ ;
	wire _w5305_ ;
	wire _w5306_ ;
	wire _w5307_ ;
	wire _w5308_ ;
	wire _w5309_ ;
	wire _w5310_ ;
	wire _w5311_ ;
	wire _w5312_ ;
	wire _w5313_ ;
	wire _w5314_ ;
	wire _w5315_ ;
	wire _w5316_ ;
	wire _w5317_ ;
	wire _w5318_ ;
	wire _w5319_ ;
	wire _w5320_ ;
	wire _w5321_ ;
	wire _w5322_ ;
	wire _w5323_ ;
	wire _w5324_ ;
	wire _w5325_ ;
	wire _w5326_ ;
	wire _w5327_ ;
	wire _w5328_ ;
	wire _w5329_ ;
	wire _w5330_ ;
	wire _w5331_ ;
	wire _w5332_ ;
	wire _w5333_ ;
	wire _w5334_ ;
	wire _w5335_ ;
	wire _w5336_ ;
	wire _w5337_ ;
	wire _w5338_ ;
	wire _w5339_ ;
	wire _w5340_ ;
	wire _w5341_ ;
	wire _w5342_ ;
	wire _w5343_ ;
	wire _w5344_ ;
	wire _w5345_ ;
	wire _w5346_ ;
	wire _w5347_ ;
	wire _w5348_ ;
	wire _w5349_ ;
	wire _w5350_ ;
	wire _w5351_ ;
	wire _w5352_ ;
	wire _w5353_ ;
	wire _w5354_ ;
	wire _w5355_ ;
	wire _w5356_ ;
	wire _w5357_ ;
	wire _w5358_ ;
	wire _w5359_ ;
	wire _w5360_ ;
	wire _w5361_ ;
	wire _w5362_ ;
	wire _w5363_ ;
	wire _w5364_ ;
	wire _w5365_ ;
	wire _w5366_ ;
	wire _w5367_ ;
	wire _w5368_ ;
	wire _w5369_ ;
	wire _w5370_ ;
	wire _w5371_ ;
	wire _w5372_ ;
	wire _w5373_ ;
	wire _w5374_ ;
	wire _w5375_ ;
	wire _w5376_ ;
	wire _w5377_ ;
	wire _w5378_ ;
	wire _w5379_ ;
	wire _w5380_ ;
	wire _w5381_ ;
	wire _w5382_ ;
	wire _w5383_ ;
	wire _w5384_ ;
	wire _w5385_ ;
	wire _w5386_ ;
	wire _w5387_ ;
	wire _w5388_ ;
	wire _w5389_ ;
	wire _w5390_ ;
	wire _w5391_ ;
	wire _w5392_ ;
	wire _w5393_ ;
	wire _w5394_ ;
	wire _w5395_ ;
	wire _w5396_ ;
	wire _w5397_ ;
	wire _w5398_ ;
	wire _w5399_ ;
	wire _w5400_ ;
	wire _w5401_ ;
	wire _w5402_ ;
	wire _w5403_ ;
	wire _w5404_ ;
	wire _w5405_ ;
	wire _w5406_ ;
	wire _w5407_ ;
	wire _w5408_ ;
	wire _w5409_ ;
	wire _w5410_ ;
	wire _w5411_ ;
	wire _w5412_ ;
	wire _w5413_ ;
	wire _w5414_ ;
	wire _w5415_ ;
	wire _w5416_ ;
	wire _w5417_ ;
	wire _w5418_ ;
	wire _w5419_ ;
	wire _w5420_ ;
	wire _w5421_ ;
	wire _w5422_ ;
	wire _w5423_ ;
	wire _w5424_ ;
	wire _w5425_ ;
	wire _w5426_ ;
	wire _w5427_ ;
	wire _w5428_ ;
	wire _w5429_ ;
	wire _w5430_ ;
	wire _w5431_ ;
	wire _w5432_ ;
	wire _w5433_ ;
	wire _w5434_ ;
	wire _w5435_ ;
	wire _w5436_ ;
	wire _w5437_ ;
	wire _w5438_ ;
	wire _w5439_ ;
	wire _w5440_ ;
	wire _w5441_ ;
	wire _w5442_ ;
	wire _w5443_ ;
	wire _w5444_ ;
	wire _w5445_ ;
	wire _w5446_ ;
	wire _w5447_ ;
	wire _w5448_ ;
	wire _w5449_ ;
	wire _w5450_ ;
	wire _w5451_ ;
	wire _w5452_ ;
	wire _w5453_ ;
	wire _w5454_ ;
	wire _w5455_ ;
	wire _w5456_ ;
	wire _w5457_ ;
	wire _w5458_ ;
	wire _w5459_ ;
	wire _w5460_ ;
	wire _w5461_ ;
	wire _w5462_ ;
	wire _w5463_ ;
	wire _w5464_ ;
	wire _w5465_ ;
	wire _w5466_ ;
	wire _w5467_ ;
	wire _w5468_ ;
	wire _w5469_ ;
	wire _w5470_ ;
	wire _w5471_ ;
	wire _w5472_ ;
	wire _w5473_ ;
	wire _w5474_ ;
	wire _w5475_ ;
	wire _w5476_ ;
	wire _w5477_ ;
	wire _w5478_ ;
	wire _w5479_ ;
	wire _w5480_ ;
	wire _w5481_ ;
	wire _w5482_ ;
	wire _w5483_ ;
	wire _w5484_ ;
	wire _w5485_ ;
	wire _w5486_ ;
	wire _w5487_ ;
	wire _w5488_ ;
	wire _w5489_ ;
	wire _w5490_ ;
	wire _w5491_ ;
	wire _w5492_ ;
	wire _w5493_ ;
	wire _w5494_ ;
	wire _w5495_ ;
	wire _w5496_ ;
	wire _w5497_ ;
	wire _w5498_ ;
	wire _w5499_ ;
	wire _w5500_ ;
	wire _w5501_ ;
	wire _w5502_ ;
	wire _w5503_ ;
	wire _w5504_ ;
	wire _w5505_ ;
	wire _w5506_ ;
	wire _w5507_ ;
	wire _w5508_ ;
	wire _w5509_ ;
	wire _w5510_ ;
	wire _w5511_ ;
	wire _w5512_ ;
	wire _w5513_ ;
	wire _w5514_ ;
	wire _w5515_ ;
	wire _w5516_ ;
	wire _w5517_ ;
	wire _w5518_ ;
	wire _w5519_ ;
	wire _w5520_ ;
	wire _w5521_ ;
	wire _w5522_ ;
	wire _w5523_ ;
	wire _w5524_ ;
	wire _w5525_ ;
	wire _w5526_ ;
	wire _w5527_ ;
	wire _w5528_ ;
	wire _w5529_ ;
	wire _w5530_ ;
	wire _w5531_ ;
	wire _w5532_ ;
	wire _w5533_ ;
	wire _w5534_ ;
	wire _w5535_ ;
	wire _w5536_ ;
	wire _w5537_ ;
	wire _w5538_ ;
	wire _w5539_ ;
	wire _w5540_ ;
	wire _w5541_ ;
	wire _w5542_ ;
	wire _w5543_ ;
	wire _w5544_ ;
	wire _w5545_ ;
	wire _w5546_ ;
	wire _w5547_ ;
	wire _w5548_ ;
	wire _w5549_ ;
	wire _w5550_ ;
	wire _w5551_ ;
	wire _w5552_ ;
	wire _w5553_ ;
	wire _w5554_ ;
	wire _w5555_ ;
	wire _w5556_ ;
	wire _w5557_ ;
	wire _w5558_ ;
	wire _w5559_ ;
	wire _w5560_ ;
	wire _w5561_ ;
	wire _w5562_ ;
	wire _w5563_ ;
	wire _w5564_ ;
	wire _w5565_ ;
	wire _w5566_ ;
	wire _w5567_ ;
	wire _w5568_ ;
	wire _w5569_ ;
	wire _w5570_ ;
	wire _w5571_ ;
	wire _w5572_ ;
	wire _w5573_ ;
	wire _w5574_ ;
	wire _w5575_ ;
	wire _w5576_ ;
	wire _w5577_ ;
	wire _w5578_ ;
	wire _w5579_ ;
	wire _w5580_ ;
	wire _w5581_ ;
	wire _w5582_ ;
	wire _w5583_ ;
	wire _w5584_ ;
	wire _w5585_ ;
	wire _w5586_ ;
	wire _w5587_ ;
	wire _w5588_ ;
	wire _w5589_ ;
	wire _w5590_ ;
	wire _w5591_ ;
	wire _w5592_ ;
	wire _w5593_ ;
	wire _w5594_ ;
	wire _w5595_ ;
	wire _w5596_ ;
	wire _w5597_ ;
	wire _w5598_ ;
	wire _w5599_ ;
	wire _w5600_ ;
	wire _w5601_ ;
	wire _w5602_ ;
	wire _w5603_ ;
	wire _w5604_ ;
	wire _w5605_ ;
	wire _w5606_ ;
	wire _w5607_ ;
	wire _w5608_ ;
	wire _w5609_ ;
	wire _w5610_ ;
	wire _w5611_ ;
	wire _w5612_ ;
	wire _w5613_ ;
	wire _w5614_ ;
	wire _w5615_ ;
	wire _w5616_ ;
	wire _w5617_ ;
	wire _w5618_ ;
	wire _w5619_ ;
	wire _w5620_ ;
	wire _w5621_ ;
	wire _w5622_ ;
	wire _w5623_ ;
	wire _w5624_ ;
	wire _w5625_ ;
	wire _w5626_ ;
	wire _w5627_ ;
	wire _w5628_ ;
	wire _w5629_ ;
	wire _w5630_ ;
	wire _w5631_ ;
	wire _w5632_ ;
	wire _w5633_ ;
	wire _w5634_ ;
	wire _w5635_ ;
	wire _w5636_ ;
	wire _w5637_ ;
	wire _w5638_ ;
	wire _w5639_ ;
	wire _w5640_ ;
	wire _w5641_ ;
	wire _w5642_ ;
	wire _w5643_ ;
	wire _w5644_ ;
	wire _w5645_ ;
	wire _w5646_ ;
	wire _w5647_ ;
	wire _w5648_ ;
	wire _w5649_ ;
	wire _w5650_ ;
	wire _w5651_ ;
	wire _w5652_ ;
	wire _w5653_ ;
	wire _w5654_ ;
	wire _w5655_ ;
	wire _w5656_ ;
	wire _w5657_ ;
	wire _w5658_ ;
	wire _w5659_ ;
	wire _w5660_ ;
	wire _w5661_ ;
	wire _w5662_ ;
	wire _w5663_ ;
	wire _w5664_ ;
	wire _w5665_ ;
	wire _w5666_ ;
	wire _w5667_ ;
	wire _w5668_ ;
	wire _w5669_ ;
	wire _w5670_ ;
	wire _w5671_ ;
	wire _w5672_ ;
	wire _w5673_ ;
	wire _w5674_ ;
	wire _w5675_ ;
	wire _w5676_ ;
	wire _w5677_ ;
	wire _w5678_ ;
	wire _w5679_ ;
	wire _w5680_ ;
	wire _w5681_ ;
	wire _w5682_ ;
	wire _w5683_ ;
	wire _w5684_ ;
	wire _w5685_ ;
	wire _w5686_ ;
	wire _w5687_ ;
	wire _w5688_ ;
	wire _w5689_ ;
	wire _w5690_ ;
	wire _w5691_ ;
	wire _w5692_ ;
	wire _w5693_ ;
	wire _w5694_ ;
	wire _w5695_ ;
	wire _w5696_ ;
	wire _w5697_ ;
	wire _w5698_ ;
	wire _w5699_ ;
	wire _w5700_ ;
	wire _w5701_ ;
	wire _w5702_ ;
	wire _w5703_ ;
	wire _w5704_ ;
	wire _w5705_ ;
	wire _w5706_ ;
	wire _w5707_ ;
	wire _w5708_ ;
	wire _w5709_ ;
	wire _w5710_ ;
	wire _w5711_ ;
	wire _w5712_ ;
	wire _w5713_ ;
	wire _w5714_ ;
	wire _w5715_ ;
	wire _w5716_ ;
	wire _w5717_ ;
	wire _w5718_ ;
	wire _w5719_ ;
	wire _w5720_ ;
	wire _w5721_ ;
	wire _w5722_ ;
	wire _w5723_ ;
	wire _w5724_ ;
	wire _w5725_ ;
	wire _w5726_ ;
	wire _w5727_ ;
	wire _w5728_ ;
	wire _w5729_ ;
	wire _w5730_ ;
	wire _w5731_ ;
	wire _w5732_ ;
	wire _w5733_ ;
	wire _w5734_ ;
	wire _w5735_ ;
	wire _w5736_ ;
	wire _w5737_ ;
	wire _w5738_ ;
	wire _w5739_ ;
	wire _w5740_ ;
	wire _w5741_ ;
	wire _w5742_ ;
	wire _w5743_ ;
	wire _w5744_ ;
	wire _w5745_ ;
	wire _w5746_ ;
	wire _w5747_ ;
	wire _w5748_ ;
	wire _w5749_ ;
	wire _w5750_ ;
	wire _w5751_ ;
	wire _w5752_ ;
	wire _w5753_ ;
	wire _w5754_ ;
	wire _w5755_ ;
	wire _w5756_ ;
	wire _w5757_ ;
	wire _w5758_ ;
	wire _w5759_ ;
	wire _w5760_ ;
	wire _w5761_ ;
	wire _w5762_ ;
	wire _w5763_ ;
	wire _w5764_ ;
	wire _w5765_ ;
	wire _w5766_ ;
	wire _w5767_ ;
	wire _w5768_ ;
	wire _w5769_ ;
	wire _w5770_ ;
	wire _w5771_ ;
	wire _w5772_ ;
	wire _w5773_ ;
	wire _w5774_ ;
	wire _w5775_ ;
	wire _w5776_ ;
	wire _w5777_ ;
	wire _w5778_ ;
	wire _w5779_ ;
	wire _w5780_ ;
	wire _w5781_ ;
	wire _w5782_ ;
	wire _w5783_ ;
	wire _w5784_ ;
	wire _w5785_ ;
	wire _w5786_ ;
	wire _w5787_ ;
	wire _w5788_ ;
	wire _w5789_ ;
	wire _w5790_ ;
	wire _w5791_ ;
	wire _w5792_ ;
	wire _w5793_ ;
	wire _w5794_ ;
	wire _w5795_ ;
	wire _w5796_ ;
	wire _w5797_ ;
	wire _w5798_ ;
	wire _w5799_ ;
	wire _w5800_ ;
	wire _w5801_ ;
	wire _w5802_ ;
	wire _w5803_ ;
	wire _w5804_ ;
	wire _w5805_ ;
	wire _w5806_ ;
	wire _w5807_ ;
	wire _w5808_ ;
	wire _w5809_ ;
	wire _w5810_ ;
	wire _w5811_ ;
	wire _w5812_ ;
	wire _w5813_ ;
	wire _w5814_ ;
	wire _w5815_ ;
	wire _w5816_ ;
	wire _w5817_ ;
	wire _w5818_ ;
	wire _w5819_ ;
	wire _w5820_ ;
	wire _w5821_ ;
	wire _w5822_ ;
	wire _w5823_ ;
	wire _w5824_ ;
	wire _w5825_ ;
	wire _w5826_ ;
	wire _w5827_ ;
	wire _w5828_ ;
	wire _w5829_ ;
	wire _w5830_ ;
	wire _w5831_ ;
	wire _w5832_ ;
	wire _w5833_ ;
	wire _w5834_ ;
	wire _w5835_ ;
	wire _w5836_ ;
	wire _w5837_ ;
	wire _w5838_ ;
	wire _w5839_ ;
	wire _w5840_ ;
	wire _w5841_ ;
	wire _w5842_ ;
	wire _w5843_ ;
	wire _w5844_ ;
	wire _w5845_ ;
	wire _w5846_ ;
	wire _w5847_ ;
	wire _w5848_ ;
	wire _w5849_ ;
	wire _w5850_ ;
	wire _w5851_ ;
	wire _w5852_ ;
	wire _w5853_ ;
	wire _w5854_ ;
	wire _w5855_ ;
	wire _w5856_ ;
	wire _w5857_ ;
	wire _w5858_ ;
	wire _w5859_ ;
	wire _w5860_ ;
	wire _w5861_ ;
	wire _w5862_ ;
	wire _w5863_ ;
	wire _w5864_ ;
	wire _w5865_ ;
	wire _w5866_ ;
	wire _w5867_ ;
	wire _w5868_ ;
	wire _w5869_ ;
	wire _w5870_ ;
	wire _w5871_ ;
	wire _w5872_ ;
	wire _w5873_ ;
	wire _w5874_ ;
	wire _w5875_ ;
	wire _w5876_ ;
	wire _w5877_ ;
	wire _w5878_ ;
	wire _w5879_ ;
	wire _w5880_ ;
	wire _w5881_ ;
	wire _w5882_ ;
	wire _w5883_ ;
	wire _w5884_ ;
	wire _w5885_ ;
	wire _w5886_ ;
	wire _w5887_ ;
	wire _w5888_ ;
	wire _w5889_ ;
	wire _w5890_ ;
	wire _w5891_ ;
	wire _w5892_ ;
	wire _w5893_ ;
	wire _w5894_ ;
	wire _w5895_ ;
	wire _w5896_ ;
	wire _w5897_ ;
	wire _w5898_ ;
	wire _w5899_ ;
	wire _w5900_ ;
	wire _w5901_ ;
	wire _w5902_ ;
	wire _w5903_ ;
	wire _w5904_ ;
	wire _w5905_ ;
	wire _w5906_ ;
	wire _w5907_ ;
	wire _w5908_ ;
	wire _w5909_ ;
	wire _w5910_ ;
	wire _w5911_ ;
	wire _w5912_ ;
	wire _w5913_ ;
	wire _w5914_ ;
	wire _w5915_ ;
	wire _w5916_ ;
	wire _w5917_ ;
	wire _w5918_ ;
	wire _w5919_ ;
	wire _w5920_ ;
	wire _w5921_ ;
	wire _w5922_ ;
	wire _w5923_ ;
	wire _w5924_ ;
	wire _w5925_ ;
	wire _w5926_ ;
	wire _w5927_ ;
	wire _w5928_ ;
	wire _w5929_ ;
	wire _w5930_ ;
	wire _w5931_ ;
	wire _w5932_ ;
	wire _w5933_ ;
	wire _w5934_ ;
	wire _w5935_ ;
	wire _w5936_ ;
	wire _w5937_ ;
	wire _w5938_ ;
	wire _w5939_ ;
	wire _w5940_ ;
	wire _w5941_ ;
	wire _w5942_ ;
	wire _w5943_ ;
	wire _w5944_ ;
	wire _w5945_ ;
	wire _w5946_ ;
	wire _w5947_ ;
	wire _w5948_ ;
	wire _w5949_ ;
	wire _w5950_ ;
	wire _w5951_ ;
	wire _w5952_ ;
	wire _w5953_ ;
	wire _w5954_ ;
	wire _w5955_ ;
	wire _w5956_ ;
	wire _w5957_ ;
	wire _w5958_ ;
	wire _w5959_ ;
	wire _w5960_ ;
	wire _w5961_ ;
	wire _w5962_ ;
	wire _w5963_ ;
	wire _w5964_ ;
	wire _w5965_ ;
	wire _w5966_ ;
	wire _w5967_ ;
	wire _w5968_ ;
	wire _w5969_ ;
	wire _w5970_ ;
	wire _w5971_ ;
	wire _w5972_ ;
	wire _w5973_ ;
	wire _w5974_ ;
	wire _w5975_ ;
	wire _w5976_ ;
	wire _w5977_ ;
	wire _w5978_ ;
	wire _w5979_ ;
	wire _w5980_ ;
	wire _w5981_ ;
	wire _w5982_ ;
	wire _w5983_ ;
	wire _w5984_ ;
	wire _w5985_ ;
	wire _w5986_ ;
	wire _w5987_ ;
	wire _w5988_ ;
	wire _w5989_ ;
	wire _w5990_ ;
	wire _w5991_ ;
	wire _w5992_ ;
	wire _w5993_ ;
	wire _w5994_ ;
	wire _w5995_ ;
	wire _w5996_ ;
	wire _w5997_ ;
	wire _w5998_ ;
	wire _w5999_ ;
	wire _w6000_ ;
	wire _w6001_ ;
	wire _w6002_ ;
	wire _w6003_ ;
	wire _w6004_ ;
	wire _w6005_ ;
	wire _w6006_ ;
	wire _w6007_ ;
	wire _w6008_ ;
	wire _w6009_ ;
	wire _w6010_ ;
	wire _w6011_ ;
	wire _w6012_ ;
	wire _w6013_ ;
	wire _w6014_ ;
	wire _w6015_ ;
	wire _w6016_ ;
	wire _w6017_ ;
	wire _w6018_ ;
	wire _w6019_ ;
	wire _w6020_ ;
	wire _w6021_ ;
	wire _w6022_ ;
	wire _w6023_ ;
	wire _w6024_ ;
	wire _w6025_ ;
	wire _w6026_ ;
	wire _w6027_ ;
	wire _w6028_ ;
	wire _w6029_ ;
	wire _w6030_ ;
	wire _w6031_ ;
	wire _w6032_ ;
	wire _w6033_ ;
	wire _w6034_ ;
	wire _w6035_ ;
	wire _w6036_ ;
	wire _w6037_ ;
	wire _w6038_ ;
	wire _w6039_ ;
	wire _w6040_ ;
	wire _w6041_ ;
	wire _w6042_ ;
	wire _w6043_ ;
	wire _w6044_ ;
	wire _w6045_ ;
	wire _w6046_ ;
	wire _w6047_ ;
	wire _w6048_ ;
	wire _w6049_ ;
	wire _w6050_ ;
	wire _w6051_ ;
	wire _w6052_ ;
	wire _w6053_ ;
	wire _w6054_ ;
	wire _w6055_ ;
	wire _w6056_ ;
	wire _w6057_ ;
	wire _w6058_ ;
	wire _w6059_ ;
	wire _w6060_ ;
	wire _w6061_ ;
	wire _w6062_ ;
	wire _w6063_ ;
	wire _w6064_ ;
	wire _w6065_ ;
	wire _w6066_ ;
	wire _w6067_ ;
	wire _w6068_ ;
	wire _w6069_ ;
	wire _w6070_ ;
	wire _w6071_ ;
	wire _w6072_ ;
	wire _w6073_ ;
	wire _w6074_ ;
	wire _w6075_ ;
	wire _w6076_ ;
	wire _w6077_ ;
	wire _w6078_ ;
	wire _w6079_ ;
	wire _w6080_ ;
	wire _w6081_ ;
	wire _w6082_ ;
	wire _w6083_ ;
	wire _w6084_ ;
	wire _w6085_ ;
	wire _w6086_ ;
	wire _w6087_ ;
	wire _w6088_ ;
	wire _w6089_ ;
	wire _w6090_ ;
	wire _w6091_ ;
	wire _w6092_ ;
	wire _w6093_ ;
	wire _w6094_ ;
	wire _w6095_ ;
	wire _w6096_ ;
	wire _w6097_ ;
	wire _w6098_ ;
	wire _w6099_ ;
	wire _w6100_ ;
	wire _w6101_ ;
	wire _w6102_ ;
	wire _w6103_ ;
	wire _w6104_ ;
	wire _w6105_ ;
	wire _w6106_ ;
	wire _w6107_ ;
	wire _w6108_ ;
	wire _w6109_ ;
	wire _w6110_ ;
	wire _w6111_ ;
	wire _w6112_ ;
	wire _w6113_ ;
	wire _w6114_ ;
	wire _w6115_ ;
	wire _w6116_ ;
	wire _w6117_ ;
	wire _w6118_ ;
	wire _w6119_ ;
	wire _w6120_ ;
	wire _w6121_ ;
	wire _w6122_ ;
	wire _w6123_ ;
	wire _w6124_ ;
	wire _w6125_ ;
	wire _w6126_ ;
	wire _w6127_ ;
	wire _w6128_ ;
	wire _w6129_ ;
	wire _w6130_ ;
	wire _w6131_ ;
	wire _w6132_ ;
	wire _w6133_ ;
	wire _w6134_ ;
	wire _w6135_ ;
	wire _w6136_ ;
	wire _w6137_ ;
	wire _w6138_ ;
	wire _w6139_ ;
	wire _w6140_ ;
	wire _w6141_ ;
	wire _w6142_ ;
	wire _w6143_ ;
	wire _w6144_ ;
	wire _w6145_ ;
	wire _w6146_ ;
	wire _w6147_ ;
	wire _w6148_ ;
	wire _w6149_ ;
	wire _w6150_ ;
	wire _w6151_ ;
	wire _w6152_ ;
	wire _w6153_ ;
	wire _w6154_ ;
	wire _w6155_ ;
	wire _w6156_ ;
	wire _w6157_ ;
	wire _w6158_ ;
	wire _w6159_ ;
	wire _w6160_ ;
	wire _w6161_ ;
	wire _w6162_ ;
	wire _w6163_ ;
	wire _w6164_ ;
	wire _w6165_ ;
	wire _w6166_ ;
	wire _w6167_ ;
	wire _w6168_ ;
	wire _w6169_ ;
	wire _w6170_ ;
	wire _w6171_ ;
	wire _w6172_ ;
	wire _w6173_ ;
	wire _w6174_ ;
	wire _w6175_ ;
	wire _w6176_ ;
	wire _w6177_ ;
	wire _w6178_ ;
	wire _w6179_ ;
	wire _w6180_ ;
	wire _w6181_ ;
	wire _w6182_ ;
	wire _w6183_ ;
	wire _w6184_ ;
	wire _w6185_ ;
	wire _w6186_ ;
	wire _w6187_ ;
	wire _w6188_ ;
	wire _w6189_ ;
	wire _w6190_ ;
	wire _w6191_ ;
	wire _w6192_ ;
	wire _w6193_ ;
	wire _w6194_ ;
	wire _w6195_ ;
	wire _w6196_ ;
	wire _w6197_ ;
	wire _w6198_ ;
	wire _w6199_ ;
	wire _w6200_ ;
	wire _w6201_ ;
	wire _w6202_ ;
	wire _w6203_ ;
	wire _w6204_ ;
	wire _w6205_ ;
	wire _w6206_ ;
	wire _w6207_ ;
	wire _w6208_ ;
	wire _w6209_ ;
	wire _w6210_ ;
	wire _w6211_ ;
	wire _w6212_ ;
	wire _w6213_ ;
	wire _w6214_ ;
	wire _w6215_ ;
	wire _w6216_ ;
	wire _w6217_ ;
	wire _w6218_ ;
	wire _w6219_ ;
	wire _w6220_ ;
	wire _w6221_ ;
	wire _w6222_ ;
	wire _w6223_ ;
	wire _w6224_ ;
	wire _w6225_ ;
	wire _w6226_ ;
	wire _w6227_ ;
	wire _w6228_ ;
	wire _w6229_ ;
	wire _w6230_ ;
	wire _w6231_ ;
	wire _w6232_ ;
	wire _w6233_ ;
	wire _w6234_ ;
	wire _w6235_ ;
	wire _w6236_ ;
	wire _w6237_ ;
	wire _w6238_ ;
	wire _w6239_ ;
	wire _w6240_ ;
	wire _w6241_ ;
	wire _w6242_ ;
	wire _w6243_ ;
	wire _w6244_ ;
	wire _w6245_ ;
	wire _w6246_ ;
	wire _w6247_ ;
	wire _w6248_ ;
	wire _w6249_ ;
	wire _w6250_ ;
	wire _w6251_ ;
	wire _w6252_ ;
	wire _w6253_ ;
	wire _w6254_ ;
	wire _w6255_ ;
	wire _w6256_ ;
	wire _w6257_ ;
	wire _w6258_ ;
	wire _w6259_ ;
	wire _w6260_ ;
	wire _w6261_ ;
	wire _w6262_ ;
	wire _w6263_ ;
	wire _w6264_ ;
	wire _w6265_ ;
	wire _w6266_ ;
	wire _w6267_ ;
	wire _w6268_ ;
	wire _w6269_ ;
	wire _w6270_ ;
	wire _w6271_ ;
	wire _w6272_ ;
	wire _w6273_ ;
	wire _w6274_ ;
	wire _w6275_ ;
	wire _w6276_ ;
	wire _w6277_ ;
	wire _w6278_ ;
	wire _w6279_ ;
	wire _w6280_ ;
	wire _w6281_ ;
	wire _w6282_ ;
	wire _w6283_ ;
	wire _w6284_ ;
	wire _w6285_ ;
	wire _w6286_ ;
	wire _w6287_ ;
	wire _w6288_ ;
	wire _w6289_ ;
	wire _w6290_ ;
	wire _w6291_ ;
	wire _w6292_ ;
	wire _w6293_ ;
	wire _w6294_ ;
	wire _w6295_ ;
	wire _w6296_ ;
	wire _w6297_ ;
	wire _w6298_ ;
	wire _w6299_ ;
	wire _w6300_ ;
	wire _w6301_ ;
	wire _w6302_ ;
	wire _w6303_ ;
	wire _w6304_ ;
	wire _w6305_ ;
	wire _w6306_ ;
	wire _w6307_ ;
	wire _w6308_ ;
	wire _w6309_ ;
	wire _w6310_ ;
	wire _w6311_ ;
	wire _w6312_ ;
	wire _w6313_ ;
	wire _w6314_ ;
	wire _w6315_ ;
	wire _w6316_ ;
	wire _w6317_ ;
	wire _w6318_ ;
	wire _w6319_ ;
	wire _w6320_ ;
	wire _w6321_ ;
	wire _w6322_ ;
	wire _w6323_ ;
	wire _w6324_ ;
	wire _w6325_ ;
	wire _w6326_ ;
	wire _w6327_ ;
	wire _w6328_ ;
	wire _w6329_ ;
	wire _w6330_ ;
	wire _w6331_ ;
	wire _w6332_ ;
	wire _w6333_ ;
	wire _w6334_ ;
	wire _w6335_ ;
	wire _w6336_ ;
	wire _w6337_ ;
	wire _w6338_ ;
	wire _w6339_ ;
	wire _w6340_ ;
	wire _w6341_ ;
	wire _w6342_ ;
	wire _w6343_ ;
	wire _w6344_ ;
	wire _w6345_ ;
	wire _w6346_ ;
	wire _w6347_ ;
	wire _w6348_ ;
	wire _w6349_ ;
	wire _w6350_ ;
	wire _w6351_ ;
	wire _w6352_ ;
	wire _w6353_ ;
	wire _w6354_ ;
	wire _w6355_ ;
	wire _w6356_ ;
	wire _w6357_ ;
	wire _w6358_ ;
	wire _w6359_ ;
	wire _w6360_ ;
	wire _w6361_ ;
	wire _w6362_ ;
	wire _w6363_ ;
	wire _w6364_ ;
	wire _w6365_ ;
	wire _w6366_ ;
	wire _w6367_ ;
	wire _w6368_ ;
	wire _w6369_ ;
	wire _w6370_ ;
	wire _w6371_ ;
	wire _w6372_ ;
	wire _w6373_ ;
	wire _w6374_ ;
	wire _w6375_ ;
	wire _w6376_ ;
	wire _w6377_ ;
	wire _w6378_ ;
	wire _w6379_ ;
	wire _w6380_ ;
	wire _w6381_ ;
	wire _w6382_ ;
	wire _w6383_ ;
	wire _w6384_ ;
	wire _w6385_ ;
	wire _w6386_ ;
	wire _w6387_ ;
	wire _w6388_ ;
	wire _w6389_ ;
	wire _w6390_ ;
	wire _w6391_ ;
	wire _w6392_ ;
	wire _w6393_ ;
	wire _w6394_ ;
	wire _w6395_ ;
	wire _w6396_ ;
	wire _w6397_ ;
	wire _w6398_ ;
	wire _w6399_ ;
	wire _w6400_ ;
	wire _w6401_ ;
	wire _w6402_ ;
	wire _w6403_ ;
	wire _w6404_ ;
	wire _w6405_ ;
	wire _w6406_ ;
	wire _w6407_ ;
	wire _w6408_ ;
	wire _w6409_ ;
	wire _w6410_ ;
	wire _w6411_ ;
	wire _w6412_ ;
	wire _w6413_ ;
	wire _w6414_ ;
	wire _w6415_ ;
	wire _w6416_ ;
	wire _w6417_ ;
	wire _w6418_ ;
	wire _w6419_ ;
	wire _w6420_ ;
	wire _w6421_ ;
	wire _w6422_ ;
	wire _w6423_ ;
	wire _w6424_ ;
	wire _w6425_ ;
	wire _w6426_ ;
	wire _w6427_ ;
	wire _w6428_ ;
	wire _w6429_ ;
	wire _w6430_ ;
	wire _w6431_ ;
	wire _w6432_ ;
	wire _w6433_ ;
	wire _w6434_ ;
	wire _w6435_ ;
	wire _w6436_ ;
	wire _w6437_ ;
	wire _w6438_ ;
	wire _w6439_ ;
	wire _w6440_ ;
	wire _w6441_ ;
	wire _w6442_ ;
	wire _w6443_ ;
	wire _w6444_ ;
	wire _w6445_ ;
	wire _w6446_ ;
	wire _w6447_ ;
	wire _w6448_ ;
	wire _w6449_ ;
	wire _w6450_ ;
	wire _w6451_ ;
	wire _w6452_ ;
	wire _w6453_ ;
	wire _w6454_ ;
	wire _w6455_ ;
	wire _w6456_ ;
	wire _w6457_ ;
	wire _w6458_ ;
	wire _w6459_ ;
	wire _w6460_ ;
	wire _w6461_ ;
	wire _w6462_ ;
	wire _w6463_ ;
	wire _w6464_ ;
	wire _w6465_ ;
	wire _w6466_ ;
	wire _w6467_ ;
	wire _w6468_ ;
	wire _w6469_ ;
	wire _w6470_ ;
	wire _w6471_ ;
	wire _w6472_ ;
	wire _w6473_ ;
	wire _w6474_ ;
	wire _w6475_ ;
	wire _w6476_ ;
	wire _w6477_ ;
	wire _w6478_ ;
	wire _w6479_ ;
	wire _w6480_ ;
	wire _w6481_ ;
	wire _w6482_ ;
	wire _w6483_ ;
	wire _w6484_ ;
	wire _w6485_ ;
	wire _w6486_ ;
	wire _w6487_ ;
	wire _w6488_ ;
	wire _w6489_ ;
	wire _w6490_ ;
	wire _w6491_ ;
	wire _w6492_ ;
	wire _w6493_ ;
	wire _w6494_ ;
	wire _w6495_ ;
	wire _w6496_ ;
	wire _w6497_ ;
	wire _w6498_ ;
	wire _w6499_ ;
	wire _w6500_ ;
	wire _w6501_ ;
	wire _w6502_ ;
	wire _w6503_ ;
	wire _w6504_ ;
	wire _w6505_ ;
	wire _w6506_ ;
	wire _w6507_ ;
	wire _w6508_ ;
	wire _w6509_ ;
	wire _w6510_ ;
	wire _w6511_ ;
	wire _w6512_ ;
	wire _w6513_ ;
	wire _w6514_ ;
	wire _w6515_ ;
	wire _w6516_ ;
	wire _w6517_ ;
	wire _w6518_ ;
	wire _w6519_ ;
	wire _w6520_ ;
	wire _w6521_ ;
	wire _w6522_ ;
	wire _w6523_ ;
	wire _w6524_ ;
	wire _w6525_ ;
	wire _w6526_ ;
	wire _w6527_ ;
	wire _w6528_ ;
	wire _w6529_ ;
	wire _w6530_ ;
	wire _w6531_ ;
	wire _w6532_ ;
	wire _w6533_ ;
	wire _w6534_ ;
	wire _w6535_ ;
	wire _w6536_ ;
	wire _w6537_ ;
	wire _w6538_ ;
	wire _w6539_ ;
	wire _w6540_ ;
	wire _w6541_ ;
	wire _w6542_ ;
	wire _w6543_ ;
	wire _w6544_ ;
	wire _w6545_ ;
	wire _w6546_ ;
	wire _w6547_ ;
	wire _w6548_ ;
	wire _w6549_ ;
	wire _w6550_ ;
	wire _w6551_ ;
	wire _w6552_ ;
	wire _w6553_ ;
	wire _w6554_ ;
	wire _w6555_ ;
	wire _w6556_ ;
	wire _w6557_ ;
	wire _w6558_ ;
	wire _w6559_ ;
	wire _w6560_ ;
	wire _w6561_ ;
	wire _w6562_ ;
	wire _w6563_ ;
	wire _w6564_ ;
	wire _w6565_ ;
	wire _w6566_ ;
	wire _w6567_ ;
	wire _w6568_ ;
	wire _w6569_ ;
	wire _w6570_ ;
	wire _w6571_ ;
	wire _w6572_ ;
	wire _w6573_ ;
	wire _w6574_ ;
	wire _w6575_ ;
	wire _w6576_ ;
	wire _w6577_ ;
	wire _w6578_ ;
	wire _w6579_ ;
	wire _w6580_ ;
	wire _w6581_ ;
	wire _w6582_ ;
	wire _w6583_ ;
	wire _w6584_ ;
	wire _w6585_ ;
	wire _w6586_ ;
	wire _w6587_ ;
	wire _w6588_ ;
	wire _w6589_ ;
	wire _w6590_ ;
	wire _w6591_ ;
	wire _w6592_ ;
	wire _w6593_ ;
	wire _w6594_ ;
	wire _w6595_ ;
	wire _w6596_ ;
	wire _w6597_ ;
	wire _w6598_ ;
	wire _w6599_ ;
	wire _w6600_ ;
	wire _w6601_ ;
	wire _w6602_ ;
	wire _w6603_ ;
	wire _w6604_ ;
	wire _w6605_ ;
	wire _w6606_ ;
	wire _w6607_ ;
	wire _w6608_ ;
	wire _w6609_ ;
	wire _w6610_ ;
	wire _w6611_ ;
	wire _w6612_ ;
	wire _w6613_ ;
	wire _w6614_ ;
	wire _w6615_ ;
	wire _w6616_ ;
	wire _w6617_ ;
	wire _w6618_ ;
	wire _w6619_ ;
	wire _w6620_ ;
	wire _w6621_ ;
	wire _w6622_ ;
	wire _w6623_ ;
	wire _w6624_ ;
	wire _w6625_ ;
	wire _w6626_ ;
	wire _w6627_ ;
	wire _w6628_ ;
	wire _w6629_ ;
	wire _w6630_ ;
	wire _w6631_ ;
	wire _w6632_ ;
	wire _w6633_ ;
	wire _w6634_ ;
	wire _w6635_ ;
	wire _w6636_ ;
	wire _w6637_ ;
	wire _w6638_ ;
	wire _w6639_ ;
	wire _w6640_ ;
	wire _w6641_ ;
	wire _w6642_ ;
	wire _w6643_ ;
	wire _w6644_ ;
	wire _w6645_ ;
	wire _w6646_ ;
	wire _w6647_ ;
	wire _w6648_ ;
	wire _w6649_ ;
	wire _w6650_ ;
	wire _w6651_ ;
	wire _w6652_ ;
	wire _w6653_ ;
	wire _w6654_ ;
	wire _w6655_ ;
	wire _w6656_ ;
	wire _w6657_ ;
	wire _w6658_ ;
	wire _w6659_ ;
	wire _w6660_ ;
	wire _w6661_ ;
	wire _w6662_ ;
	wire _w6663_ ;
	wire _w6664_ ;
	wire _w6665_ ;
	wire _w6666_ ;
	wire _w6667_ ;
	wire _w6668_ ;
	wire _w6669_ ;
	wire _w6670_ ;
	wire _w6671_ ;
	wire _w6672_ ;
	wire _w6673_ ;
	wire _w6674_ ;
	wire _w6675_ ;
	wire _w6676_ ;
	wire _w6677_ ;
	wire _w6678_ ;
	wire _w6679_ ;
	wire _w6680_ ;
	wire _w6681_ ;
	wire _w6682_ ;
	wire _w6683_ ;
	wire _w6684_ ;
	wire _w6685_ ;
	wire _w6686_ ;
	wire _w6687_ ;
	wire _w6688_ ;
	wire _w6689_ ;
	wire _w6690_ ;
	wire _w6691_ ;
	wire _w6692_ ;
	wire _w6693_ ;
	wire _w6694_ ;
	wire _w6695_ ;
	wire _w6696_ ;
	wire _w6697_ ;
	wire _w6698_ ;
	wire _w6699_ ;
	wire _w6700_ ;
	wire _w6701_ ;
	wire _w6702_ ;
	wire _w6703_ ;
	wire _w6704_ ;
	wire _w6705_ ;
	wire _w6706_ ;
	wire _w6707_ ;
	wire _w6708_ ;
	wire _w6709_ ;
	wire _w6710_ ;
	wire _w6711_ ;
	wire _w6712_ ;
	wire _w6713_ ;
	wire _w6714_ ;
	wire _w6715_ ;
	wire _w6716_ ;
	wire _w6717_ ;
	wire _w6718_ ;
	wire _w6719_ ;
	wire _w6720_ ;
	wire _w6721_ ;
	wire _w6722_ ;
	wire _w6723_ ;
	wire _w6724_ ;
	wire _w6725_ ;
	wire _w6726_ ;
	wire _w6727_ ;
	wire _w6728_ ;
	wire _w6729_ ;
	wire _w6730_ ;
	wire _w6731_ ;
	wire _w6732_ ;
	wire _w6733_ ;
	wire _w6734_ ;
	wire _w6735_ ;
	wire _w6736_ ;
	wire _w6737_ ;
	wire _w6738_ ;
	wire _w6739_ ;
	wire _w6740_ ;
	wire _w6741_ ;
	wire _w6742_ ;
	wire _w6743_ ;
	wire _w6744_ ;
	wire _w6745_ ;
	wire _w6746_ ;
	wire _w6747_ ;
	wire _w6748_ ;
	wire _w6749_ ;
	wire _w6750_ ;
	wire _w6751_ ;
	wire _w6752_ ;
	wire _w6753_ ;
	wire _w6754_ ;
	wire _w6755_ ;
	wire _w6756_ ;
	wire _w6757_ ;
	wire _w6758_ ;
	wire _w6759_ ;
	wire _w6760_ ;
	wire _w6761_ ;
	wire _w6762_ ;
	wire _w6763_ ;
	wire _w6764_ ;
	wire _w6765_ ;
	wire _w6766_ ;
	wire _w6767_ ;
	wire _w6768_ ;
	wire _w6769_ ;
	wire _w6770_ ;
	wire _w6771_ ;
	wire _w6772_ ;
	wire _w6773_ ;
	wire _w6774_ ;
	wire _w6775_ ;
	wire _w6776_ ;
	wire _w6777_ ;
	wire _w6778_ ;
	wire _w6779_ ;
	wire _w6780_ ;
	wire _w6781_ ;
	wire _w6782_ ;
	wire _w6783_ ;
	wire _w6784_ ;
	wire _w6785_ ;
	wire _w6786_ ;
	wire _w6787_ ;
	wire _w6788_ ;
	wire _w6789_ ;
	wire _w6790_ ;
	wire _w6791_ ;
	wire _w6792_ ;
	wire _w6793_ ;
	wire _w6794_ ;
	wire _w6795_ ;
	wire _w6796_ ;
	wire _w6797_ ;
	wire _w6798_ ;
	wire _w6799_ ;
	wire _w6800_ ;
	wire _w6801_ ;
	wire _w6802_ ;
	wire _w6803_ ;
	wire _w6804_ ;
	wire _w6805_ ;
	wire _w6806_ ;
	wire _w6807_ ;
	wire _w6808_ ;
	wire _w6809_ ;
	wire _w6810_ ;
	wire _w6811_ ;
	wire _w6812_ ;
	wire _w6813_ ;
	wire _w6814_ ;
	wire _w6815_ ;
	wire _w6816_ ;
	wire _w6817_ ;
	wire _w6818_ ;
	wire _w6819_ ;
	wire _w6820_ ;
	wire _w6821_ ;
	wire _w6822_ ;
	wire _w6823_ ;
	wire _w6824_ ;
	wire _w6825_ ;
	wire _w6826_ ;
	wire _w6827_ ;
	wire _w6828_ ;
	wire _w6829_ ;
	wire _w6830_ ;
	wire _w6831_ ;
	wire _w6832_ ;
	wire _w6833_ ;
	wire _w6834_ ;
	wire _w6835_ ;
	wire _w6836_ ;
	wire _w6837_ ;
	wire _w6838_ ;
	wire _w6839_ ;
	wire _w6840_ ;
	wire _w6841_ ;
	wire _w6842_ ;
	wire _w6843_ ;
	wire _w6844_ ;
	wire _w6845_ ;
	wire _w6846_ ;
	wire _w6847_ ;
	wire _w6848_ ;
	wire _w6849_ ;
	wire _w6850_ ;
	wire _w6851_ ;
	wire _w6852_ ;
	wire _w6853_ ;
	wire _w6854_ ;
	wire _w6855_ ;
	wire _w6856_ ;
	wire _w6857_ ;
	wire _w6858_ ;
	wire _w6859_ ;
	wire _w6860_ ;
	wire _w6861_ ;
	wire _w6862_ ;
	wire _w6863_ ;
	wire _w6864_ ;
	wire _w6865_ ;
	wire _w6866_ ;
	wire _w6867_ ;
	wire _w6868_ ;
	wire _w6869_ ;
	wire _w6870_ ;
	wire _w6871_ ;
	wire _w6872_ ;
	wire _w6873_ ;
	wire _w6874_ ;
	wire _w6875_ ;
	wire _w6876_ ;
	wire _w6877_ ;
	wire _w6878_ ;
	wire _w6879_ ;
	wire _w6880_ ;
	wire _w6881_ ;
	wire _w6882_ ;
	wire _w6883_ ;
	wire _w6884_ ;
	wire _w6885_ ;
	wire _w6886_ ;
	wire _w6887_ ;
	wire _w6888_ ;
	wire _w6889_ ;
	wire _w6890_ ;
	wire _w6891_ ;
	wire _w6892_ ;
	wire _w6893_ ;
	wire _w6894_ ;
	wire _w6895_ ;
	wire _w6896_ ;
	wire _w6897_ ;
	wire _w6898_ ;
	wire _w6899_ ;
	wire _w6900_ ;
	wire _w6901_ ;
	wire _w6902_ ;
	wire _w6903_ ;
	wire _w6904_ ;
	wire _w6905_ ;
	wire _w6906_ ;
	wire _w6907_ ;
	wire _w6908_ ;
	wire _w6909_ ;
	wire _w6910_ ;
	wire _w6911_ ;
	wire _w6912_ ;
	wire _w6913_ ;
	wire _w6914_ ;
	wire _w6915_ ;
	wire _w6916_ ;
	wire _w6917_ ;
	wire _w6918_ ;
	wire _w6919_ ;
	wire _w6920_ ;
	wire _w6921_ ;
	wire _w6922_ ;
	wire _w6923_ ;
	wire _w6924_ ;
	wire _w6925_ ;
	wire _w6926_ ;
	wire _w6927_ ;
	wire _w6928_ ;
	wire _w6929_ ;
	wire _w6930_ ;
	wire _w6931_ ;
	wire _w6932_ ;
	wire _w6933_ ;
	wire _w6934_ ;
	wire _w6935_ ;
	wire _w6936_ ;
	wire _w6937_ ;
	wire _w6938_ ;
	wire _w6939_ ;
	wire _w6940_ ;
	wire _w6941_ ;
	wire _w6942_ ;
	wire _w6943_ ;
	wire _w6944_ ;
	wire _w6945_ ;
	wire _w6946_ ;
	wire _w6947_ ;
	wire _w6948_ ;
	wire _w6949_ ;
	wire _w6950_ ;
	wire _w6951_ ;
	wire _w6952_ ;
	wire _w6953_ ;
	wire _w6954_ ;
	wire _w6955_ ;
	wire _w6956_ ;
	wire _w6957_ ;
	wire _w6958_ ;
	wire _w6959_ ;
	wire _w6960_ ;
	wire _w6961_ ;
	wire _w6962_ ;
	wire _w6963_ ;
	wire _w6964_ ;
	wire _w6965_ ;
	wire _w6966_ ;
	wire _w6967_ ;
	wire _w6968_ ;
	wire _w6969_ ;
	wire _w6970_ ;
	wire _w6971_ ;
	wire _w6972_ ;
	wire _w6973_ ;
	wire _w6974_ ;
	wire _w6975_ ;
	wire _w6976_ ;
	wire _w6977_ ;
	wire _w6978_ ;
	wire _w6979_ ;
	wire _w6980_ ;
	wire _w6981_ ;
	wire _w6982_ ;
	wire _w6983_ ;
	wire _w6984_ ;
	wire _w6985_ ;
	wire _w6986_ ;
	wire _w6987_ ;
	wire _w6988_ ;
	wire _w6989_ ;
	wire _w6990_ ;
	wire _w6991_ ;
	wire _w6992_ ;
	wire _w6993_ ;
	wire _w6994_ ;
	wire _w6995_ ;
	wire _w6996_ ;
	wire _w6997_ ;
	wire _w6998_ ;
	wire _w6999_ ;
	wire _w7000_ ;
	wire _w7001_ ;
	wire _w7002_ ;
	wire _w7003_ ;
	wire _w7004_ ;
	wire _w7005_ ;
	wire _w7006_ ;
	wire _w7007_ ;
	wire _w7008_ ;
	wire _w7009_ ;
	wire _w7010_ ;
	wire _w7011_ ;
	wire _w7012_ ;
	wire _w7013_ ;
	wire _w7014_ ;
	wire _w7015_ ;
	wire _w7016_ ;
	wire _w7017_ ;
	wire _w7018_ ;
	wire _w7019_ ;
	wire _w7020_ ;
	wire _w7021_ ;
	wire _w7022_ ;
	wire _w7023_ ;
	wire _w7024_ ;
	wire _w7025_ ;
	wire _w7026_ ;
	wire _w7027_ ;
	wire _w7028_ ;
	wire _w7029_ ;
	wire _w7030_ ;
	wire _w7031_ ;
	wire _w7032_ ;
	wire _w7033_ ;
	wire _w7034_ ;
	wire _w7035_ ;
	wire _w7036_ ;
	wire _w7037_ ;
	wire _w7038_ ;
	wire _w7039_ ;
	wire _w7040_ ;
	wire _w7041_ ;
	wire _w7042_ ;
	wire _w7043_ ;
	wire _w7044_ ;
	wire _w7045_ ;
	wire _w7046_ ;
	wire _w7047_ ;
	wire _w7048_ ;
	wire _w7049_ ;
	wire _w7050_ ;
	wire _w7051_ ;
	wire _w7052_ ;
	wire _w7053_ ;
	wire _w7054_ ;
	wire _w7055_ ;
	wire _w7056_ ;
	wire _w7057_ ;
	wire _w7058_ ;
	wire _w7059_ ;
	wire _w7060_ ;
	wire _w7061_ ;
	wire _w7062_ ;
	wire _w7063_ ;
	wire _w7064_ ;
	wire _w7065_ ;
	wire _w7066_ ;
	wire _w7067_ ;
	wire _w7068_ ;
	wire _w7069_ ;
	wire _w7070_ ;
	wire _w7071_ ;
	wire _w7072_ ;
	wire _w7073_ ;
	wire _w7074_ ;
	wire _w7075_ ;
	wire _w7076_ ;
	wire _w7077_ ;
	wire _w7078_ ;
	wire _w7079_ ;
	wire _w7080_ ;
	wire _w7081_ ;
	wire _w7082_ ;
	wire _w7083_ ;
	wire _w7084_ ;
	wire _w7085_ ;
	wire _w7086_ ;
	wire _w7087_ ;
	wire _w7088_ ;
	wire _w7089_ ;
	wire _w7090_ ;
	wire _w7091_ ;
	wire _w7092_ ;
	wire _w7093_ ;
	wire _w7094_ ;
	wire _w7095_ ;
	wire _w7096_ ;
	wire _w7097_ ;
	wire _w7098_ ;
	wire _w7099_ ;
	wire _w7100_ ;
	wire _w7101_ ;
	wire _w7102_ ;
	wire _w7103_ ;
	wire _w7104_ ;
	wire _w7105_ ;
	wire _w7106_ ;
	wire _w7107_ ;
	wire _w7108_ ;
	wire _w7109_ ;
	wire _w7110_ ;
	wire _w7111_ ;
	wire _w7112_ ;
	wire _w7113_ ;
	wire _w7114_ ;
	wire _w7115_ ;
	wire _w7116_ ;
	wire _w7117_ ;
	wire _w7118_ ;
	wire _w7119_ ;
	wire _w7120_ ;
	wire _w7121_ ;
	wire _w7122_ ;
	wire _w7123_ ;
	wire _w7124_ ;
	wire _w7125_ ;
	wire _w7126_ ;
	wire _w7127_ ;
	wire _w7128_ ;
	wire _w7129_ ;
	wire _w7130_ ;
	wire _w7131_ ;
	wire _w7132_ ;
	wire _w7133_ ;
	wire _w7134_ ;
	wire _w7135_ ;
	wire _w7136_ ;
	wire _w7137_ ;
	wire _w7138_ ;
	wire _w7139_ ;
	wire _w7140_ ;
	wire _w7141_ ;
	wire _w7142_ ;
	wire _w7143_ ;
	wire _w7144_ ;
	wire _w7145_ ;
	wire _w7146_ ;
	wire _w7147_ ;
	wire _w7148_ ;
	wire _w7149_ ;
	wire _w7150_ ;
	wire _w7151_ ;
	wire _w7152_ ;
	wire _w7153_ ;
	wire _w7154_ ;
	wire _w7155_ ;
	wire _w7156_ ;
	wire _w7157_ ;
	wire _w7158_ ;
	wire _w7159_ ;
	wire _w7160_ ;
	wire _w7161_ ;
	wire _w7162_ ;
	wire _w7163_ ;
	wire _w7164_ ;
	wire _w7165_ ;
	wire _w7166_ ;
	wire _w7167_ ;
	wire _w7168_ ;
	wire _w7169_ ;
	wire _w7170_ ;
	wire _w7171_ ;
	wire _w7172_ ;
	wire _w7173_ ;
	wire _w7174_ ;
	wire _w7175_ ;
	wire _w7176_ ;
	wire _w7177_ ;
	wire _w7178_ ;
	wire _w7179_ ;
	wire _w7180_ ;
	wire _w7181_ ;
	wire _w7182_ ;
	wire _w7183_ ;
	wire _w7184_ ;
	wire _w7185_ ;
	wire _w7186_ ;
	wire _w7187_ ;
	wire _w7188_ ;
	wire _w7189_ ;
	wire _w7190_ ;
	wire _w7191_ ;
	wire _w7192_ ;
	wire _w7193_ ;
	wire _w7194_ ;
	wire _w7195_ ;
	wire _w7196_ ;
	wire _w7197_ ;
	wire _w7198_ ;
	wire _w7199_ ;
	wire _w7200_ ;
	wire _w7201_ ;
	wire _w7202_ ;
	wire _w7203_ ;
	wire _w7204_ ;
	wire _w7205_ ;
	wire _w7206_ ;
	wire _w7207_ ;
	wire _w7208_ ;
	wire _w7209_ ;
	wire _w7210_ ;
	wire _w7211_ ;
	wire _w7212_ ;
	wire _w7213_ ;
	wire _w7214_ ;
	wire _w7215_ ;
	wire _w7216_ ;
	wire _w7217_ ;
	wire _w7218_ ;
	wire _w7219_ ;
	wire _w7220_ ;
	wire _w7221_ ;
	wire _w7222_ ;
	wire _w7223_ ;
	wire _w7224_ ;
	wire _w7225_ ;
	wire _w7226_ ;
	wire _w7227_ ;
	wire _w7228_ ;
	wire _w7229_ ;
	wire _w7230_ ;
	wire _w7231_ ;
	wire _w7232_ ;
	wire _w7233_ ;
	wire _w7234_ ;
	wire _w7235_ ;
	wire _w7236_ ;
	wire _w7237_ ;
	wire _w7238_ ;
	wire _w7239_ ;
	wire _w7240_ ;
	wire _w7241_ ;
	wire _w7242_ ;
	wire _w7243_ ;
	wire _w7244_ ;
	wire _w7245_ ;
	wire _w7246_ ;
	wire _w7247_ ;
	wire _w7248_ ;
	wire _w7249_ ;
	wire _w7250_ ;
	wire _w7251_ ;
	wire _w7252_ ;
	wire _w7253_ ;
	wire _w7254_ ;
	wire _w7255_ ;
	wire _w7256_ ;
	wire _w7257_ ;
	wire _w7258_ ;
	wire _w7259_ ;
	wire _w7260_ ;
	wire _w7261_ ;
	wire _w7262_ ;
	wire _w7263_ ;
	wire _w7264_ ;
	wire _w7265_ ;
	wire _w7266_ ;
	wire _w7267_ ;
	wire _w7268_ ;
	wire _w7269_ ;
	wire _w7270_ ;
	wire _w7271_ ;
	wire _w7272_ ;
	wire _w7273_ ;
	wire _w7274_ ;
	wire _w7275_ ;
	wire _w7276_ ;
	wire _w7277_ ;
	wire _w7278_ ;
	wire _w7279_ ;
	wire _w7280_ ;
	wire _w7281_ ;
	wire _w7282_ ;
	wire _w7283_ ;
	wire _w7284_ ;
	wire _w7285_ ;
	wire _w7286_ ;
	wire _w7287_ ;
	wire _w7288_ ;
	wire _w7289_ ;
	wire _w7290_ ;
	wire _w7291_ ;
	wire _w7292_ ;
	wire _w7293_ ;
	wire _w7294_ ;
	wire _w7295_ ;
	wire _w7296_ ;
	wire _w7297_ ;
	wire _w7298_ ;
	wire _w7299_ ;
	wire _w7300_ ;
	wire _w7301_ ;
	wire _w7302_ ;
	wire _w7303_ ;
	wire _w7304_ ;
	wire _w7305_ ;
	wire _w7306_ ;
	wire _w7307_ ;
	wire _w7308_ ;
	wire _w7309_ ;
	wire _w7310_ ;
	wire _w7311_ ;
	wire _w7312_ ;
	wire _w7313_ ;
	wire _w7314_ ;
	wire _w7315_ ;
	wire _w7316_ ;
	wire _w7317_ ;
	wire _w7318_ ;
	wire _w7319_ ;
	wire _w7320_ ;
	wire _w7321_ ;
	wire _w7322_ ;
	wire _w7323_ ;
	wire _w7324_ ;
	wire _w7325_ ;
	wire _w7326_ ;
	wire _w7327_ ;
	wire _w7328_ ;
	wire _w7329_ ;
	wire _w7330_ ;
	wire _w7331_ ;
	wire _w7332_ ;
	wire _w7333_ ;
	wire _w7334_ ;
	wire _w7335_ ;
	wire _w7336_ ;
	wire _w7337_ ;
	wire _w7338_ ;
	wire _w7339_ ;
	wire _w7340_ ;
	wire _w7341_ ;
	wire _w7342_ ;
	wire _w7343_ ;
	wire _w7344_ ;
	wire _w7345_ ;
	wire _w7346_ ;
	wire _w7347_ ;
	wire _w7348_ ;
	wire _w7349_ ;
	wire _w7350_ ;
	wire _w7351_ ;
	wire _w7352_ ;
	wire _w7353_ ;
	wire _w7354_ ;
	wire _w7355_ ;
	wire _w7356_ ;
	wire _w7357_ ;
	wire _w7358_ ;
	wire _w7359_ ;
	wire _w7360_ ;
	wire _w7361_ ;
	wire _w7362_ ;
	wire _w7363_ ;
	wire _w7364_ ;
	wire _w7365_ ;
	wire _w7366_ ;
	wire _w7367_ ;
	wire _w7368_ ;
	wire _w7369_ ;
	wire _w7370_ ;
	wire _w7371_ ;
	wire _w7372_ ;
	wire _w7373_ ;
	wire _w7374_ ;
	wire _w7375_ ;
	wire _w7376_ ;
	wire _w7377_ ;
	wire _w7378_ ;
	wire _w7379_ ;
	wire _w7380_ ;
	wire _w7381_ ;
	wire _w7382_ ;
	wire _w7383_ ;
	wire _w7384_ ;
	wire _w7385_ ;
	wire _w7386_ ;
	wire _w7387_ ;
	wire _w7388_ ;
	wire _w7389_ ;
	wire _w7390_ ;
	wire _w7391_ ;
	wire _w7392_ ;
	wire _w7393_ ;
	wire _w7394_ ;
	wire _w7395_ ;
	wire _w7396_ ;
	wire _w7397_ ;
	wire _w7398_ ;
	wire _w7399_ ;
	wire _w7400_ ;
	wire _w7401_ ;
	wire _w7402_ ;
	wire _w7403_ ;
	wire _w7404_ ;
	wire _w7405_ ;
	wire _w7406_ ;
	wire _w7407_ ;
	wire _w7408_ ;
	wire _w7409_ ;
	wire _w7410_ ;
	wire _w7411_ ;
	wire _w7412_ ;
	wire _w7413_ ;
	wire _w7414_ ;
	wire _w7415_ ;
	wire _w7416_ ;
	wire _w7417_ ;
	wire _w7418_ ;
	wire _w7419_ ;
	wire _w7420_ ;
	wire _w7421_ ;
	wire _w7422_ ;
	wire _w7423_ ;
	wire _w7424_ ;
	wire _w7425_ ;
	wire _w7426_ ;
	wire _w7427_ ;
	wire _w7428_ ;
	wire _w7429_ ;
	wire _w7430_ ;
	wire _w7431_ ;
	wire _w7432_ ;
	wire _w7433_ ;
	wire _w7434_ ;
	wire _w7435_ ;
	wire _w7436_ ;
	wire _w7437_ ;
	wire _w7438_ ;
	wire _w7439_ ;
	wire _w7440_ ;
	wire _w7441_ ;
	wire _w7442_ ;
	wire _w7443_ ;
	wire _w7444_ ;
	wire _w7445_ ;
	wire _w7446_ ;
	wire _w7447_ ;
	wire _w7448_ ;
	wire _w7449_ ;
	wire _w7450_ ;
	wire _w7451_ ;
	wire _w7452_ ;
	wire _w7453_ ;
	wire _w7454_ ;
	wire _w7455_ ;
	wire _w7456_ ;
	wire _w7457_ ;
	wire _w7458_ ;
	wire _w7459_ ;
	wire _w7460_ ;
	wire _w7461_ ;
	wire _w7462_ ;
	wire _w7463_ ;
	wire _w7464_ ;
	wire _w7465_ ;
	wire _w7466_ ;
	wire _w7467_ ;
	wire _w7468_ ;
	wire _w7469_ ;
	wire _w7470_ ;
	wire _w7471_ ;
	wire _w7472_ ;
	wire _w7473_ ;
	wire _w7474_ ;
	wire _w7475_ ;
	wire _w7476_ ;
	wire _w7477_ ;
	wire _w7478_ ;
	wire _w7479_ ;
	wire _w7480_ ;
	wire _w7481_ ;
	wire _w7482_ ;
	wire _w7483_ ;
	wire _w7484_ ;
	wire _w7485_ ;
	wire _w7486_ ;
	wire _w7487_ ;
	wire _w7488_ ;
	wire _w7489_ ;
	wire _w7490_ ;
	wire _w7491_ ;
	wire _w7492_ ;
	wire _w7493_ ;
	wire _w7494_ ;
	wire _w7495_ ;
	wire _w7496_ ;
	wire _w7497_ ;
	wire _w7498_ ;
	wire _w7499_ ;
	wire _w7500_ ;
	wire _w7501_ ;
	wire _w7502_ ;
	wire _w7503_ ;
	wire _w7504_ ;
	wire _w7505_ ;
	wire _w7506_ ;
	wire _w7507_ ;
	wire _w7508_ ;
	wire _w7509_ ;
	wire _w7510_ ;
	wire _w7511_ ;
	wire _w7512_ ;
	wire _w7513_ ;
	wire _w7514_ ;
	wire _w7515_ ;
	wire _w7516_ ;
	wire _w7517_ ;
	wire _w7518_ ;
	wire _w7519_ ;
	wire _w7520_ ;
	wire _w7521_ ;
	wire _w7522_ ;
	wire _w7523_ ;
	wire _w7524_ ;
	wire _w7525_ ;
	wire _w7526_ ;
	wire _w7527_ ;
	wire _w7528_ ;
	wire _w7529_ ;
	wire _w7530_ ;
	wire _w7531_ ;
	wire _w7532_ ;
	wire _w7533_ ;
	wire _w7534_ ;
	wire _w7535_ ;
	wire _w7536_ ;
	wire _w7537_ ;
	wire _w7538_ ;
	wire _w7539_ ;
	wire _w7540_ ;
	wire _w7541_ ;
	wire _w7542_ ;
	wire _w7543_ ;
	wire _w7544_ ;
	wire _w7545_ ;
	wire _w7546_ ;
	wire _w7547_ ;
	wire _w7548_ ;
	wire _w7549_ ;
	wire _w7550_ ;
	wire _w7551_ ;
	wire _w7552_ ;
	wire _w7553_ ;
	wire _w7554_ ;
	wire _w7555_ ;
	wire _w7556_ ;
	wire _w7557_ ;
	wire _w7558_ ;
	wire _w7559_ ;
	wire _w7560_ ;
	wire _w7561_ ;
	wire _w7562_ ;
	wire _w7563_ ;
	wire _w7564_ ;
	wire _w7565_ ;
	wire _w7566_ ;
	wire _w7567_ ;
	wire _w7568_ ;
	wire _w7569_ ;
	wire _w7570_ ;
	wire _w7571_ ;
	wire _w7572_ ;
	wire _w7573_ ;
	wire _w7574_ ;
	wire _w7575_ ;
	wire _w7576_ ;
	wire _w7577_ ;
	wire _w7578_ ;
	wire _w7579_ ;
	wire _w7580_ ;
	wire _w7581_ ;
	wire _w7582_ ;
	wire _w7583_ ;
	wire _w7584_ ;
	wire _w7585_ ;
	wire _w7586_ ;
	wire _w7587_ ;
	wire _w7588_ ;
	wire _w7589_ ;
	wire _w7590_ ;
	wire _w7591_ ;
	wire _w7592_ ;
	wire _w7593_ ;
	wire _w7594_ ;
	wire _w7595_ ;
	wire _w7596_ ;
	wire _w7597_ ;
	wire _w7598_ ;
	wire _w7599_ ;
	wire _w7600_ ;
	wire _w7601_ ;
	wire _w7602_ ;
	wire _w7603_ ;
	wire _w7604_ ;
	wire _w7605_ ;
	wire _w7606_ ;
	wire _w7607_ ;
	wire _w7608_ ;
	wire _w7609_ ;
	wire _w7610_ ;
	wire _w7611_ ;
	wire _w7612_ ;
	wire _w7613_ ;
	wire _w7614_ ;
	wire _w7615_ ;
	wire _w7616_ ;
	wire _w7617_ ;
	wire _w7618_ ;
	wire _w7619_ ;
	wire _w7620_ ;
	wire _w7621_ ;
	wire _w7622_ ;
	wire _w7623_ ;
	wire _w7624_ ;
	wire _w7625_ ;
	wire _w7626_ ;
	wire _w7627_ ;
	wire _w7628_ ;
	wire _w7629_ ;
	wire _w7630_ ;
	wire _w7631_ ;
	wire _w7632_ ;
	wire _w7633_ ;
	wire _w7634_ ;
	wire _w7635_ ;
	wire _w7636_ ;
	wire _w7637_ ;
	wire _w7638_ ;
	wire _w7639_ ;
	wire _w7640_ ;
	wire _w7641_ ;
	wire _w7642_ ;
	wire _w7643_ ;
	wire _w7644_ ;
	wire _w7645_ ;
	wire _w7646_ ;
	wire _w7647_ ;
	wire _w7648_ ;
	wire _w7649_ ;
	wire _w7650_ ;
	wire _w7651_ ;
	wire _w7652_ ;
	wire _w7653_ ;
	wire _w7654_ ;
	wire _w7655_ ;
	wire _w7656_ ;
	wire _w7657_ ;
	wire _w7658_ ;
	wire _w7659_ ;
	wire _w7660_ ;
	wire _w7661_ ;
	wire _w7662_ ;
	wire _w7663_ ;
	wire _w7664_ ;
	wire _w7665_ ;
	wire _w7666_ ;
	wire _w7667_ ;
	wire _w7668_ ;
	wire _w7669_ ;
	wire _w7670_ ;
	wire _w7671_ ;
	wire _w7672_ ;
	wire _w7673_ ;
	wire _w7674_ ;
	wire _w7675_ ;
	wire _w7676_ ;
	wire _w7677_ ;
	wire _w7678_ ;
	wire _w7679_ ;
	wire _w7680_ ;
	wire _w7681_ ;
	wire _w7682_ ;
	wire _w7683_ ;
	wire _w7684_ ;
	wire _w7685_ ;
	wire _w7686_ ;
	wire _w7687_ ;
	wire _w7688_ ;
	wire _w7689_ ;
	wire _w7690_ ;
	wire _w7691_ ;
	wire _w7692_ ;
	wire _w7693_ ;
	wire _w7694_ ;
	wire _w7695_ ;
	wire _w7696_ ;
	wire _w7697_ ;
	wire _w7698_ ;
	wire _w7699_ ;
	wire _w7700_ ;
	wire _w7701_ ;
	wire _w7702_ ;
	wire _w7703_ ;
	wire _w7704_ ;
	wire _w7705_ ;
	wire _w7706_ ;
	wire _w7707_ ;
	wire _w7708_ ;
	wire _w7709_ ;
	wire _w7710_ ;
	wire _w7711_ ;
	wire _w7712_ ;
	wire _w7713_ ;
	wire _w7714_ ;
	wire _w7715_ ;
	wire _w7716_ ;
	wire _w7717_ ;
	wire _w7718_ ;
	wire _w7719_ ;
	wire _w7720_ ;
	wire _w7721_ ;
	wire _w7722_ ;
	wire _w7723_ ;
	wire _w7724_ ;
	wire _w7725_ ;
	wire _w7726_ ;
	wire _w7727_ ;
	wire _w7728_ ;
	wire _w7729_ ;
	wire _w7730_ ;
	wire _w7731_ ;
	wire _w7732_ ;
	wire _w7733_ ;
	wire _w7734_ ;
	wire _w7735_ ;
	wire _w7736_ ;
	wire _w7737_ ;
	wire _w7738_ ;
	wire _w7739_ ;
	wire _w7740_ ;
	wire _w7741_ ;
	wire _w7742_ ;
	wire _w7743_ ;
	wire _w7744_ ;
	wire _w7745_ ;
	wire _w7746_ ;
	wire _w7747_ ;
	wire _w7748_ ;
	wire _w7749_ ;
	wire _w7750_ ;
	wire _w7751_ ;
	wire _w7752_ ;
	wire _w7753_ ;
	wire _w7754_ ;
	wire _w7755_ ;
	wire _w7756_ ;
	wire _w7757_ ;
	wire _w7758_ ;
	wire _w7759_ ;
	wire _w7760_ ;
	wire _w7761_ ;
	wire _w7762_ ;
	wire _w7763_ ;
	wire _w7764_ ;
	wire _w7765_ ;
	wire _w7766_ ;
	wire _w7767_ ;
	wire _w7768_ ;
	wire _w7769_ ;
	wire _w7770_ ;
	wire _w7771_ ;
	wire _w7772_ ;
	wire _w7773_ ;
	wire _w7774_ ;
	wire _w7775_ ;
	wire _w7776_ ;
	wire _w7777_ ;
	wire _w7778_ ;
	wire _w7779_ ;
	wire _w7780_ ;
	wire _w7781_ ;
	wire _w7782_ ;
	wire _w7783_ ;
	wire _w7784_ ;
	wire _w7785_ ;
	wire _w7786_ ;
	wire _w7787_ ;
	wire _w7788_ ;
	wire _w7789_ ;
	wire _w7790_ ;
	wire _w7791_ ;
	wire _w7792_ ;
	wire _w7793_ ;
	wire _w7794_ ;
	wire _w7795_ ;
	wire _w7796_ ;
	wire _w7797_ ;
	wire _w7798_ ;
	wire _w7799_ ;
	wire _w7800_ ;
	wire _w7801_ ;
	wire _w7802_ ;
	wire _w7803_ ;
	wire _w7804_ ;
	wire _w7805_ ;
	wire _w7806_ ;
	wire _w7807_ ;
	wire _w7808_ ;
	wire _w7809_ ;
	wire _w7810_ ;
	wire _w7811_ ;
	wire _w7812_ ;
	wire _w7813_ ;
	wire _w7814_ ;
	wire _w7815_ ;
	wire _w7816_ ;
	wire _w7817_ ;
	wire _w7818_ ;
	wire _w7819_ ;
	wire _w7820_ ;
	wire _w7821_ ;
	wire _w7822_ ;
	wire _w7823_ ;
	wire _w7824_ ;
	wire _w7825_ ;
	wire _w7826_ ;
	wire _w7827_ ;
	wire _w7828_ ;
	wire _w7829_ ;
	wire _w7830_ ;
	wire _w7831_ ;
	wire _w7832_ ;
	wire _w7833_ ;
	wire _w7834_ ;
	wire _w7835_ ;
	wire _w7836_ ;
	wire _w7837_ ;
	wire _w7838_ ;
	wire _w7839_ ;
	wire _w7840_ ;
	wire _w7841_ ;
	wire _w7842_ ;
	wire _w7843_ ;
	wire _w7844_ ;
	wire _w7845_ ;
	wire _w7846_ ;
	wire _w7847_ ;
	wire _w7848_ ;
	wire _w7849_ ;
	wire _w7850_ ;
	wire _w7851_ ;
	wire _w7852_ ;
	wire _w7853_ ;
	wire _w7854_ ;
	wire _w7855_ ;
	wire _w7856_ ;
	wire _w7857_ ;
	wire _w7858_ ;
	wire _w7859_ ;
	wire _w7860_ ;
	wire _w7861_ ;
	wire _w7862_ ;
	wire _w7863_ ;
	wire _w7864_ ;
	wire _w7865_ ;
	wire _w7866_ ;
	wire _w7867_ ;
	wire _w7868_ ;
	wire _w7869_ ;
	wire _w7870_ ;
	wire _w7871_ ;
	wire _w7872_ ;
	wire _w7873_ ;
	wire _w7874_ ;
	wire _w7875_ ;
	wire _w7876_ ;
	wire _w7877_ ;
	wire _w7878_ ;
	wire _w7879_ ;
	wire _w7880_ ;
	wire _w7881_ ;
	wire _w7882_ ;
	wire _w7883_ ;
	wire _w7884_ ;
	wire _w7885_ ;
	wire _w7886_ ;
	wire _w7887_ ;
	wire _w7888_ ;
	wire _w7889_ ;
	wire _w7890_ ;
	wire _w7891_ ;
	wire _w7892_ ;
	wire _w7893_ ;
	wire _w7894_ ;
	wire _w7895_ ;
	wire _w7896_ ;
	wire _w7897_ ;
	wire _w7898_ ;
	wire _w7899_ ;
	wire _w7900_ ;
	wire _w7901_ ;
	wire _w7902_ ;
	wire _w7903_ ;
	wire _w7904_ ;
	wire _w7905_ ;
	wire _w7906_ ;
	wire _w7907_ ;
	wire _w7908_ ;
	wire _w7909_ ;
	wire _w7910_ ;
	wire _w7911_ ;
	wire _w7912_ ;
	wire _w7913_ ;
	wire _w7914_ ;
	wire _w7915_ ;
	wire _w7916_ ;
	wire _w7917_ ;
	wire _w7918_ ;
	wire _w7919_ ;
	wire _w7920_ ;
	wire _w7921_ ;
	wire _w7922_ ;
	wire _w7923_ ;
	wire _w7924_ ;
	wire _w7925_ ;
	wire _w7926_ ;
	wire _w7927_ ;
	wire _w7928_ ;
	wire _w7929_ ;
	wire _w7930_ ;
	wire _w7931_ ;
	wire _w7932_ ;
	wire _w7933_ ;
	wire _w7934_ ;
	wire _w7935_ ;
	wire _w7936_ ;
	wire _w7937_ ;
	wire _w7938_ ;
	wire _w7939_ ;
	wire _w7940_ ;
	wire _w7941_ ;
	wire _w7942_ ;
	wire _w7943_ ;
	wire _w7944_ ;
	wire _w7945_ ;
	wire _w7946_ ;
	wire _w7947_ ;
	wire _w7948_ ;
	wire _w7949_ ;
	wire _w7950_ ;
	wire _w7951_ ;
	wire _w7952_ ;
	wire _w7953_ ;
	wire _w7954_ ;
	wire _w7955_ ;
	wire _w7956_ ;
	wire _w7957_ ;
	wire _w7958_ ;
	wire _w7959_ ;
	wire _w7960_ ;
	wire _w7961_ ;
	wire _w7962_ ;
	wire _w7963_ ;
	wire _w7964_ ;
	wire _w7965_ ;
	wire _w7966_ ;
	wire _w7967_ ;
	wire _w7968_ ;
	wire _w7969_ ;
	wire _w7970_ ;
	wire _w7971_ ;
	wire _w7972_ ;
	wire _w7973_ ;
	wire _w7974_ ;
	wire _w7975_ ;
	wire _w7976_ ;
	wire _w7977_ ;
	wire _w7978_ ;
	wire _w7979_ ;
	wire _w7980_ ;
	wire _w7981_ ;
	wire _w7982_ ;
	wire _w7983_ ;
	wire _w7984_ ;
	wire _w7985_ ;
	wire _w7986_ ;
	wire _w7987_ ;
	wire _w7988_ ;
	wire _w7989_ ;
	wire _w7990_ ;
	wire _w7991_ ;
	wire _w7992_ ;
	wire _w7993_ ;
	wire _w7994_ ;
	wire _w7995_ ;
	wire _w7996_ ;
	wire _w7997_ ;
	wire _w7998_ ;
	wire _w7999_ ;
	wire _w8000_ ;
	wire _w8001_ ;
	wire _w8002_ ;
	wire _w8003_ ;
	wire _w8004_ ;
	wire _w8005_ ;
	wire _w8006_ ;
	wire _w8007_ ;
	wire _w8008_ ;
	wire _w8009_ ;
	wire _w8010_ ;
	wire _w8011_ ;
	wire _w8012_ ;
	wire _w8013_ ;
	wire _w8014_ ;
	wire _w8015_ ;
	wire _w8016_ ;
	wire _w8017_ ;
	wire _w8018_ ;
	wire _w8019_ ;
	wire _w8020_ ;
	wire _w8021_ ;
	wire _w8022_ ;
	wire _w8023_ ;
	wire _w8024_ ;
	wire _w8025_ ;
	wire _w8026_ ;
	wire _w8027_ ;
	wire _w8028_ ;
	wire _w8029_ ;
	wire _w8030_ ;
	wire _w8031_ ;
	wire _w8032_ ;
	wire _w8033_ ;
	wire _w8034_ ;
	wire _w8035_ ;
	wire _w8036_ ;
	wire _w8037_ ;
	wire _w8038_ ;
	wire _w8039_ ;
	wire _w8040_ ;
	wire _w8041_ ;
	wire _w8042_ ;
	wire _w8043_ ;
	wire _w8044_ ;
	wire _w8045_ ;
	wire _w8046_ ;
	wire _w8047_ ;
	wire _w8048_ ;
	wire _w8049_ ;
	wire _w8050_ ;
	wire _w8051_ ;
	wire _w8052_ ;
	wire _w8053_ ;
	wire _w8054_ ;
	wire _w8055_ ;
	wire _w8056_ ;
	wire _w8057_ ;
	wire _w8058_ ;
	wire _w8059_ ;
	wire _w8060_ ;
	wire _w8061_ ;
	wire _w8062_ ;
	wire _w8063_ ;
	wire _w8064_ ;
	wire _w8065_ ;
	wire _w8066_ ;
	wire _w8067_ ;
	wire _w8068_ ;
	wire _w8069_ ;
	wire _w8070_ ;
	wire _w8071_ ;
	wire _w8072_ ;
	wire _w8073_ ;
	wire _w8074_ ;
	wire _w8075_ ;
	wire _w8076_ ;
	wire _w8077_ ;
	wire _w8078_ ;
	wire _w8079_ ;
	wire _w8080_ ;
	wire _w8081_ ;
	wire _w8082_ ;
	wire _w8083_ ;
	wire _w8084_ ;
	wire _w8085_ ;
	wire _w8086_ ;
	wire _w8087_ ;
	wire _w8088_ ;
	wire _w8089_ ;
	wire _w8090_ ;
	wire _w8091_ ;
	wire _w8092_ ;
	wire _w8093_ ;
	wire _w8094_ ;
	wire _w8095_ ;
	wire _w8096_ ;
	wire _w8097_ ;
	wire _w8098_ ;
	wire _w8099_ ;
	wire _w8100_ ;
	wire _w8101_ ;
	wire _w8102_ ;
	wire _w8103_ ;
	wire _w8104_ ;
	wire _w8105_ ;
	wire _w8106_ ;
	wire _w8107_ ;
	wire _w8108_ ;
	wire _w8109_ ;
	wire _w8110_ ;
	wire _w8111_ ;
	wire _w8112_ ;
	wire _w8113_ ;
	wire _w8114_ ;
	wire _w8115_ ;
	wire _w8116_ ;
	wire _w8117_ ;
	wire _w8118_ ;
	wire _w8119_ ;
	wire _w8120_ ;
	wire _w8121_ ;
	wire _w8122_ ;
	wire _w8123_ ;
	wire _w8124_ ;
	wire _w8125_ ;
	wire _w8126_ ;
	wire _w8127_ ;
	wire _w8128_ ;
	wire _w8129_ ;
	wire _w8130_ ;
	wire _w8131_ ;
	wire _w8132_ ;
	wire _w8133_ ;
	wire _w8134_ ;
	wire _w8135_ ;
	wire _w8136_ ;
	wire _w8137_ ;
	wire _w8138_ ;
	wire _w8139_ ;
	wire _w8140_ ;
	wire _w8141_ ;
	wire _w8142_ ;
	wire _w8143_ ;
	wire _w8144_ ;
	wire _w8145_ ;
	wire _w8146_ ;
	wire _w8147_ ;
	wire _w8148_ ;
	wire _w8149_ ;
	wire _w8150_ ;
	wire _w8151_ ;
	wire _w8152_ ;
	wire _w8153_ ;
	wire _w8154_ ;
	wire _w8155_ ;
	wire _w8156_ ;
	wire _w8157_ ;
	wire _w8158_ ;
	wire _w8159_ ;
	wire _w8160_ ;
	wire _w8161_ ;
	wire _w8162_ ;
	wire _w8163_ ;
	wire _w8164_ ;
	wire _w8165_ ;
	wire _w8166_ ;
	wire _w8167_ ;
	wire _w8168_ ;
	wire _w8169_ ;
	wire _w8170_ ;
	wire _w8171_ ;
	wire _w8172_ ;
	wire _w8173_ ;
	wire _w8174_ ;
	wire _w8175_ ;
	wire _w8176_ ;
	wire _w8177_ ;
	wire _w8178_ ;
	wire _w8179_ ;
	wire _w8180_ ;
	wire _w8181_ ;
	wire _w8182_ ;
	wire _w8183_ ;
	wire _w8184_ ;
	wire _w8185_ ;
	wire _w8186_ ;
	wire _w8187_ ;
	wire _w8188_ ;
	wire _w8189_ ;
	wire _w8190_ ;
	wire _w8191_ ;
	wire _w8192_ ;
	wire _w8193_ ;
	wire _w8194_ ;
	wire _w8195_ ;
	wire _w8196_ ;
	wire _w8197_ ;
	wire _w8198_ ;
	wire _w8199_ ;
	wire _w8200_ ;
	wire _w8201_ ;
	wire _w8202_ ;
	wire _w8203_ ;
	wire _w8204_ ;
	wire _w8205_ ;
	wire _w8206_ ;
	wire _w8207_ ;
	wire _w8208_ ;
	wire _w8209_ ;
	wire _w8210_ ;
	wire _w8211_ ;
	wire _w8212_ ;
	wire _w8213_ ;
	wire _w8214_ ;
	wire _w8215_ ;
	wire _w8216_ ;
	wire _w8217_ ;
	wire _w8218_ ;
	wire _w8219_ ;
	wire _w8220_ ;
	wire _w8221_ ;
	wire _w8222_ ;
	wire _w8223_ ;
	wire _w8224_ ;
	wire _w8225_ ;
	wire _w8226_ ;
	wire _w8227_ ;
	wire _w8228_ ;
	wire _w8229_ ;
	wire _w8230_ ;
	wire _w8231_ ;
	wire _w8232_ ;
	wire _w8233_ ;
	wire _w8234_ ;
	wire _w8235_ ;
	wire _w8236_ ;
	wire _w8237_ ;
	wire _w8238_ ;
	wire _w8239_ ;
	wire _w8240_ ;
	wire _w8241_ ;
	wire _w8242_ ;
	wire _w8243_ ;
	wire _w8244_ ;
	wire _w8245_ ;
	wire _w8246_ ;
	wire _w8247_ ;
	wire _w8248_ ;
	wire _w8249_ ;
	wire _w8250_ ;
	wire _w8251_ ;
	wire _w8252_ ;
	wire _w8253_ ;
	wire _w8254_ ;
	wire _w8255_ ;
	wire _w8256_ ;
	wire _w8257_ ;
	wire _w8258_ ;
	wire _w8259_ ;
	wire _w8260_ ;
	wire _w8261_ ;
	wire _w8262_ ;
	wire _w8263_ ;
	wire _w8264_ ;
	wire _w8265_ ;
	wire _w8266_ ;
	wire _w8267_ ;
	wire _w8268_ ;
	wire _w8269_ ;
	wire _w8270_ ;
	wire _w8271_ ;
	wire _w8272_ ;
	wire _w8273_ ;
	wire _w8274_ ;
	wire _w8275_ ;
	wire _w8276_ ;
	wire _w8277_ ;
	wire _w8278_ ;
	wire _w8279_ ;
	wire _w8280_ ;
	wire _w8281_ ;
	wire _w8282_ ;
	wire _w8283_ ;
	wire _w8284_ ;
	wire _w8285_ ;
	wire _w8286_ ;
	wire _w8287_ ;
	wire _w8288_ ;
	wire _w8289_ ;
	wire _w8290_ ;
	wire _w8291_ ;
	wire _w8292_ ;
	wire _w8293_ ;
	wire _w8294_ ;
	wire _w8295_ ;
	wire _w8296_ ;
	wire _w8297_ ;
	wire _w8298_ ;
	wire _w8299_ ;
	wire _w8300_ ;
	wire _w8301_ ;
	wire _w8302_ ;
	wire _w8303_ ;
	wire _w8304_ ;
	wire _w8305_ ;
	wire _w8306_ ;
	wire _w8307_ ;
	wire _w8308_ ;
	wire _w8309_ ;
	wire _w8310_ ;
	wire _w8311_ ;
	wire _w8312_ ;
	wire _w8313_ ;
	wire _w8314_ ;
	wire _w8315_ ;
	wire _w8316_ ;
	wire _w8317_ ;
	wire _w8318_ ;
	wire _w8319_ ;
	wire _w8320_ ;
	wire _w8321_ ;
	wire _w8322_ ;
	wire _w8323_ ;
	wire _w8324_ ;
	wire _w8325_ ;
	wire _w8326_ ;
	wire _w8327_ ;
	wire _w8328_ ;
	wire _w8329_ ;
	wire _w8330_ ;
	wire _w8331_ ;
	wire _w8332_ ;
	wire _w8333_ ;
	wire _w8334_ ;
	wire _w8335_ ;
	wire _w8336_ ;
	wire _w8337_ ;
	wire _w8338_ ;
	wire _w8339_ ;
	wire _w8340_ ;
	wire _w8341_ ;
	wire _w8342_ ;
	wire _w8343_ ;
	wire _w8344_ ;
	wire _w8345_ ;
	wire _w8346_ ;
	wire _w8347_ ;
	wire _w8348_ ;
	wire _w8349_ ;
	wire _w8350_ ;
	wire _w8351_ ;
	wire _w8352_ ;
	wire _w8353_ ;
	wire _w8354_ ;
	wire _w8355_ ;
	wire _w8356_ ;
	wire _w8357_ ;
	wire _w8358_ ;
	wire _w8359_ ;
	wire _w8360_ ;
	wire _w8361_ ;
	wire _w8362_ ;
	wire _w8363_ ;
	wire _w8364_ ;
	wire _w8365_ ;
	wire _w8366_ ;
	wire _w8367_ ;
	wire _w8368_ ;
	wire _w8369_ ;
	wire _w8370_ ;
	wire _w8371_ ;
	wire _w8372_ ;
	wire _w8373_ ;
	wire _w8374_ ;
	wire _w8375_ ;
	wire _w8376_ ;
	wire _w8377_ ;
	wire _w8378_ ;
	wire _w8379_ ;
	wire _w8380_ ;
	wire _w8381_ ;
	wire _w8382_ ;
	wire _w8383_ ;
	wire _w8384_ ;
	wire _w8385_ ;
	wire _w8386_ ;
	wire _w8387_ ;
	wire _w8388_ ;
	wire _w8389_ ;
	wire _w8390_ ;
	wire _w8391_ ;
	wire _w8392_ ;
	wire _w8393_ ;
	wire _w8394_ ;
	wire _w8395_ ;
	wire _w8396_ ;
	wire _w8397_ ;
	wire _w8398_ ;
	wire _w8399_ ;
	wire _w8400_ ;
	wire _w8401_ ;
	wire _w8402_ ;
	wire _w8403_ ;
	wire _w8404_ ;
	wire _w8405_ ;
	wire _w8406_ ;
	wire _w8407_ ;
	wire _w8408_ ;
	wire _w8409_ ;
	wire _w8410_ ;
	wire _w8411_ ;
	wire _w8412_ ;
	wire _w8413_ ;
	wire _w8414_ ;
	wire _w8415_ ;
	wire _w8416_ ;
	wire _w8417_ ;
	wire _w8418_ ;
	wire _w8419_ ;
	wire _w8420_ ;
	wire _w8421_ ;
	wire _w8422_ ;
	wire _w8423_ ;
	wire _w8424_ ;
	wire _w8425_ ;
	wire _w8426_ ;
	wire _w8427_ ;
	wire _w8428_ ;
	wire _w8429_ ;
	wire _w8430_ ;
	wire _w8431_ ;
	wire _w8432_ ;
	wire _w8433_ ;
	wire _w8434_ ;
	wire _w8435_ ;
	wire _w8436_ ;
	wire _w8437_ ;
	wire _w8438_ ;
	wire _w8439_ ;
	wire _w8440_ ;
	wire _w8441_ ;
	wire _w8442_ ;
	wire _w8443_ ;
	wire _w8444_ ;
	wire _w8445_ ;
	wire _w8446_ ;
	wire _w8447_ ;
	wire _w8448_ ;
	wire _w8449_ ;
	wire _w8450_ ;
	wire _w8451_ ;
	wire _w8452_ ;
	wire _w8453_ ;
	wire _w8454_ ;
	wire _w8455_ ;
	wire _w8456_ ;
	wire _w8457_ ;
	wire _w8458_ ;
	wire _w8459_ ;
	wire _w8460_ ;
	wire _w8461_ ;
	wire _w8462_ ;
	wire _w8463_ ;
	wire _w8464_ ;
	wire _w8465_ ;
	wire _w8466_ ;
	wire _w8467_ ;
	wire _w8468_ ;
	wire _w8469_ ;
	wire _w8470_ ;
	wire _w8471_ ;
	wire _w8472_ ;
	wire _w8473_ ;
	wire _w8474_ ;
	wire _w8475_ ;
	wire _w8476_ ;
	wire _w8477_ ;
	wire _w8478_ ;
	wire _w8479_ ;
	wire _w8480_ ;
	wire _w8481_ ;
	wire _w8482_ ;
	wire _w8483_ ;
	wire _w8484_ ;
	wire _w8485_ ;
	wire _w8486_ ;
	wire _w8487_ ;
	wire _w8488_ ;
	wire _w8489_ ;
	wire _w8490_ ;
	wire _w8491_ ;
	wire _w8492_ ;
	wire _w8493_ ;
	wire _w8494_ ;
	wire _w8495_ ;
	wire _w8496_ ;
	wire _w8497_ ;
	wire _w8498_ ;
	wire _w8499_ ;
	wire _w8500_ ;
	wire _w8501_ ;
	wire _w8502_ ;
	wire _w8503_ ;
	wire _w8504_ ;
	wire _w8505_ ;
	wire _w8506_ ;
	wire _w8507_ ;
	wire _w8508_ ;
	wire _w8509_ ;
	wire _w8510_ ;
	wire _w8511_ ;
	wire _w8512_ ;
	wire _w8513_ ;
	wire _w8514_ ;
	wire _w8515_ ;
	wire _w8516_ ;
	wire _w8517_ ;
	wire _w8518_ ;
	wire _w8519_ ;
	wire _w8520_ ;
	wire _w8521_ ;
	wire _w8522_ ;
	wire _w8523_ ;
	wire _w8524_ ;
	wire _w8525_ ;
	wire _w8526_ ;
	wire _w8527_ ;
	wire _w8528_ ;
	wire _w8529_ ;
	wire _w8530_ ;
	wire _w8531_ ;
	wire _w8532_ ;
	wire _w8533_ ;
	wire _w8534_ ;
	wire _w8535_ ;
	wire _w8536_ ;
	wire _w8537_ ;
	wire _w8538_ ;
	wire _w8539_ ;
	wire _w8540_ ;
	wire _w8541_ ;
	wire _w8542_ ;
	wire _w8543_ ;
	wire _w8544_ ;
	wire _w8545_ ;
	wire _w8546_ ;
	wire _w8547_ ;
	wire _w8548_ ;
	wire _w8549_ ;
	wire _w8550_ ;
	wire _w8551_ ;
	wire _w8552_ ;
	wire _w8553_ ;
	wire _w8554_ ;
	wire _w8555_ ;
	wire _w8556_ ;
	wire _w8557_ ;
	wire _w8558_ ;
	wire _w8559_ ;
	wire _w8560_ ;
	wire _w8561_ ;
	wire _w8562_ ;
	wire _w8563_ ;
	wire _w8564_ ;
	wire _w8565_ ;
	wire _w8566_ ;
	wire _w8567_ ;
	wire _w8568_ ;
	wire _w8569_ ;
	wire _w8570_ ;
	wire _w8571_ ;
	wire _w8572_ ;
	wire _w8573_ ;
	wire _w8574_ ;
	wire _w8575_ ;
	wire _w8576_ ;
	wire _w8577_ ;
	wire _w8578_ ;
	wire _w8579_ ;
	wire _w8580_ ;
	wire _w8581_ ;
	wire _w8582_ ;
	wire _w8583_ ;
	wire _w8584_ ;
	wire _w8585_ ;
	wire _w8586_ ;
	wire _w8587_ ;
	wire _w8588_ ;
	wire _w8589_ ;
	wire _w8590_ ;
	wire _w8591_ ;
	wire _w8592_ ;
	wire _w8593_ ;
	wire _w8594_ ;
	wire _w8595_ ;
	wire _w8596_ ;
	wire _w8597_ ;
	wire _w8598_ ;
	wire _w8599_ ;
	wire _w8600_ ;
	wire _w8601_ ;
	wire _w8602_ ;
	wire _w8603_ ;
	wire _w8604_ ;
	wire _w8605_ ;
	wire _w8606_ ;
	wire _w8607_ ;
	wire _w8608_ ;
	wire _w8609_ ;
	wire _w8610_ ;
	wire _w8611_ ;
	wire _w8612_ ;
	wire _w8613_ ;
	wire _w8614_ ;
	wire _w8615_ ;
	wire _w8616_ ;
	wire _w8617_ ;
	wire _w8618_ ;
	wire _w8619_ ;
	wire _w8620_ ;
	wire _w8621_ ;
	wire _w8622_ ;
	wire _w8623_ ;
	wire _w8624_ ;
	wire _w8625_ ;
	wire _w8626_ ;
	wire _w8627_ ;
	wire _w8628_ ;
	wire _w8629_ ;
	wire _w8630_ ;
	wire _w8631_ ;
	wire _w8632_ ;
	wire _w8633_ ;
	wire _w8634_ ;
	wire _w8635_ ;
	wire _w8636_ ;
	wire _w8637_ ;
	wire _w8638_ ;
	wire _w8639_ ;
	wire _w8640_ ;
	wire _w8641_ ;
	wire _w8642_ ;
	wire _w8643_ ;
	wire _w8644_ ;
	wire _w8645_ ;
	wire _w8646_ ;
	wire _w8647_ ;
	wire _w8648_ ;
	wire _w8649_ ;
	wire _w8650_ ;
	wire _w8651_ ;
	wire _w8652_ ;
	wire _w8653_ ;
	wire _w8654_ ;
	wire _w8655_ ;
	wire _w8656_ ;
	wire _w8657_ ;
	wire _w8658_ ;
	wire _w8659_ ;
	wire _w8660_ ;
	wire _w8661_ ;
	wire _w8662_ ;
	wire _w8663_ ;
	wire _w8664_ ;
	wire _w8665_ ;
	wire _w8666_ ;
	wire _w8667_ ;
	wire _w8668_ ;
	wire _w8669_ ;
	wire _w8670_ ;
	wire _w8671_ ;
	wire _w8672_ ;
	wire _w8673_ ;
	wire _w8674_ ;
	wire _w8675_ ;
	wire _w8676_ ;
	wire _w8677_ ;
	wire _w8678_ ;
	wire _w8679_ ;
	wire _w8680_ ;
	wire _w8681_ ;
	wire _w8682_ ;
	wire _w8683_ ;
	wire _w8684_ ;
	wire _w8685_ ;
	wire _w8686_ ;
	wire _w8687_ ;
	wire _w8688_ ;
	wire _w8689_ ;
	wire _w8690_ ;
	wire _w8691_ ;
	wire _w8692_ ;
	wire _w8693_ ;
	wire _w8694_ ;
	wire _w8695_ ;
	wire _w8696_ ;
	wire _w8697_ ;
	wire _w8698_ ;
	wire _w8699_ ;
	wire _w8700_ ;
	wire _w8701_ ;
	wire _w8702_ ;
	wire _w8703_ ;
	wire _w8704_ ;
	wire _w8705_ ;
	wire _w8706_ ;
	wire _w8707_ ;
	wire _w8708_ ;
	wire _w8709_ ;
	wire _w8710_ ;
	wire _w8711_ ;
	wire _w8712_ ;
	wire _w8713_ ;
	wire _w8714_ ;
	wire _w8715_ ;
	wire _w8716_ ;
	wire _w8717_ ;
	wire _w8718_ ;
	wire _w8719_ ;
	wire _w8720_ ;
	wire _w8721_ ;
	wire _w8722_ ;
	wire _w8723_ ;
	wire _w8724_ ;
	wire _w8725_ ;
	wire _w8726_ ;
	wire _w8727_ ;
	wire _w8728_ ;
	wire _w8729_ ;
	wire _w8730_ ;
	wire _w8731_ ;
	wire _w8732_ ;
	wire _w8733_ ;
	wire _w8734_ ;
	wire _w8735_ ;
	wire _w8736_ ;
	wire _w8737_ ;
	wire _w8738_ ;
	wire _w8739_ ;
	wire _w8740_ ;
	wire _w8741_ ;
	wire _w8742_ ;
	wire _w8743_ ;
	wire _w8744_ ;
	wire _w8745_ ;
	wire _w8746_ ;
	wire _w8747_ ;
	wire _w8748_ ;
	wire _w8749_ ;
	wire _w8750_ ;
	wire _w8751_ ;
	wire _w8752_ ;
	wire _w8753_ ;
	wire _w8754_ ;
	wire _w8755_ ;
	wire _w8756_ ;
	wire _w8757_ ;
	wire _w8758_ ;
	wire _w8759_ ;
	wire _w8760_ ;
	wire _w8761_ ;
	wire _w8762_ ;
	wire _w8763_ ;
	wire _w8764_ ;
	wire _w8765_ ;
	wire _w8766_ ;
	wire _w8767_ ;
	wire _w8768_ ;
	wire _w8769_ ;
	wire _w8770_ ;
	wire _w8771_ ;
	wire _w8772_ ;
	wire _w8773_ ;
	wire _w8774_ ;
	wire _w8775_ ;
	wire _w8776_ ;
	wire _w8777_ ;
	wire _w8778_ ;
	wire _w8779_ ;
	wire _w8780_ ;
	wire _w8781_ ;
	wire _w8782_ ;
	wire _w8783_ ;
	wire _w8784_ ;
	wire _w8785_ ;
	wire _w8786_ ;
	wire _w8787_ ;
	wire _w8788_ ;
	wire _w8789_ ;
	wire _w8790_ ;
	wire _w8791_ ;
	wire _w8792_ ;
	wire _w8793_ ;
	wire _w8794_ ;
	wire _w8795_ ;
	wire _w8796_ ;
	wire _w8797_ ;
	wire _w8798_ ;
	wire _w8799_ ;
	wire _w8800_ ;
	wire _w8801_ ;
	wire _w8802_ ;
	wire _w8803_ ;
	wire _w8804_ ;
	wire _w8805_ ;
	wire _w8806_ ;
	wire _w8807_ ;
	wire _w8808_ ;
	wire _w8809_ ;
	wire _w8810_ ;
	wire _w8811_ ;
	wire _w8812_ ;
	wire _w8813_ ;
	wire _w8814_ ;
	wire _w8815_ ;
	wire _w8816_ ;
	wire _w8817_ ;
	wire _w8818_ ;
	wire _w8819_ ;
	wire _w8820_ ;
	wire _w8821_ ;
	wire _w8822_ ;
	wire _w8823_ ;
	wire _w8824_ ;
	wire _w8825_ ;
	wire _w8826_ ;
	wire _w8827_ ;
	wire _w8828_ ;
	wire _w8829_ ;
	wire _w8830_ ;
	wire _w8831_ ;
	wire _w8832_ ;
	wire _w8833_ ;
	wire _w8834_ ;
	wire _w8835_ ;
	wire _w8836_ ;
	wire _w8837_ ;
	wire _w8838_ ;
	wire _w8839_ ;
	wire _w8840_ ;
	wire _w8841_ ;
	wire _w8842_ ;
	wire _w8843_ ;
	wire _w8844_ ;
	wire _w8845_ ;
	wire _w8846_ ;
	wire _w8847_ ;
	wire _w8848_ ;
	wire _w8849_ ;
	wire _w8850_ ;
	wire _w8851_ ;
	wire _w8852_ ;
	wire _w8853_ ;
	wire _w8854_ ;
	wire _w8855_ ;
	wire _w8856_ ;
	wire _w8857_ ;
	wire _w8858_ ;
	wire _w8859_ ;
	wire _w8860_ ;
	wire _w8861_ ;
	wire _w8862_ ;
	wire _w8863_ ;
	wire _w8864_ ;
	wire _w8865_ ;
	wire _w8866_ ;
	wire _w8867_ ;
	wire _w8868_ ;
	wire _w8869_ ;
	wire _w8870_ ;
	wire _w8871_ ;
	wire _w8872_ ;
	wire _w8873_ ;
	wire _w8874_ ;
	wire _w8875_ ;
	wire _w8876_ ;
	wire _w8877_ ;
	wire _w8878_ ;
	wire _w8879_ ;
	wire _w8880_ ;
	wire _w8881_ ;
	wire _w8882_ ;
	wire _w8883_ ;
	wire _w8884_ ;
	wire _w8885_ ;
	wire _w8886_ ;
	wire _w8887_ ;
	wire _w8888_ ;
	wire _w8889_ ;
	wire _w8890_ ;
	wire _w8891_ ;
	wire _w8892_ ;
	wire _w8893_ ;
	wire _w8894_ ;
	wire _w8895_ ;
	wire _w8896_ ;
	wire _w8897_ ;
	wire _w8898_ ;
	wire _w8899_ ;
	wire _w8900_ ;
	wire _w8901_ ;
	wire _w8902_ ;
	wire _w8903_ ;
	wire _w8904_ ;
	wire _w8905_ ;
	wire _w8906_ ;
	wire _w8907_ ;
	wire _w8908_ ;
	wire _w8909_ ;
	wire _w8910_ ;
	wire _w8911_ ;
	wire _w8912_ ;
	wire _w8913_ ;
	wire _w8914_ ;
	wire _w8915_ ;
	wire _w8916_ ;
	wire _w8917_ ;
	wire _w8918_ ;
	wire _w8919_ ;
	wire _w8920_ ;
	wire _w8921_ ;
	wire _w8922_ ;
	wire _w8923_ ;
	wire _w8924_ ;
	wire _w8925_ ;
	wire _w8926_ ;
	wire _w8927_ ;
	wire _w8928_ ;
	wire _w8929_ ;
	wire _w8930_ ;
	wire _w8931_ ;
	wire _w8932_ ;
	wire _w8933_ ;
	wire _w8934_ ;
	wire _w8935_ ;
	wire _w8936_ ;
	wire _w8937_ ;
	wire _w8938_ ;
	wire _w8939_ ;
	wire _w8940_ ;
	wire _w8941_ ;
	wire _w8942_ ;
	wire _w8943_ ;
	wire _w8944_ ;
	wire _w8945_ ;
	wire _w8946_ ;
	wire _w8947_ ;
	wire _w8948_ ;
	wire _w8949_ ;
	wire _w8950_ ;
	wire _w8951_ ;
	wire _w8952_ ;
	wire _w8953_ ;
	wire _w8954_ ;
	wire _w8955_ ;
	wire _w8956_ ;
	wire _w8957_ ;
	wire _w8958_ ;
	wire _w8959_ ;
	wire _w8960_ ;
	wire _w8961_ ;
	wire _w8962_ ;
	wire _w8963_ ;
	wire _w8964_ ;
	wire _w8965_ ;
	wire _w8966_ ;
	wire _w8967_ ;
	wire _w8968_ ;
	wire _w8969_ ;
	wire _w8970_ ;
	wire _w8971_ ;
	wire _w8972_ ;
	wire _w8973_ ;
	wire _w8974_ ;
	wire _w8975_ ;
	wire _w8976_ ;
	wire _w8977_ ;
	wire _w8978_ ;
	wire _w8979_ ;
	wire _w8980_ ;
	wire _w8981_ ;
	wire _w8982_ ;
	wire _w8983_ ;
	wire _w8984_ ;
	wire _w8985_ ;
	wire _w8986_ ;
	wire _w8987_ ;
	wire _w8988_ ;
	wire _w8989_ ;
	wire _w8990_ ;
	wire _w8991_ ;
	wire _w8992_ ;
	wire _w8993_ ;
	wire _w8994_ ;
	wire _w8995_ ;
	wire _w8996_ ;
	wire _w8997_ ;
	wire _w8998_ ;
	wire _w8999_ ;
	wire _w9000_ ;
	wire _w9001_ ;
	wire _w9002_ ;
	wire _w9003_ ;
	wire _w9004_ ;
	wire _w9005_ ;
	wire _w9006_ ;
	wire _w9007_ ;
	wire _w9008_ ;
	wire _w9009_ ;
	wire _w9010_ ;
	wire _w9011_ ;
	wire _w9012_ ;
	wire _w9013_ ;
	wire _w9014_ ;
	wire _w9015_ ;
	wire _w9016_ ;
	wire _w9017_ ;
	wire _w9018_ ;
	wire _w9019_ ;
	wire _w9020_ ;
	wire _w9021_ ;
	wire _w9022_ ;
	wire _w9023_ ;
	wire _w9024_ ;
	wire _w9025_ ;
	wire _w9026_ ;
	wire _w9027_ ;
	wire _w9028_ ;
	wire _w9029_ ;
	wire _w9030_ ;
	wire _w9031_ ;
	wire _w9032_ ;
	wire _w9033_ ;
	wire _w9034_ ;
	wire _w9035_ ;
	wire _w9036_ ;
	wire _w9037_ ;
	wire _w9038_ ;
	wire _w9039_ ;
	wire _w9040_ ;
	wire _w9041_ ;
	wire _w9042_ ;
	wire _w9043_ ;
	wire _w9044_ ;
	wire _w9045_ ;
	wire _w9046_ ;
	wire _w9047_ ;
	wire _w9048_ ;
	wire _w9049_ ;
	wire _w9050_ ;
	wire _w9051_ ;
	wire _w9052_ ;
	wire _w9053_ ;
	wire _w9054_ ;
	wire _w9055_ ;
	wire _w9056_ ;
	wire _w9057_ ;
	wire _w9058_ ;
	wire _w9059_ ;
	wire _w9060_ ;
	wire _w9061_ ;
	wire _w9062_ ;
	wire _w9063_ ;
	wire _w9064_ ;
	wire _w9065_ ;
	wire _w9066_ ;
	wire _w9067_ ;
	wire _w9068_ ;
	wire _w9069_ ;
	wire _w9070_ ;
	wire _w9071_ ;
	wire _w9072_ ;
	wire _w9073_ ;
	wire _w9074_ ;
	wire _w9075_ ;
	wire _w9076_ ;
	wire _w9077_ ;
	wire _w9078_ ;
	wire _w9079_ ;
	wire _w9080_ ;
	wire _w9081_ ;
	wire _w9082_ ;
	wire _w9083_ ;
	wire _w9084_ ;
	wire _w9085_ ;
	wire _w9086_ ;
	wire _w9087_ ;
	wire _w9088_ ;
	wire _w9089_ ;
	wire _w9090_ ;
	wire _w9091_ ;
	wire _w9092_ ;
	wire _w9093_ ;
	wire _w9094_ ;
	wire _w9095_ ;
	wire _w9096_ ;
	wire _w9097_ ;
	wire _w9098_ ;
	wire _w9099_ ;
	wire _w9100_ ;
	wire _w9101_ ;
	wire _w9102_ ;
	wire _w9103_ ;
	wire _w9104_ ;
	wire _w9105_ ;
	wire _w9106_ ;
	wire _w9107_ ;
	wire _w9108_ ;
	wire _w9109_ ;
	wire _w9110_ ;
	wire _w9111_ ;
	wire _w9112_ ;
	wire _w9113_ ;
	wire _w9114_ ;
	wire _w9115_ ;
	wire _w9116_ ;
	wire _w9117_ ;
	wire _w9118_ ;
	wire _w9119_ ;
	wire _w9120_ ;
	wire _w9121_ ;
	wire _w9122_ ;
	wire _w9123_ ;
	wire _w9124_ ;
	wire _w9125_ ;
	wire _w9126_ ;
	wire _w9127_ ;
	wire _w9128_ ;
	wire _w9129_ ;
	wire _w9130_ ;
	wire _w9131_ ;
	wire _w9132_ ;
	wire _w9133_ ;
	wire _w9134_ ;
	wire _w9135_ ;
	wire _w9136_ ;
	wire _w9137_ ;
	wire _w9138_ ;
	wire _w9139_ ;
	wire _w9140_ ;
	wire _w9141_ ;
	wire _w9142_ ;
	wire _w9143_ ;
	wire _w9144_ ;
	wire _w9145_ ;
	wire _w9146_ ;
	wire _w9147_ ;
	wire _w9148_ ;
	wire _w9149_ ;
	wire _w9150_ ;
	wire _w9151_ ;
	wire _w9152_ ;
	wire _w9153_ ;
	wire _w9154_ ;
	wire _w9155_ ;
	wire _w9156_ ;
	wire _w9157_ ;
	wire _w9158_ ;
	wire _w9159_ ;
	wire _w9160_ ;
	wire _w9161_ ;
	wire _w9162_ ;
	wire _w9163_ ;
	wire _w9164_ ;
	wire _w9165_ ;
	wire _w9166_ ;
	wire _w9167_ ;
	wire _w9168_ ;
	wire _w9169_ ;
	wire _w9170_ ;
	wire _w9171_ ;
	wire _w9172_ ;
	wire _w9173_ ;
	wire _w9174_ ;
	wire _w9175_ ;
	wire _w9176_ ;
	wire _w9177_ ;
	wire _w9178_ ;
	wire _w9179_ ;
	wire _w9180_ ;
	wire _w9181_ ;
	wire _w9182_ ;
	wire _w9183_ ;
	wire _w9184_ ;
	wire _w9185_ ;
	wire _w9186_ ;
	wire _w9187_ ;
	wire _w9188_ ;
	wire _w9189_ ;
	wire _w9190_ ;
	wire _w9191_ ;
	wire _w9192_ ;
	wire _w9193_ ;
	wire _w9194_ ;
	wire _w9195_ ;
	wire _w9196_ ;
	wire _w9197_ ;
	wire _w9198_ ;
	wire _w9199_ ;
	wire _w9200_ ;
	wire _w9201_ ;
	wire _w9202_ ;
	wire _w9203_ ;
	wire _w9204_ ;
	wire _w9205_ ;
	wire _w9206_ ;
	wire _w9207_ ;
	wire _w9208_ ;
	wire _w9209_ ;
	wire _w9210_ ;
	wire _w9211_ ;
	wire _w9212_ ;
	wire _w9213_ ;
	wire _w9214_ ;
	wire _w9215_ ;
	wire _w9216_ ;
	wire _w9217_ ;
	wire _w9218_ ;
	wire _w9219_ ;
	wire _w9220_ ;
	wire _w9221_ ;
	wire _w9222_ ;
	wire _w9223_ ;
	wire _w9224_ ;
	wire _w9225_ ;
	wire _w9226_ ;
	wire _w9227_ ;
	wire _w9228_ ;
	wire _w9229_ ;
	wire _w9230_ ;
	wire _w9231_ ;
	wire _w9232_ ;
	wire _w9233_ ;
	wire _w9234_ ;
	wire _w9235_ ;
	wire _w9236_ ;
	wire _w9237_ ;
	wire _w9238_ ;
	wire _w9239_ ;
	wire _w9240_ ;
	wire _w9241_ ;
	wire _w9242_ ;
	wire _w9243_ ;
	wire _w9244_ ;
	wire _w9245_ ;
	wire _w9246_ ;
	wire _w9247_ ;
	wire _w9248_ ;
	wire _w9249_ ;
	wire _w9250_ ;
	wire _w9251_ ;
	wire _w9252_ ;
	wire _w9253_ ;
	wire _w9254_ ;
	wire _w9255_ ;
	wire _w9256_ ;
	wire _w9257_ ;
	wire _w9258_ ;
	wire _w9259_ ;
	wire _w9260_ ;
	wire _w9261_ ;
	wire _w9262_ ;
	wire _w9263_ ;
	wire _w9264_ ;
	wire _w9265_ ;
	wire _w9266_ ;
	wire _w9267_ ;
	wire _w9268_ ;
	wire _w9269_ ;
	wire _w9270_ ;
	wire _w9271_ ;
	wire _w9272_ ;
	wire _w9273_ ;
	wire _w9274_ ;
	wire _w9275_ ;
	wire _w9276_ ;
	wire _w9277_ ;
	wire _w9278_ ;
	wire _w9279_ ;
	wire _w9280_ ;
	wire _w9281_ ;
	wire _w9282_ ;
	wire _w9283_ ;
	wire _w9284_ ;
	wire _w9285_ ;
	wire _w9286_ ;
	wire _w9287_ ;
	wire _w9288_ ;
	wire _w9289_ ;
	wire _w9290_ ;
	wire _w9291_ ;
	wire _w9292_ ;
	wire _w9293_ ;
	wire _w9294_ ;
	wire _w9295_ ;
	wire _w9296_ ;
	wire _w9297_ ;
	wire _w9298_ ;
	wire _w9299_ ;
	wire _w9300_ ;
	wire _w9301_ ;
	wire _w9302_ ;
	wire _w9303_ ;
	wire _w9304_ ;
	wire _w9305_ ;
	wire _w9306_ ;
	wire _w9307_ ;
	wire _w9308_ ;
	wire _w9309_ ;
	wire _w9310_ ;
	wire _w9311_ ;
	wire _w9312_ ;
	wire _w9313_ ;
	wire _w9314_ ;
	wire _w9315_ ;
	wire _w9316_ ;
	wire _w9317_ ;
	wire _w9318_ ;
	wire _w9319_ ;
	wire _w9320_ ;
	wire _w9321_ ;
	wire _w9322_ ;
	wire _w9323_ ;
	wire _w9324_ ;
	wire _w9325_ ;
	wire _w9326_ ;
	wire _w9327_ ;
	wire _w9328_ ;
	wire _w9329_ ;
	wire _w9330_ ;
	wire _w9331_ ;
	wire _w9332_ ;
	wire _w9333_ ;
	wire _w9334_ ;
	wire _w9335_ ;
	wire _w9336_ ;
	wire _w9337_ ;
	wire _w9338_ ;
	wire _w9339_ ;
	wire _w9340_ ;
	wire _w9341_ ;
	wire _w9342_ ;
	wire _w9343_ ;
	wire _w9344_ ;
	wire _w9345_ ;
	wire _w9346_ ;
	wire _w9347_ ;
	wire _w9348_ ;
	wire _w9349_ ;
	wire _w9350_ ;
	wire _w9351_ ;
	wire _w9352_ ;
	wire _w9353_ ;
	wire _w9354_ ;
	wire _w9355_ ;
	wire _w9356_ ;
	wire _w9357_ ;
	wire _w9358_ ;
	wire _w9359_ ;
	wire _w9360_ ;
	wire _w9361_ ;
	wire _w9362_ ;
	wire _w9363_ ;
	wire _w9364_ ;
	wire _w9365_ ;
	wire _w9366_ ;
	wire _w9367_ ;
	wire _w9368_ ;
	wire _w9369_ ;
	wire _w9370_ ;
	wire _w9371_ ;
	wire _w9372_ ;
	wire _w9373_ ;
	wire _w9374_ ;
	wire _w9375_ ;
	wire _w9376_ ;
	wire _w9377_ ;
	wire _w9378_ ;
	wire _w9379_ ;
	wire _w9380_ ;
	wire _w9381_ ;
	wire _w9382_ ;
	wire _w9383_ ;
	wire _w9384_ ;
	wire _w9385_ ;
	wire _w9386_ ;
	wire _w9387_ ;
	wire _w9388_ ;
	wire _w9389_ ;
	wire _w9390_ ;
	wire _w9391_ ;
	wire _w9392_ ;
	wire _w9393_ ;
	wire _w9394_ ;
	wire _w9395_ ;
	wire _w9396_ ;
	wire _w9397_ ;
	wire _w9398_ ;
	wire _w9399_ ;
	wire _w9400_ ;
	wire _w9401_ ;
	wire _w9402_ ;
	wire _w9403_ ;
	wire _w9404_ ;
	wire _w9405_ ;
	wire _w9406_ ;
	wire _w9407_ ;
	wire _w9408_ ;
	wire _w9409_ ;
	wire _w9410_ ;
	wire _w9411_ ;
	wire _w9412_ ;
	wire _w9413_ ;
	wire _w9414_ ;
	wire _w9415_ ;
	wire _w9416_ ;
	wire _w9417_ ;
	wire _w9418_ ;
	wire _w9419_ ;
	wire _w9420_ ;
	wire _w9421_ ;
	wire _w9422_ ;
	wire _w9423_ ;
	wire _w9424_ ;
	wire _w9425_ ;
	wire _w9426_ ;
	wire _w9427_ ;
	wire _w9428_ ;
	wire _w9429_ ;
	wire _w9430_ ;
	wire _w9431_ ;
	wire _w9432_ ;
	wire _w9433_ ;
	wire _w9434_ ;
	wire _w9435_ ;
	wire _w9436_ ;
	wire _w9437_ ;
	wire _w9438_ ;
	wire _w9439_ ;
	wire _w9440_ ;
	wire _w9441_ ;
	wire _w9442_ ;
	wire _w9443_ ;
	wire _w9444_ ;
	wire _w9445_ ;
	wire _w9446_ ;
	wire _w9447_ ;
	wire _w9448_ ;
	wire _w9449_ ;
	wire _w9450_ ;
	wire _w9451_ ;
	wire _w9452_ ;
	wire _w9453_ ;
	wire _w9454_ ;
	wire _w9455_ ;
	wire _w9456_ ;
	wire _w9457_ ;
	wire _w9458_ ;
	wire _w9459_ ;
	wire _w9460_ ;
	wire _w9461_ ;
	wire _w9462_ ;
	wire _w9463_ ;
	wire _w9464_ ;
	wire _w9465_ ;
	wire _w9466_ ;
	wire _w9467_ ;
	wire _w9468_ ;
	wire _w9469_ ;
	wire _w9470_ ;
	wire _w9471_ ;
	wire _w9472_ ;
	wire _w9473_ ;
	wire _w9474_ ;
	wire _w9475_ ;
	wire _w9476_ ;
	wire _w9477_ ;
	wire _w9478_ ;
	wire _w9479_ ;
	wire _w9480_ ;
	wire _w9481_ ;
	wire _w9482_ ;
	wire _w9483_ ;
	wire _w9484_ ;
	wire _w9485_ ;
	wire _w9486_ ;
	wire _w9487_ ;
	wire _w9488_ ;
	wire _w9489_ ;
	wire _w9490_ ;
	wire _w9491_ ;
	wire _w9492_ ;
	wire _w9493_ ;
	wire _w9494_ ;
	wire _w9495_ ;
	wire _w9496_ ;
	wire _w9497_ ;
	wire _w9498_ ;
	wire _w9499_ ;
	wire _w9500_ ;
	wire _w9501_ ;
	wire _w9502_ ;
	wire _w9503_ ;
	wire _w9504_ ;
	wire _w9505_ ;
	wire _w9506_ ;
	wire _w9507_ ;
	wire _w9508_ ;
	wire _w9509_ ;
	wire _w9510_ ;
	wire _w9511_ ;
	wire _w9512_ ;
	wire _w9513_ ;
	wire _w9514_ ;
	wire _w9515_ ;
	wire _w9516_ ;
	wire _w9517_ ;
	wire _w9518_ ;
	wire _w9519_ ;
	wire _w9520_ ;
	wire _w9521_ ;
	wire _w9522_ ;
	wire _w9523_ ;
	wire _w9524_ ;
	wire _w9525_ ;
	wire _w9526_ ;
	wire _w9527_ ;
	wire _w9528_ ;
	wire _w9529_ ;
	wire _w9530_ ;
	wire _w9531_ ;
	wire _w9532_ ;
	wire _w9533_ ;
	wire _w9534_ ;
	wire _w9535_ ;
	wire _w9536_ ;
	wire _w9537_ ;
	wire _w9538_ ;
	wire _w9539_ ;
	wire _w9540_ ;
	wire _w9541_ ;
	wire _w9542_ ;
	wire _w9543_ ;
	wire _w9544_ ;
	wire _w9545_ ;
	wire _w9546_ ;
	wire _w9547_ ;
	wire _w9548_ ;
	wire _w9549_ ;
	wire _w9550_ ;
	wire _w9551_ ;
	wire _w9552_ ;
	wire _w9553_ ;
	wire _w9554_ ;
	wire _w9555_ ;
	wire _w9556_ ;
	wire _w9557_ ;
	wire _w9558_ ;
	wire _w9559_ ;
	wire _w9560_ ;
	wire _w9561_ ;
	wire _w9562_ ;
	wire _w9563_ ;
	wire _w9564_ ;
	wire _w9565_ ;
	wire _w9566_ ;
	wire _w9567_ ;
	wire _w9568_ ;
	wire _w9569_ ;
	wire _w9570_ ;
	wire _w9571_ ;
	wire _w9572_ ;
	wire _w9573_ ;
	wire _w9574_ ;
	wire _w9575_ ;
	wire _w9576_ ;
	wire _w9577_ ;
	wire _w9578_ ;
	wire _w9579_ ;
	wire _w9580_ ;
	wire _w9581_ ;
	wire _w9582_ ;
	wire _w9583_ ;
	wire _w9584_ ;
	wire _w9585_ ;
	wire _w9586_ ;
	wire _w9587_ ;
	wire _w9588_ ;
	wire _w9589_ ;
	wire _w9590_ ;
	wire _w9591_ ;
	wire _w9592_ ;
	wire _w9593_ ;
	wire _w9594_ ;
	wire _w9595_ ;
	wire _w9596_ ;
	wire _w9597_ ;
	wire _w9598_ ;
	wire _w9599_ ;
	wire _w9600_ ;
	wire _w9601_ ;
	wire _w9602_ ;
	wire _w9603_ ;
	wire _w9604_ ;
	wire _w9605_ ;
	wire _w9606_ ;
	wire _w9607_ ;
	wire _w9608_ ;
	wire _w9609_ ;
	wire _w9610_ ;
	wire _w9611_ ;
	wire _w9612_ ;
	wire _w9613_ ;
	wire _w9614_ ;
	wire _w9615_ ;
	wire _w9616_ ;
	wire _w9617_ ;
	wire _w9618_ ;
	wire _w9619_ ;
	wire _w9620_ ;
	wire _w9621_ ;
	wire _w9622_ ;
	wire _w9623_ ;
	wire _w9624_ ;
	wire _w9625_ ;
	wire _w9626_ ;
	wire _w9627_ ;
	wire _w9628_ ;
	wire _w9629_ ;
	wire _w9630_ ;
	wire _w9631_ ;
	wire _w9632_ ;
	wire _w9633_ ;
	wire _w9634_ ;
	wire _w9635_ ;
	wire _w9636_ ;
	wire _w9637_ ;
	wire _w9638_ ;
	wire _w9639_ ;
	wire _w9640_ ;
	wire _w9641_ ;
	wire _w9642_ ;
	wire _w9643_ ;
	wire _w9644_ ;
	wire _w9645_ ;
	wire _w9646_ ;
	wire _w9647_ ;
	wire _w9648_ ;
	wire _w9649_ ;
	wire _w9650_ ;
	wire _w9651_ ;
	wire _w9652_ ;
	wire _w9653_ ;
	wire _w9654_ ;
	wire _w9655_ ;
	wire _w9656_ ;
	wire _w9657_ ;
	wire _w9658_ ;
	wire _w9659_ ;
	wire _w9660_ ;
	wire _w9661_ ;
	wire _w9662_ ;
	wire _w9663_ ;
	wire _w9664_ ;
	wire _w9665_ ;
	wire _w9666_ ;
	wire _w9667_ ;
	wire _w9668_ ;
	wire _w9669_ ;
	wire _w9670_ ;
	wire _w9671_ ;
	wire _w9672_ ;
	wire _w9673_ ;
	wire _w9674_ ;
	wire _w9675_ ;
	wire _w9676_ ;
	wire _w9677_ ;
	wire _w9678_ ;
	wire _w9679_ ;
	wire _w9680_ ;
	wire _w9681_ ;
	wire _w9682_ ;
	wire _w9683_ ;
	wire _w9684_ ;
	wire _w9685_ ;
	wire _w9686_ ;
	wire _w9687_ ;
	wire _w9688_ ;
	wire _w9689_ ;
	wire _w9690_ ;
	wire _w9691_ ;
	wire _w9692_ ;
	wire _w9693_ ;
	wire _w9694_ ;
	wire _w9695_ ;
	wire _w9696_ ;
	wire _w9697_ ;
	wire _w9698_ ;
	wire _w9699_ ;
	wire _w9700_ ;
	wire _w9701_ ;
	wire _w9702_ ;
	wire _w9703_ ;
	wire _w9704_ ;
	wire _w9705_ ;
	wire _w9706_ ;
	wire _w9707_ ;
	wire _w9708_ ;
	wire _w9709_ ;
	wire _w9710_ ;
	wire _w9711_ ;
	wire _w9712_ ;
	wire _w9713_ ;
	wire _w9714_ ;
	wire _w9715_ ;
	wire _w9716_ ;
	wire _w9717_ ;
	wire _w9718_ ;
	wire _w9719_ ;
	wire _w9720_ ;
	wire _w9721_ ;
	wire _w9722_ ;
	wire _w9723_ ;
	wire _w9724_ ;
	wire _w9725_ ;
	wire _w9726_ ;
	wire _w9727_ ;
	wire _w9728_ ;
	wire _w9729_ ;
	wire _w9730_ ;
	wire _w9731_ ;
	wire _w9732_ ;
	wire _w9733_ ;
	wire _w9734_ ;
	wire _w9735_ ;
	wire _w9736_ ;
	wire _w9737_ ;
	wire _w9738_ ;
	wire _w9739_ ;
	wire _w9740_ ;
	wire _w9741_ ;
	wire _w9742_ ;
	wire _w9743_ ;
	wire _w9744_ ;
	wire _w9745_ ;
	wire _w9746_ ;
	wire _w9747_ ;
	wire _w9748_ ;
	wire _w9749_ ;
	wire _w9750_ ;
	wire _w9751_ ;
	wire _w9752_ ;
	wire _w9753_ ;
	wire _w9754_ ;
	wire _w9755_ ;
	wire _w9756_ ;
	wire _w9757_ ;
	wire _w9758_ ;
	wire _w9759_ ;
	wire _w9760_ ;
	wire _w9761_ ;
	wire _w9762_ ;
	wire _w9763_ ;
	wire _w9764_ ;
	wire _w9765_ ;
	wire _w9766_ ;
	wire _w9767_ ;
	wire _w9768_ ;
	wire _w9769_ ;
	wire _w9770_ ;
	wire _w9771_ ;
	wire _w9772_ ;
	wire _w9773_ ;
	wire _w9774_ ;
	wire _w9775_ ;
	wire _w9776_ ;
	wire _w9777_ ;
	wire _w9778_ ;
	wire _w9779_ ;
	wire _w9780_ ;
	wire _w9781_ ;
	wire _w9782_ ;
	wire _w9783_ ;
	wire _w9784_ ;
	wire _w9785_ ;
	wire _w9786_ ;
	wire _w9787_ ;
	wire _w9788_ ;
	wire _w9789_ ;
	wire _w9790_ ;
	wire _w9791_ ;
	wire _w9792_ ;
	wire _w9793_ ;
	wire _w9794_ ;
	wire _w9795_ ;
	wire _w9796_ ;
	wire _w9797_ ;
	wire _w9798_ ;
	wire _w9799_ ;
	wire _w9800_ ;
	wire _w9801_ ;
	wire _w9802_ ;
	wire _w9803_ ;
	wire _w9804_ ;
	wire _w9805_ ;
	wire _w9806_ ;
	wire _w9807_ ;
	wire _w9808_ ;
	wire _w9809_ ;
	wire _w9810_ ;
	wire _w9811_ ;
	wire _w9812_ ;
	wire _w9813_ ;
	wire _w9814_ ;
	wire _w9815_ ;
	wire _w9816_ ;
	wire _w9817_ ;
	wire _w9818_ ;
	wire _w9819_ ;
	wire _w9820_ ;
	wire _w9821_ ;
	wire _w9822_ ;
	wire _w9823_ ;
	wire _w9824_ ;
	wire _w9825_ ;
	wire _w9826_ ;
	wire _w9827_ ;
	wire _w9828_ ;
	wire _w9829_ ;
	wire _w9830_ ;
	wire _w9831_ ;
	wire _w9832_ ;
	wire _w9833_ ;
	wire _w9834_ ;
	wire _w9835_ ;
	wire _w9836_ ;
	wire _w9837_ ;
	wire _w9838_ ;
	wire _w9839_ ;
	wire _w9840_ ;
	wire _w9841_ ;
	wire _w9842_ ;
	wire _w9843_ ;
	wire _w9844_ ;
	wire _w9845_ ;
	wire _w9846_ ;
	wire _w9847_ ;
	wire _w9848_ ;
	wire _w9849_ ;
	wire _w9850_ ;
	wire _w9851_ ;
	wire _w9852_ ;
	wire _w9853_ ;
	wire _w9854_ ;
	wire _w9855_ ;
	wire _w9856_ ;
	wire _w9857_ ;
	wire _w9858_ ;
	wire _w9859_ ;
	wire _w9860_ ;
	wire _w9861_ ;
	wire _w9862_ ;
	wire _w9863_ ;
	wire _w9864_ ;
	wire _w9865_ ;
	wire _w9866_ ;
	wire _w9867_ ;
	wire _w9868_ ;
	wire _w9869_ ;
	wire _w9870_ ;
	wire _w9871_ ;
	wire _w9872_ ;
	wire _w9873_ ;
	wire _w9874_ ;
	wire _w9875_ ;
	wire _w9876_ ;
	wire _w9877_ ;
	wire _w9878_ ;
	wire _w9879_ ;
	wire _w9880_ ;
	wire _w9881_ ;
	wire _w9882_ ;
	wire _w9883_ ;
	wire _w9884_ ;
	wire _w9885_ ;
	wire _w9886_ ;
	wire _w9887_ ;
	wire _w9888_ ;
	wire _w9889_ ;
	wire _w9890_ ;
	wire _w9891_ ;
	wire _w9892_ ;
	wire _w9893_ ;
	wire _w9894_ ;
	wire _w9895_ ;
	wire _w9896_ ;
	wire _w9897_ ;
	wire _w9898_ ;
	wire _w9899_ ;
	wire _w9900_ ;
	wire _w9901_ ;
	wire _w9902_ ;
	wire _w9903_ ;
	wire _w9904_ ;
	wire _w9905_ ;
	wire _w9906_ ;
	wire _w9907_ ;
	wire _w9908_ ;
	wire _w9909_ ;
	wire _w9910_ ;
	wire _w9911_ ;
	wire _w9912_ ;
	wire _w9913_ ;
	wire _w9914_ ;
	wire _w9915_ ;
	wire _w9916_ ;
	wire _w9917_ ;
	wire _w9918_ ;
	wire _w9919_ ;
	wire _w9920_ ;
	wire _w9921_ ;
	wire _w9922_ ;
	wire _w9923_ ;
	wire _w9924_ ;
	wire _w9925_ ;
	wire _w9926_ ;
	wire _w9927_ ;
	wire _w9928_ ;
	wire _w9929_ ;
	wire _w9930_ ;
	wire _w9931_ ;
	wire _w9932_ ;
	wire _w9933_ ;
	wire _w9934_ ;
	wire _w9935_ ;
	wire _w9936_ ;
	wire _w9937_ ;
	wire _w9938_ ;
	wire _w9939_ ;
	wire _w9940_ ;
	wire _w9941_ ;
	wire _w9942_ ;
	wire _w9943_ ;
	wire _w9944_ ;
	wire _w9945_ ;
	wire _w9946_ ;
	wire _w9947_ ;
	wire _w9948_ ;
	wire _w9949_ ;
	wire _w9950_ ;
	wire _w9951_ ;
	wire _w9952_ ;
	wire _w9953_ ;
	wire _w9954_ ;
	wire _w9955_ ;
	wire _w9956_ ;
	wire _w9957_ ;
	wire _w9958_ ;
	wire _w9959_ ;
	wire _w9960_ ;
	wire _w9961_ ;
	wire _w9962_ ;
	wire _w9963_ ;
	wire _w9964_ ;
	wire _w9965_ ;
	wire _w9966_ ;
	wire _w9967_ ;
	wire _w9968_ ;
	wire _w9969_ ;
	wire _w9970_ ;
	wire _w9971_ ;
	wire _w9972_ ;
	wire _w9973_ ;
	wire _w9974_ ;
	wire _w9975_ ;
	wire _w9976_ ;
	wire _w9977_ ;
	wire _w9978_ ;
	wire _w9979_ ;
	wire _w9980_ ;
	wire _w9981_ ;
	wire _w9982_ ;
	wire _w9983_ ;
	wire _w9984_ ;
	wire _w9985_ ;
	wire _w9986_ ;
	wire _w9987_ ;
	wire _w9988_ ;
	wire _w9989_ ;
	wire _w9990_ ;
	wire _w9991_ ;
	wire _w9992_ ;
	wire _w9993_ ;
	wire _w9994_ ;
	wire _w9995_ ;
	wire _w9996_ ;
	wire _w9997_ ;
	wire _w9998_ ;
	wire _w9999_ ;
	wire _w10000_ ;
	wire _w10001_ ;
	wire _w10002_ ;
	wire _w10003_ ;
	wire _w10004_ ;
	wire _w10005_ ;
	wire _w10006_ ;
	wire _w10007_ ;
	wire _w10008_ ;
	wire _w10009_ ;
	wire _w10010_ ;
	wire _w10011_ ;
	wire _w10012_ ;
	wire _w10013_ ;
	wire _w10014_ ;
	wire _w10015_ ;
	wire _w10016_ ;
	wire _w10017_ ;
	wire _w10018_ ;
	wire _w10019_ ;
	wire _w10020_ ;
	wire _w10021_ ;
	wire _w10022_ ;
	wire _w10023_ ;
	wire _w10024_ ;
	wire _w10025_ ;
	wire _w10026_ ;
	wire _w10027_ ;
	wire _w10028_ ;
	wire _w10029_ ;
	wire _w10030_ ;
	wire _w10031_ ;
	wire _w10032_ ;
	wire _w10033_ ;
	wire _w10034_ ;
	wire _w10035_ ;
	wire _w10036_ ;
	wire _w10037_ ;
	wire _w10038_ ;
	wire _w10039_ ;
	wire _w10040_ ;
	wire _w10041_ ;
	wire _w10042_ ;
	wire _w10043_ ;
	wire _w10044_ ;
	wire _w10045_ ;
	wire _w10046_ ;
	wire _w10047_ ;
	wire _w10048_ ;
	wire _w10049_ ;
	wire _w10050_ ;
	wire _w10051_ ;
	wire _w10052_ ;
	wire _w10053_ ;
	wire _w10054_ ;
	wire _w10055_ ;
	wire _w10056_ ;
	wire _w10057_ ;
	wire _w10058_ ;
	wire _w10059_ ;
	wire _w10060_ ;
	wire _w10061_ ;
	wire _w10062_ ;
	wire _w10063_ ;
	wire _w10064_ ;
	wire _w10065_ ;
	wire _w10066_ ;
	wire _w10067_ ;
	wire _w10068_ ;
	wire _w10069_ ;
	wire _w10070_ ;
	wire _w10071_ ;
	wire _w10072_ ;
	wire _w10073_ ;
	wire _w10074_ ;
	wire _w10075_ ;
	wire _w10076_ ;
	wire _w10077_ ;
	wire _w10078_ ;
	wire _w10079_ ;
	wire _w10080_ ;
	wire _w10081_ ;
	wire _w10082_ ;
	wire _w10083_ ;
	wire _w10084_ ;
	wire _w10085_ ;
	wire _w10086_ ;
	wire _w10087_ ;
	wire _w10088_ ;
	wire _w10089_ ;
	wire _w10090_ ;
	wire _w10091_ ;
	wire _w10092_ ;
	wire _w10093_ ;
	wire _w10094_ ;
	wire _w10095_ ;
	wire _w10096_ ;
	wire _w10097_ ;
	wire _w10098_ ;
	wire _w10099_ ;
	wire _w10100_ ;
	wire _w10101_ ;
	wire _w10102_ ;
	wire _w10103_ ;
	wire _w10104_ ;
	wire _w10105_ ;
	wire _w10106_ ;
	wire _w10107_ ;
	wire _w10108_ ;
	wire _w10109_ ;
	wire _w10110_ ;
	wire _w10111_ ;
	wire _w10112_ ;
	wire _w10113_ ;
	wire _w10114_ ;
	wire _w10115_ ;
	wire _w10116_ ;
	wire _w10117_ ;
	wire _w10118_ ;
	wire _w10119_ ;
	wire _w10120_ ;
	wire _w10121_ ;
	wire _w10122_ ;
	wire _w10123_ ;
	wire _w10124_ ;
	wire _w10125_ ;
	wire _w10126_ ;
	wire _w10127_ ;
	wire _w10128_ ;
	wire _w10129_ ;
	wire _w10130_ ;
	wire _w10131_ ;
	wire _w10132_ ;
	wire _w10133_ ;
	wire _w10134_ ;
	wire _w10135_ ;
	wire _w10136_ ;
	wire _w10137_ ;
	wire _w10138_ ;
	wire _w10139_ ;
	wire _w10140_ ;
	wire _w10141_ ;
	wire _w10142_ ;
	wire _w10143_ ;
	wire _w10144_ ;
	wire _w10145_ ;
	wire _w10146_ ;
	wire _w10147_ ;
	wire _w10148_ ;
	wire _w10149_ ;
	wire _w10150_ ;
	wire _w10151_ ;
	wire _w10152_ ;
	wire _w10153_ ;
	wire _w10154_ ;
	wire _w10155_ ;
	wire _w10156_ ;
	wire _w10157_ ;
	wire _w10158_ ;
	wire _w10159_ ;
	wire _w10160_ ;
	wire _w10161_ ;
	wire _w10162_ ;
	wire _w10163_ ;
	wire _w10164_ ;
	wire _w10165_ ;
	wire _w10166_ ;
	wire _w10167_ ;
	wire _w10168_ ;
	wire _w10169_ ;
	wire _w10170_ ;
	wire _w10171_ ;
	wire _w10172_ ;
	wire _w10173_ ;
	wire _w10174_ ;
	wire _w10175_ ;
	wire _w10176_ ;
	wire _w10177_ ;
	wire _w10178_ ;
	wire _w10179_ ;
	wire _w10180_ ;
	wire _w10181_ ;
	wire _w10182_ ;
	wire _w10183_ ;
	wire _w10184_ ;
	wire _w10185_ ;
	wire _w10186_ ;
	wire _w10187_ ;
	wire _w10188_ ;
	wire _w10189_ ;
	wire _w10190_ ;
	wire _w10191_ ;
	wire _w10192_ ;
	wire _w10193_ ;
	wire _w10194_ ;
	wire _w10195_ ;
	wire _w10196_ ;
	wire _w10197_ ;
	wire _w10198_ ;
	wire _w10199_ ;
	wire _w10200_ ;
	wire _w10201_ ;
	wire _w10202_ ;
	wire _w10203_ ;
	wire _w10204_ ;
	wire _w10205_ ;
	wire _w10206_ ;
	wire _w10207_ ;
	wire _w10208_ ;
	wire _w10209_ ;
	wire _w10210_ ;
	wire _w10211_ ;
	wire _w10212_ ;
	wire _w10213_ ;
	wire _w10214_ ;
	wire _w10215_ ;
	wire _w10216_ ;
	wire _w10217_ ;
	wire _w10218_ ;
	wire _w10219_ ;
	wire _w10220_ ;
	wire _w10221_ ;
	wire _w10222_ ;
	wire _w10223_ ;
	wire _w10224_ ;
	wire _w10225_ ;
	wire _w10226_ ;
	wire _w10227_ ;
	wire _w10228_ ;
	wire _w10229_ ;
	wire _w10230_ ;
	wire _w10231_ ;
	wire _w10232_ ;
	wire _w10233_ ;
	wire _w10234_ ;
	wire _w10235_ ;
	wire _w10236_ ;
	wire _w10237_ ;
	wire _w10238_ ;
	wire _w10239_ ;
	wire _w10240_ ;
	wire _w10241_ ;
	wire _w10242_ ;
	wire _w10243_ ;
	wire _w10244_ ;
	wire _w10245_ ;
	wire _w10246_ ;
	wire _w10247_ ;
	wire _w10248_ ;
	wire _w10249_ ;
	wire _w10250_ ;
	wire _w10251_ ;
	wire _w10252_ ;
	wire _w10253_ ;
	wire _w10254_ ;
	wire _w10255_ ;
	wire _w10256_ ;
	wire _w10257_ ;
	wire _w10258_ ;
	wire _w10259_ ;
	wire _w10260_ ;
	wire _w10261_ ;
	wire _w10262_ ;
	wire _w10263_ ;
	wire _w10264_ ;
	wire _w10265_ ;
	wire _w10266_ ;
	wire _w10267_ ;
	wire _w10268_ ;
	wire _w10269_ ;
	wire _w10270_ ;
	wire _w10271_ ;
	wire _w10272_ ;
	wire _w10273_ ;
	wire _w10274_ ;
	wire _w10275_ ;
	wire _w10276_ ;
	wire _w10277_ ;
	wire _w10278_ ;
	wire _w10279_ ;
	wire _w10280_ ;
	wire _w10281_ ;
	wire _w10282_ ;
	wire _w10283_ ;
	wire _w10284_ ;
	wire _w10285_ ;
	wire _w10286_ ;
	wire _w10287_ ;
	wire _w10288_ ;
	wire _w10289_ ;
	wire _w10290_ ;
	wire _w10291_ ;
	wire _w10292_ ;
	wire _w10293_ ;
	wire _w10294_ ;
	wire _w10295_ ;
	wire _w10296_ ;
	wire _w10297_ ;
	wire _w10298_ ;
	wire _w10299_ ;
	wire _w10300_ ;
	wire _w10301_ ;
	wire _w10302_ ;
	wire _w10303_ ;
	wire _w10304_ ;
	wire _w10305_ ;
	wire _w10306_ ;
	LUT2 #(
		.INIT('h9)
	) name0 (
		\a[2] ,
		\a[3] ,
		_w34_
	);
	LUT4 #(
		.INIT('h0660)
	) name1 (
		\a[2] ,
		\a[3] ,
		\a[4] ,
		\a[5] ,
		_w35_
	);
	LUT2 #(
		.INIT('h9)
	) name2 (
		\a[20] ,
		\a[21] ,
		_w36_
	);
	LUT4 #(
		.INIT('h0660)
	) name3 (
		\a[20] ,
		\a[21] ,
		\a[22] ,
		\a[23] ,
		_w37_
	);
	LUT4 #(
		.INIT('h0010)
	) name4 (
		\a[23] ,
		\a[24] ,
		\a[25] ,
		\a[26] ,
		_w38_
	);
	LUT4 #(
		.INIT('h0040)
	) name5 (
		\a[27] ,
		\a[28] ,
		\a[29] ,
		\a[30] ,
		_w39_
	);
	LUT2 #(
		.INIT('h8)
	) name6 (
		_w38_,
		_w39_,
		_w40_
	);
	LUT4 #(
		.INIT('h4000)
	) name7 (
		\a[23] ,
		\a[24] ,
		\a[25] ,
		\a[26] ,
		_w41_
	);
	LUT3 #(
		.INIT('h1f)
	) name8 (
		_w38_,
		_w41_,
		_w39_,
		_w42_
	);
	LUT4 #(
		.INIT('h0020)
	) name9 (
		\a[27] ,
		\a[28] ,
		\a[29] ,
		\a[30] ,
		_w43_
	);
	LUT4 #(
		.INIT('h0400)
	) name10 (
		\a[23] ,
		\a[24] ,
		\a[25] ,
		\a[26] ,
		_w44_
	);
	LUT2 #(
		.INIT('h8)
	) name11 (
		_w43_,
		_w44_,
		_w45_
	);
	LUT4 #(
		.INIT('h8000)
	) name12 (
		\a[23] ,
		\a[24] ,
		\a[25] ,
		\a[26] ,
		_w46_
	);
	LUT4 #(
		.INIT('h0002)
	) name13 (
		\a[23] ,
		\a[24] ,
		\a[25] ,
		\a[26] ,
		_w47_
	);
	LUT4 #(
		.INIT('h135f)
	) name14 (
		_w47_,
		_w39_,
		_w43_,
		_w46_,
		_w48_
	);
	LUT3 #(
		.INIT('h40)
	) name15 (
		_w45_,
		_w48_,
		_w42_,
		_w49_
	);
	LUT4 #(
		.INIT('h0800)
	) name16 (
		\a[23] ,
		\a[24] ,
		\a[25] ,
		\a[26] ,
		_w50_
	);
	LUT2 #(
		.INIT('h8)
	) name17 (
		_w50_,
		_w43_,
		_w51_
	);
	LUT4 #(
		.INIT('h0040)
	) name18 (
		\a[23] ,
		\a[24] ,
		\a[25] ,
		\a[26] ,
		_w52_
	);
	LUT2 #(
		.INIT('h8)
	) name19 (
		_w52_,
		_w43_,
		_w53_
	);
	LUT3 #(
		.INIT('h1f)
	) name20 (
		_w52_,
		_w50_,
		_w43_,
		_w54_
	);
	LUT4 #(
		.INIT('h0020)
	) name21 (
		\a[23] ,
		\a[24] ,
		\a[25] ,
		\a[26] ,
		_w55_
	);
	LUT4 #(
		.INIT('h2000)
	) name22 (
		\a[23] ,
		\a[24] ,
		\a[25] ,
		\a[26] ,
		_w56_
	);
	LUT2 #(
		.INIT('h8)
	) name23 (
		_w56_,
		_w39_,
		_w57_
	);
	LUT3 #(
		.INIT('h1f)
	) name24 (
		_w55_,
		_w56_,
		_w39_,
		_w58_
	);
	LUT4 #(
		.INIT('h0100)
	) name25 (
		\a[23] ,
		\a[24] ,
		\a[25] ,
		\a[26] ,
		_w59_
	);
	LUT2 #(
		.INIT('h8)
	) name26 (
		_w59_,
		_w43_,
		_w60_
	);
	LUT2 #(
		.INIT('h8)
	) name27 (
		_w52_,
		_w39_,
		_w61_
	);
	LUT4 #(
		.INIT('h135f)
	) name28 (
		_w52_,
		_w59_,
		_w39_,
		_w43_,
		_w62_
	);
	LUT3 #(
		.INIT('h80)
	) name29 (
		_w58_,
		_w54_,
		_w62_,
		_w63_
	);
	LUT2 #(
		.INIT('h8)
	) name30 (
		_w43_,
		_w46_,
		_w64_
	);
	LUT4 #(
		.INIT('h0001)
	) name31 (
		\a[23] ,
		\a[24] ,
		\a[25] ,
		\a[26] ,
		_w65_
	);
	LUT3 #(
		.INIT('h37)
	) name32 (
		_w47_,
		_w39_,
		_w65_,
		_w66_
	);
	LUT4 #(
		.INIT('h0008)
	) name33 (
		\a[23] ,
		\a[24] ,
		\a[25] ,
		\a[26] ,
		_w67_
	);
	LUT3 #(
		.INIT('h37)
	) name34 (
		_w67_,
		_w39_,
		_w44_,
		_w68_
	);
	LUT2 #(
		.INIT('h8)
	) name35 (
		_w41_,
		_w43_,
		_w69_
	);
	LUT3 #(
		.INIT('h1f)
	) name36 (
		_w38_,
		_w41_,
		_w43_,
		_w70_
	);
	LUT4 #(
		.INIT('h4000)
	) name37 (
		_w64_,
		_w66_,
		_w68_,
		_w70_,
		_w71_
	);
	LUT4 #(
		.INIT('h0010)
	) name38 (
		\a[27] ,
		\a[28] ,
		\a[29] ,
		\a[30] ,
		_w72_
	);
	LUT2 #(
		.INIT('h8)
	) name39 (
		_w72_,
		_w44_,
		_w73_
	);
	LUT2 #(
		.INIT('h8)
	) name40 (
		_w43_,
		_w65_,
		_w74_
	);
	LUT4 #(
		.INIT('h153f)
	) name41 (
		_w72_,
		_w43_,
		_w65_,
		_w44_,
		_w75_
	);
	LUT4 #(
		.INIT('h8000)
	) name42 (
		_w49_,
		_w63_,
		_w71_,
		_w75_,
		_w76_
	);
	LUT2 #(
		.INIT('h8)
	) name43 (
		_w67_,
		_w72_,
		_w77_
	);
	LUT4 #(
		.INIT('h0008)
	) name44 (
		\a[27] ,
		\a[28] ,
		\a[29] ,
		\a[30] ,
		_w78_
	);
	LUT2 #(
		.INIT('h8)
	) name45 (
		_w78_,
		_w41_,
		_w79_
	);
	LUT2 #(
		.INIT('h8)
	) name46 (
		_w47_,
		_w72_,
		_w80_
	);
	LUT4 #(
		.INIT('h135f)
	) name47 (
		_w78_,
		_w47_,
		_w41_,
		_w72_,
		_w81_
	);
	LUT2 #(
		.INIT('h4)
	) name48 (
		_w77_,
		_w81_,
		_w82_
	);
	LUT2 #(
		.INIT('h8)
	) name49 (
		_w72_,
		_w46_,
		_w83_
	);
	LUT2 #(
		.INIT('h8)
	) name50 (
		_w55_,
		_w72_,
		_w84_
	);
	LUT4 #(
		.INIT('h0080)
	) name51 (
		\a[23] ,
		\a[24] ,
		\a[25] ,
		\a[26] ,
		_w85_
	);
	LUT2 #(
		.INIT('h8)
	) name52 (
		_w85_,
		_w72_,
		_w86_
	);
	LUT3 #(
		.INIT('h1f)
	) name53 (
		_w55_,
		_w85_,
		_w72_,
		_w87_
	);
	LUT4 #(
		.INIT('h0f1f)
	) name54 (
		_w55_,
		_w85_,
		_w72_,
		_w46_,
		_w88_
	);
	LUT4 #(
		.INIT('h153f)
	) name55 (
		_w78_,
		_w72_,
		_w65_,
		_w46_,
		_w89_
	);
	LUT4 #(
		.INIT('h0200)
	) name56 (
		\a[23] ,
		\a[24] ,
		\a[25] ,
		\a[26] ,
		_w90_
	);
	LUT2 #(
		.INIT('h8)
	) name57 (
		_w90_,
		_w72_,
		_w91_
	);
	LUT3 #(
		.INIT('h08)
	) name58 (
		_w89_,
		_w88_,
		_w91_,
		_w92_
	);
	LUT4 #(
		.INIT('h1000)
	) name59 (
		\a[23] ,
		\a[24] ,
		\a[25] ,
		\a[26] ,
		_w93_
	);
	LUT2 #(
		.INIT('h8)
	) name60 (
		_w72_,
		_w93_,
		_w94_
	);
	LUT3 #(
		.INIT('h57)
	) name61 (
		_w72_,
		_w50_,
		_w93_,
		_w95_
	);
	LUT3 #(
		.INIT('h1f)
	) name62 (
		_w38_,
		_w59_,
		_w72_,
		_w96_
	);
	LUT2 #(
		.INIT('h8)
	) name63 (
		_w52_,
		_w72_,
		_w97_
	);
	LUT3 #(
		.INIT('h1f)
	) name64 (
		_w52_,
		_w56_,
		_w72_,
		_w98_
	);
	LUT3 #(
		.INIT('h80)
	) name65 (
		_w96_,
		_w95_,
		_w98_,
		_w99_
	);
	LUT3 #(
		.INIT('h80)
	) name66 (
		_w82_,
		_w92_,
		_w99_,
		_w100_
	);
	LUT2 #(
		.INIT('h8)
	) name67 (
		_w56_,
		_w43_,
		_w101_
	);
	LUT2 #(
		.INIT('h8)
	) name68 (
		_w90_,
		_w39_,
		_w102_
	);
	LUT3 #(
		.INIT('h1f)
	) name69 (
		_w85_,
		_w90_,
		_w39_,
		_w103_
	);
	LUT2 #(
		.INIT('h8)
	) name70 (
		_w90_,
		_w43_,
		_w104_
	);
	LUT3 #(
		.INIT('h37)
	) name71 (
		_w90_,
		_w43_,
		_w93_,
		_w105_
	);
	LUT4 #(
		.INIT('h0080)
	) name72 (
		\a[27] ,
		\a[28] ,
		\a[29] ,
		\a[30] ,
		_w106_
	);
	LUT2 #(
		.INIT('h8)
	) name73 (
		_w106_,
		_w65_,
		_w107_
	);
	LUT4 #(
		.INIT('h153f)
	) name74 (
		_w106_,
		_w67_,
		_w43_,
		_w65_,
		_w108_
	);
	LUT4 #(
		.INIT('h4000)
	) name75 (
		_w101_,
		_w105_,
		_w108_,
		_w103_,
		_w109_
	);
	LUT4 #(
		.INIT('h0004)
	) name76 (
		\a[23] ,
		\a[24] ,
		\a[25] ,
		\a[26] ,
		_w110_
	);
	LUT2 #(
		.INIT('h8)
	) name77 (
		_w110_,
		_w39_,
		_w111_
	);
	LUT3 #(
		.INIT('h57)
	) name78 (
		_w110_,
		_w39_,
		_w43_,
		_w112_
	);
	LUT4 #(
		.INIT('h1537)
	) name79 (
		_w110_,
		_w39_,
		_w50_,
		_w43_,
		_w113_
	);
	LUT2 #(
		.INIT('h8)
	) name80 (
		_w59_,
		_w39_,
		_w114_
	);
	LUT3 #(
		.INIT('h37)
	) name81 (
		_w59_,
		_w39_,
		_w93_,
		_w115_
	);
	LUT3 #(
		.INIT('h1f)
	) name82 (
		_w55_,
		_w85_,
		_w43_,
		_w116_
	);
	LUT3 #(
		.INIT('h80)
	) name83 (
		_w113_,
		_w115_,
		_w116_,
		_w117_
	);
	LUT2 #(
		.INIT('h8)
	) name84 (
		_w41_,
		_w72_,
		_w118_
	);
	LUT3 #(
		.INIT('h1f)
	) name85 (
		_w110_,
		_w41_,
		_w72_,
		_w119_
	);
	LUT3 #(
		.INIT('h80)
	) name86 (
		_w109_,
		_w117_,
		_w119_,
		_w120_
	);
	LUT3 #(
		.INIT('h80)
	) name87 (
		_w76_,
		_w100_,
		_w120_,
		_w121_
	);
	LUT4 #(
		.INIT('h0001)
	) name88 (
		\a[27] ,
		\a[28] ,
		\a[29] ,
		\a[30] ,
		_w122_
	);
	LUT3 #(
		.INIT('h57)
	) name89 (
		_w122_,
		_w55_,
		_w52_,
		_w123_
	);
	LUT2 #(
		.INIT('h8)
	) name90 (
		_w122_,
		_w110_,
		_w124_
	);
	LUT3 #(
		.INIT('h57)
	) name91 (
		_w122_,
		_w110_,
		_w67_,
		_w125_
	);
	LUT4 #(
		.INIT('h5557)
	) name92 (
		_w122_,
		_w59_,
		_w110_,
		_w67_,
		_w126_
	);
	LUT2 #(
		.INIT('h8)
	) name93 (
		_w123_,
		_w126_,
		_w127_
	);
	LUT2 #(
		.INIT('h8)
	) name94 (
		_w38_,
		_w122_,
		_w128_
	);
	LUT2 #(
		.INIT('h8)
	) name95 (
		_w106_,
		_w55_,
		_w129_
	);
	LUT3 #(
		.INIT('h57)
	) name96 (
		_w106_,
		_w55_,
		_w85_,
		_w130_
	);
	LUT4 #(
		.INIT('h5557)
	) name97 (
		_w106_,
		_w55_,
		_w85_,
		_w52_,
		_w131_
	);
	LUT3 #(
		.INIT('h37)
	) name98 (
		_w38_,
		_w106_,
		_w59_,
		_w132_
	);
	LUT3 #(
		.INIT('h40)
	) name99 (
		_w128_,
		_w131_,
		_w132_,
		_w133_
	);
	LUT2 #(
		.INIT('h8)
	) name100 (
		_w127_,
		_w133_,
		_w134_
	);
	LUT2 #(
		.INIT('h8)
	) name101 (
		_w59_,
		_w78_,
		_w135_
	);
	LUT4 #(
		.INIT('h0f1f)
	) name102 (
		_w55_,
		_w59_,
		_w78_,
		_w50_,
		_w136_
	);
	LUT2 #(
		.INIT('h8)
	) name103 (
		_w52_,
		_w78_,
		_w137_
	);
	LUT3 #(
		.INIT('h1f)
	) name104 (
		_w85_,
		_w52_,
		_w78_,
		_w138_
	);
	LUT3 #(
		.INIT('h57)
	) name105 (
		_w78_,
		_w93_,
		_w44_,
		_w139_
	);
	LUT3 #(
		.INIT('h80)
	) name106 (
		_w138_,
		_w139_,
		_w136_,
		_w140_
	);
	LUT2 #(
		.INIT('h8)
	) name107 (
		_w122_,
		_w65_,
		_w141_
	);
	LUT2 #(
		.INIT('h8)
	) name108 (
		_w106_,
		_w110_,
		_w142_
	);
	LUT3 #(
		.INIT('h57)
	) name109 (
		_w106_,
		_w67_,
		_w47_,
		_w143_
	);
	LUT4 #(
		.INIT('h5557)
	) name110 (
		_w106_,
		_w110_,
		_w67_,
		_w47_,
		_w144_
	);
	LUT2 #(
		.INIT('h4)
	) name111 (
		_w141_,
		_w144_,
		_w145_
	);
	LUT2 #(
		.INIT('h8)
	) name112 (
		_w122_,
		_w85_,
		_w146_
	);
	LUT2 #(
		.INIT('h8)
	) name113 (
		_w122_,
		_w90_,
		_w147_
	);
	LUT3 #(
		.INIT('h57)
	) name114 (
		_w122_,
		_w90_,
		_w47_,
		_w148_
	);
	LUT4 #(
		.INIT('h5557)
	) name115 (
		_w122_,
		_w85_,
		_w90_,
		_w47_,
		_w149_
	);
	LUT3 #(
		.INIT('h1f)
	) name116 (
		_w38_,
		_w67_,
		_w78_,
		_w150_
	);
	LUT2 #(
		.INIT('h8)
	) name117 (
		_w78_,
		_w90_,
		_w151_
	);
	LUT2 #(
		.INIT('h8)
	) name118 (
		_w78_,
		_w56_,
		_w152_
	);
	LUT3 #(
		.INIT('h57)
	) name119 (
		_w78_,
		_w90_,
		_w56_,
		_w153_
	);
	LUT3 #(
		.INIT('h80)
	) name120 (
		_w149_,
		_w150_,
		_w153_,
		_w154_
	);
	LUT3 #(
		.INIT('h80)
	) name121 (
		_w145_,
		_w140_,
		_w154_,
		_w155_
	);
	LUT2 #(
		.INIT('h8)
	) name122 (
		_w134_,
		_w155_,
		_w156_
	);
	LUT2 #(
		.INIT('h8)
	) name123 (
		_w121_,
		_w156_,
		_w157_
	);
	LUT4 #(
		.INIT('h8000)
	) name124 (
		\a[27] ,
		\a[28] ,
		\a[29] ,
		\a[30] ,
		_w158_
	);
	LUT2 #(
		.INIT('h8)
	) name125 (
		_w52_,
		_w158_,
		_w159_
	);
	LUT2 #(
		.INIT('h8)
	) name126 (
		_w67_,
		_w158_,
		_w160_
	);
	LUT2 #(
		.INIT('h8)
	) name127 (
		_w59_,
		_w158_,
		_w161_
	);
	LUT2 #(
		.INIT('h8)
	) name128 (
		_w85_,
		_w158_,
		_w162_
	);
	LUT4 #(
		.INIT('h01ff)
	) name129 (
		_w85_,
		_w59_,
		_w67_,
		_w158_,
		_w163_
	);
	LUT2 #(
		.INIT('h8)
	) name130 (
		_w55_,
		_w158_,
		_w164_
	);
	LUT2 #(
		.INIT('h8)
	) name131 (
		_w110_,
		_w158_,
		_w165_
	);
	LUT4 #(
		.INIT('h4000)
	) name132 (
		\a[27] ,
		\a[28] ,
		\a[29] ,
		\a[30] ,
		_w166_
	);
	LUT2 #(
		.INIT('h8)
	) name133 (
		_w56_,
		_w166_,
		_w167_
	);
	LUT4 #(
		.INIT('h153f)
	) name134 (
		_w110_,
		_w56_,
		_w166_,
		_w158_,
		_w168_
	);
	LUT2 #(
		.INIT('h8)
	) name135 (
		_w38_,
		_w158_,
		_w169_
	);
	LUT2 #(
		.INIT('h8)
	) name136 (
		_w47_,
		_w158_,
		_w170_
	);
	LUT3 #(
		.INIT('h1f)
	) name137 (
		_w38_,
		_w47_,
		_w158_,
		_w171_
	);
	LUT4 #(
		.INIT('h153f)
	) name138 (
		_w65_,
		_w46_,
		_w166_,
		_w158_,
		_w172_
	);
	LUT4 #(
		.INIT('h4000)
	) name139 (
		_w164_,
		_w168_,
		_w171_,
		_w172_,
		_w173_
	);
	LUT3 #(
		.INIT('h40)
	) name140 (
		_w159_,
		_w163_,
		_w173_,
		_w174_
	);
	LUT4 #(
		.INIT('h1000)
	) name141 (
		_w146_,
		_w159_,
		_w163_,
		_w173_,
		_w175_
	);
	LUT4 #(
		.INIT('h0004)
	) name142 (
		\a[27] ,
		\a[28] ,
		\a[29] ,
		\a[30] ,
		_w176_
	);
	LUT2 #(
		.INIT('h8)
	) name143 (
		_w85_,
		_w176_,
		_w177_
	);
	LUT2 #(
		.INIT('h2)
	) name144 (
		_w144_,
		_w177_,
		_w178_
	);
	LUT2 #(
		.INIT('h8)
	) name145 (
		_w175_,
		_w178_,
		_w179_
	);
	LUT2 #(
		.INIT('h8)
	) name146 (
		_w90_,
		_w166_,
		_w180_
	);
	LUT3 #(
		.INIT('h1f)
	) name147 (
		_w38_,
		_w90_,
		_w166_,
		_w181_
	);
	LUT2 #(
		.INIT('h8)
	) name148 (
		_w65_,
		_w166_,
		_w182_
	);
	LUT3 #(
		.INIT('h1f)
	) name149 (
		_w67_,
		_w65_,
		_w166_,
		_w183_
	);
	LUT4 #(
		.INIT('h2000)
	) name150 (
		\a[27] ,
		\a[28] ,
		\a[29] ,
		\a[30] ,
		_w184_
	);
	LUT2 #(
		.INIT('h8)
	) name151 (
		_w46_,
		_w184_,
		_w185_
	);
	LUT2 #(
		.INIT('h8)
	) name152 (
		_w59_,
		_w166_,
		_w186_
	);
	LUT4 #(
		.INIT('h153f)
	) name153 (
		_w59_,
		_w46_,
		_w184_,
		_w166_,
		_w187_
	);
	LUT3 #(
		.INIT('h80)
	) name154 (
		_w181_,
		_w183_,
		_w187_,
		_w188_
	);
	LUT2 #(
		.INIT('h8)
	) name155 (
		_w41_,
		_w184_,
		_w189_
	);
	LUT2 #(
		.INIT('h8)
	) name156 (
		_w93_,
		_w184_,
		_w190_
	);
	LUT4 #(
		.INIT('h153f)
	) name157 (
		_w47_,
		_w93_,
		_w184_,
		_w166_,
		_w191_
	);
	LUT2 #(
		.INIT('h4)
	) name158 (
		_w189_,
		_w191_,
		_w192_
	);
	LUT2 #(
		.INIT('h8)
	) name159 (
		_w50_,
		_w166_,
		_w193_
	);
	LUT2 #(
		.INIT('h8)
	) name160 (
		_w85_,
		_w166_,
		_w194_
	);
	LUT4 #(
		.INIT('h153f)
	) name161 (
		_w85_,
		_w56_,
		_w184_,
		_w166_,
		_w195_
	);
	LUT3 #(
		.INIT('h1f)
	) name162 (
		_w55_,
		_w52_,
		_w166_,
		_w196_
	);
	LUT2 #(
		.INIT('h8)
	) name163 (
		_w110_,
		_w166_,
		_w197_
	);
	LUT3 #(
		.INIT('h1f)
	) name164 (
		_w110_,
		_w44_,
		_w166_,
		_w198_
	);
	LUT4 #(
		.INIT('h0800)
	) name165 (
		_w196_,
		_w198_,
		_w193_,
		_w195_,
		_w199_
	);
	LUT3 #(
		.INIT('h80)
	) name166 (
		_w192_,
		_w188_,
		_w199_,
		_w200_
	);
	LUT4 #(
		.INIT('h1000)
	) name167 (
		\a[27] ,
		\a[28] ,
		\a[29] ,
		\a[30] ,
		_w201_
	);
	LUT2 #(
		.INIT('h8)
	) name168 (
		_w46_,
		_w201_,
		_w202_
	);
	LUT2 #(
		.INIT('h8)
	) name169 (
		_w44_,
		_w201_,
		_w203_
	);
	LUT3 #(
		.INIT('h1f)
	) name170 (
		_w44_,
		_w46_,
		_w201_,
		_w204_
	);
	LUT2 #(
		.INIT('h8)
	) name171 (
		_w38_,
		_w184_,
		_w205_
	);
	LUT2 #(
		.INIT('h8)
	) name172 (
		_w50_,
		_w201_,
		_w206_
	);
	LUT4 #(
		.INIT('h135f)
	) name173 (
		_w38_,
		_w50_,
		_w184_,
		_w201_,
		_w207_
	);
	LUT2 #(
		.INIT('h8)
	) name174 (
		_w204_,
		_w207_,
		_w208_
	);
	LUT2 #(
		.INIT('h8)
	) name175 (
		_w52_,
		_w184_,
		_w209_
	);
	LUT2 #(
		.INIT('h8)
	) name176 (
		_w50_,
		_w184_,
		_w210_
	);
	LUT3 #(
		.INIT('h1f)
	) name177 (
		_w52_,
		_w50_,
		_w184_,
		_w211_
	);
	LUT2 #(
		.INIT('h8)
	) name178 (
		_w90_,
		_w184_,
		_w212_
	);
	LUT3 #(
		.INIT('h1f)
	) name179 (
		_w55_,
		_w90_,
		_w184_,
		_w213_
	);
	LUT2 #(
		.INIT('h8)
	) name180 (
		_w41_,
		_w201_,
		_w214_
	);
	LUT2 #(
		.INIT('h8)
	) name181 (
		_w110_,
		_w184_,
		_w215_
	);
	LUT4 #(
		.INIT('h135f)
	) name182 (
		_w110_,
		_w41_,
		_w184_,
		_w201_,
		_w216_
	);
	LUT3 #(
		.INIT('h80)
	) name183 (
		_w213_,
		_w216_,
		_w211_,
		_w217_
	);
	LUT2 #(
		.INIT('h8)
	) name184 (
		_w56_,
		_w201_,
		_w218_
	);
	LUT4 #(
		.INIT('h135f)
	) name185 (
		_w85_,
		_w56_,
		_w184_,
		_w201_,
		_w219_
	);
	LUT2 #(
		.INIT('h8)
	) name186 (
		_w59_,
		_w201_,
		_w220_
	);
	LUT2 #(
		.INIT('h8)
	) name187 (
		_w44_,
		_w184_,
		_w221_
	);
	LUT4 #(
		.INIT('h153f)
	) name188 (
		_w59_,
		_w44_,
		_w184_,
		_w201_,
		_w222_
	);
	LUT2 #(
		.INIT('h8)
	) name189 (
		_w67_,
		_w184_,
		_w223_
	);
	LUT2 #(
		.INIT('h8)
	) name190 (
		_w65_,
		_w184_,
		_w224_
	);
	LUT3 #(
		.INIT('h1f)
	) name191 (
		_w67_,
		_w65_,
		_w184_,
		_w225_
	);
	LUT2 #(
		.INIT('h8)
	) name192 (
		_w59_,
		_w184_,
		_w226_
	);
	LUT2 #(
		.INIT('h8)
	) name193 (
		_w93_,
		_w201_,
		_w227_
	);
	LUT4 #(
		.INIT('h135f)
	) name194 (
		_w59_,
		_w93_,
		_w184_,
		_w201_,
		_w228_
	);
	LUT4 #(
		.INIT('h8000)
	) name195 (
		_w225_,
		_w219_,
		_w222_,
		_w228_,
		_w229_
	);
	LUT2 #(
		.INIT('h8)
	) name196 (
		_w90_,
		_w201_,
		_w230_
	);
	LUT4 #(
		.INIT('h153f)
	) name197 (
		_w90_,
		_w47_,
		_w184_,
		_w201_,
		_w231_
	);
	LUT3 #(
		.INIT('h57)
	) name198 (
		_w122_,
		_w47_,
		_w65_,
		_w232_
	);
	LUT3 #(
		.INIT('h80)
	) name199 (
		_w125_,
		_w231_,
		_w232_,
		_w233_
	);
	LUT4 #(
		.INIT('h8000)
	) name200 (
		_w208_,
		_w217_,
		_w229_,
		_w233_,
		_w234_
	);
	LUT2 #(
		.INIT('h8)
	) name201 (
		_w55_,
		_w201_,
		_w235_
	);
	LUT4 #(
		.INIT('h0800)
	) name202 (
		\a[27] ,
		\a[28] ,
		\a[29] ,
		\a[30] ,
		_w236_
	);
	LUT2 #(
		.INIT('h8)
	) name203 (
		_w41_,
		_w236_,
		_w237_
	);
	LUT4 #(
		.INIT('h135f)
	) name204 (
		_w55_,
		_w41_,
		_w201_,
		_w236_,
		_w238_
	);
	LUT2 #(
		.INIT('h8)
	) name205 (
		_w93_,
		_w236_,
		_w239_
	);
	LUT4 #(
		.INIT('h135f)
	) name206 (
		_w38_,
		_w93_,
		_w201_,
		_w236_,
		_w240_
	);
	LUT2 #(
		.INIT('h8)
	) name207 (
		_w46_,
		_w236_,
		_w241_
	);
	LUT3 #(
		.INIT('h08)
	) name208 (
		_w240_,
		_w238_,
		_w241_,
		_w242_
	);
	LUT2 #(
		.INIT('h8)
	) name209 (
		_w52_,
		_w201_,
		_w243_
	);
	LUT2 #(
		.INIT('h8)
	) name210 (
		_w65_,
		_w201_,
		_w244_
	);
	LUT3 #(
		.INIT('h1f)
	) name211 (
		_w52_,
		_w65_,
		_w201_,
		_w245_
	);
	LUT2 #(
		.INIT('h8)
	) name212 (
		_w67_,
		_w201_,
		_w246_
	);
	LUT2 #(
		.INIT('h8)
	) name213 (
		_w110_,
		_w201_,
		_w247_
	);
	LUT3 #(
		.INIT('h1f)
	) name214 (
		_w110_,
		_w67_,
		_w201_,
		_w248_
	);
	LUT2 #(
		.INIT('h8)
	) name215 (
		_w245_,
		_w248_,
		_w249_
	);
	LUT2 #(
		.INIT('h8)
	) name216 (
		_w56_,
		_w236_,
		_w250_
	);
	LUT2 #(
		.INIT('h8)
	) name217 (
		_w85_,
		_w201_,
		_w251_
	);
	LUT4 #(
		.INIT('h135f)
	) name218 (
		_w85_,
		_w56_,
		_w201_,
		_w236_,
		_w252_
	);
	LUT2 #(
		.INIT('h8)
	) name219 (
		_w47_,
		_w201_,
		_w253_
	);
	LUT4 #(
		.INIT('h135f)
	) name220 (
		_w47_,
		_w50_,
		_w201_,
		_w236_,
		_w254_
	);
	LUT3 #(
		.INIT('h40)
	) name221 (
		_w128_,
		_w252_,
		_w254_,
		_w255_
	);
	LUT3 #(
		.INIT('h80)
	) name222 (
		_w242_,
		_w249_,
		_w255_,
		_w256_
	);
	LUT3 #(
		.INIT('h80)
	) name223 (
		_w234_,
		_w200_,
		_w256_,
		_w257_
	);
	LUT2 #(
		.INIT('h8)
	) name224 (
		_w41_,
		_w176_,
		_w258_
	);
	LUT4 #(
		.INIT('h0002)
	) name225 (
		\a[27] ,
		\a[28] ,
		\a[29] ,
		\a[30] ,
		_w259_
	);
	LUT4 #(
		.INIT('h135f)
	) name226 (
		_w56_,
		_w41_,
		_w259_,
		_w176_,
		_w260_
	);
	LUT2 #(
		.INIT('h8)
	) name227 (
		_w65_,
		_w176_,
		_w261_
	);
	LUT4 #(
		.INIT('h153f)
	) name228 (
		_w65_,
		_w46_,
		_w259_,
		_w176_,
		_w262_
	);
	LUT2 #(
		.INIT('h8)
	) name229 (
		_w38_,
		_w176_,
		_w263_
	);
	LUT2 #(
		.INIT('h8)
	) name230 (
		_w52_,
		_w176_,
		_w264_
	);
	LUT3 #(
		.INIT('h1f)
	) name231 (
		_w38_,
		_w52_,
		_w176_,
		_w265_
	);
	LUT3 #(
		.INIT('h80)
	) name232 (
		_w262_,
		_w265_,
		_w260_,
		_w266_
	);
	LUT2 #(
		.INIT('h8)
	) name233 (
		_w93_,
		_w176_,
		_w267_
	);
	LUT2 #(
		.INIT('h8)
	) name234 (
		_w110_,
		_w78_,
		_w268_
	);
	LUT4 #(
		.INIT('h0777)
	) name235 (
		_w110_,
		_w78_,
		_w93_,
		_w176_,
		_w269_
	);
	LUT2 #(
		.INIT('h8)
	) name236 (
		_w55_,
		_w176_,
		_w270_
	);
	LUT2 #(
		.INIT('h8)
	) name237 (
		_w59_,
		_w176_,
		_w271_
	);
	LUT3 #(
		.INIT('h1f)
	) name238 (
		_w55_,
		_w59_,
		_w176_,
		_w272_
	);
	LUT2 #(
		.INIT('h8)
	) name239 (
		_w46_,
		_w176_,
		_w273_
	);
	LUT3 #(
		.INIT('h1f)
	) name240 (
		_w110_,
		_w46_,
		_w176_,
		_w274_
	);
	LUT2 #(
		.INIT('h8)
	) name241 (
		_w90_,
		_w176_,
		_w275_
	);
	LUT2 #(
		.INIT('h8)
	) name242 (
		_w78_,
		_w65_,
		_w276_
	);
	LUT4 #(
		.INIT('h135f)
	) name243 (
		_w78_,
		_w90_,
		_w65_,
		_w176_,
		_w277_
	);
	LUT4 #(
		.INIT('h8000)
	) name244 (
		_w274_,
		_w277_,
		_w269_,
		_w272_,
		_w278_
	);
	LUT2 #(
		.INIT('h8)
	) name245 (
		_w266_,
		_w278_,
		_w279_
	);
	LUT4 #(
		.INIT('h0777)
	) name246 (
		_w106_,
		_w59_,
		_w39_,
		_w44_,
		_w280_
	);
	LUT4 #(
		.INIT('h135f)
	) name247 (
		_w122_,
		_w52_,
		_w90_,
		_w39_,
		_w281_
	);
	LUT2 #(
		.INIT('h8)
	) name248 (
		_w67_,
		_w176_,
		_w282_
	);
	LUT4 #(
		.INIT('h0777)
	) name249 (
		_w122_,
		_w52_,
		_w67_,
		_w176_,
		_w283_
	);
	LUT4 #(
		.INIT('h8000)
	) name250 (
		_w66_,
		_w281_,
		_w283_,
		_w280_,
		_w284_
	);
	LUT2 #(
		.INIT('h8)
	) name251 (
		_w78_,
		_w47_,
		_w285_
	);
	LUT2 #(
		.INIT('h8)
	) name252 (
		_w44_,
		_w176_,
		_w286_
	);
	LUT3 #(
		.INIT('h1f)
	) name253 (
		_w50_,
		_w44_,
		_w176_,
		_w287_
	);
	LUT2 #(
		.INIT('h8)
	) name254 (
		_w55_,
		_w236_,
		_w288_
	);
	LUT3 #(
		.INIT('h1f)
	) name255 (
		_w38_,
		_w59_,
		_w43_,
		_w289_
	);
	LUT4 #(
		.INIT('h0400)
	) name256 (
		_w285_,
		_w287_,
		_w288_,
		_w289_,
		_w290_
	);
	LUT2 #(
		.INIT('h8)
	) name257 (
		_w38_,
		_w236_,
		_w291_
	);
	LUT4 #(
		.INIT('h153f)
	) name258 (
		_w38_,
		_w43_,
		_w46_,
		_w236_,
		_w292_
	);
	LUT2 #(
		.INIT('h8)
	) name259 (
		_w54_,
		_w292_,
		_w293_
	);
	LUT2 #(
		.INIT('h8)
	) name260 (
		_w52_,
		_w236_,
		_w294_
	);
	LUT2 #(
		.INIT('h8)
	) name261 (
		_w59_,
		_w236_,
		_w295_
	);
	LUT3 #(
		.INIT('h1f)
	) name262 (
		_w59_,
		_w90_,
		_w236_,
		_w296_
	);
	LUT4 #(
		.INIT('h01ff)
	) name263 (
		_w52_,
		_w59_,
		_w90_,
		_w236_,
		_w297_
	);
	LUT2 #(
		.INIT('h8)
	) name264 (
		_w85_,
		_w236_,
		_w298_
	);
	LUT3 #(
		.INIT('h08)
	) name265 (
		_w58_,
		_w297_,
		_w298_,
		_w299_
	);
	LUT4 #(
		.INIT('h8000)
	) name266 (
		_w293_,
		_w284_,
		_w290_,
		_w299_,
		_w300_
	);
	LUT2 #(
		.INIT('h8)
	) name267 (
		_w44_,
		_w158_,
		_w301_
	);
	LUT3 #(
		.INIT('h1f)
	) name268 (
		_w93_,
		_w44_,
		_w158_,
		_w302_
	);
	LUT2 #(
		.INIT('h8)
	) name269 (
		_w50_,
		_w158_,
		_w303_
	);
	LUT2 #(
		.INIT('h8)
	) name270 (
		_w46_,
		_w158_,
		_w304_
	);
	LUT3 #(
		.INIT('h1f)
	) name271 (
		_w50_,
		_w46_,
		_w158_,
		_w305_
	);
	LUT2 #(
		.INIT('h8)
	) name272 (
		_w302_,
		_w305_,
		_w306_
	);
	LUT3 #(
		.INIT('h80)
	) name273 (
		_w109_,
		_w117_,
		_w306_,
		_w307_
	);
	LUT2 #(
		.INIT('h8)
	) name274 (
		_w67_,
		_w236_,
		_w308_
	);
	LUT3 #(
		.INIT('h57)
	) name275 (
		_w67_,
		_w39_,
		_w236_,
		_w309_
	);
	LUT2 #(
		.INIT('h8)
	) name276 (
		_w56_,
		_w176_,
		_w310_
	);
	LUT4 #(
		.INIT('h0777)
	) name277 (
		_w122_,
		_w55_,
		_w56_,
		_w176_,
		_w311_
	);
	LUT4 #(
		.INIT('h0777)
	) name278 (
		_w38_,
		_w106_,
		_w41_,
		_w43_,
		_w312_
	);
	LUT3 #(
		.INIT('h80)
	) name279 (
		_w311_,
		_w312_,
		_w309_,
		_w313_
	);
	LUT2 #(
		.INIT('h8)
	) name280 (
		_w41_,
		_w259_,
		_w314_
	);
	LUT2 #(
		.INIT('h8)
	) name281 (
		_w44_,
		_w236_,
		_w315_
	);
	LUT4 #(
		.INIT('h153f)
	) name282 (
		_w41_,
		_w44_,
		_w236_,
		_w259_,
		_w316_
	);
	LUT2 #(
		.INIT('h8)
	) name283 (
		_w47_,
		_w176_,
		_w317_
	);
	LUT4 #(
		.INIT('h0777)
	) name284 (
		_w122_,
		_w59_,
		_w47_,
		_w176_,
		_w318_
	);
	LUT3 #(
		.INIT('h80)
	) name285 (
		_w131_,
		_w316_,
		_w318_,
		_w319_
	);
	LUT2 #(
		.INIT('h8)
	) name286 (
		_w41_,
		_w158_,
		_w320_
	);
	LUT2 #(
		.INIT('h8)
	) name287 (
		_w93_,
		_w166_,
		_w321_
	);
	LUT4 #(
		.INIT('h153f)
	) name288 (
		_w41_,
		_w93_,
		_w166_,
		_w158_,
		_w322_
	);
	LUT2 #(
		.INIT('h8)
	) name289 (
		_w41_,
		_w166_,
		_w323_
	);
	LUT2 #(
		.INIT('h8)
	) name290 (
		_w90_,
		_w158_,
		_w324_
	);
	LUT2 #(
		.INIT('h8)
	) name291 (
		_w56_,
		_w158_,
		_w325_
	);
	LUT3 #(
		.INIT('h1f)
	) name292 (
		_w90_,
		_w56_,
		_w158_,
		_w326_
	);
	LUT3 #(
		.INIT('h20)
	) name293 (
		_w322_,
		_w323_,
		_w326_,
		_w327_
	);
	LUT4 #(
		.INIT('h8000)
	) name294 (
		_w49_,
		_w327_,
		_w313_,
		_w319_,
		_w328_
	);
	LUT4 #(
		.INIT('h8000)
	) name295 (
		_w307_,
		_w328_,
		_w279_,
		_w300_,
		_w329_
	);
	LUT3 #(
		.INIT('h80)
	) name296 (
		_w257_,
		_w179_,
		_w329_,
		_w330_
	);
	LUT2 #(
		.INIT('h4)
	) name297 (
		_w157_,
		_w330_,
		_w331_
	);
	LUT2 #(
		.INIT('h2)
	) name298 (
		_w157_,
		_w330_,
		_w332_
	);
	LUT2 #(
		.INIT('h9)
	) name299 (
		_w157_,
		_w330_,
		_w333_
	);
	LUT2 #(
		.INIT('h8)
	) name300 (
		_w55_,
		_w259_,
		_w334_
	);
	LUT2 #(
		.INIT('h8)
	) name301 (
		_w90_,
		_w259_,
		_w335_
	);
	LUT3 #(
		.INIT('h1f)
	) name302 (
		_w90_,
		_w44_,
		_w259_,
		_w336_
	);
	LUT2 #(
		.INIT('h8)
	) name303 (
		_w59_,
		_w259_,
		_w337_
	);
	LUT2 #(
		.INIT('h8)
	) name304 (
		_w85_,
		_w259_,
		_w338_
	);
	LUT2 #(
		.INIT('h8)
	) name305 (
		_w52_,
		_w259_,
		_w339_
	);
	LUT4 #(
		.INIT('h01ff)
	) name306 (
		_w85_,
		_w52_,
		_w59_,
		_w259_,
		_w340_
	);
	LUT3 #(
		.INIT('h40)
	) name307 (
		_w334_,
		_w336_,
		_w340_,
		_w341_
	);
	LUT3 #(
		.INIT('h1f)
	) name308 (
		_w67_,
		_w47_,
		_w176_,
		_w342_
	);
	LUT4 #(
		.INIT('h0777)
	) name309 (
		_w78_,
		_w90_,
		_w41_,
		_w259_,
		_w343_
	);
	LUT3 #(
		.INIT('h1f)
	) name310 (
		_w85_,
		_w56_,
		_w176_,
		_w344_
	);
	LUT3 #(
		.INIT('h80)
	) name311 (
		_w343_,
		_w344_,
		_w342_,
		_w345_
	);
	LUT2 #(
		.INIT('h8)
	) name312 (
		_w93_,
		_w259_,
		_w346_
	);
	LUT2 #(
		.INIT('h8)
	) name313 (
		_w50_,
		_w259_,
		_w347_
	);
	LUT3 #(
		.INIT('h1f)
	) name314 (
		_w50_,
		_w93_,
		_w259_,
		_w348_
	);
	LUT4 #(
		.INIT('h2000)
	) name315 (
		_w150_,
		_w285_,
		_w287_,
		_w348_,
		_w349_
	);
	LUT3 #(
		.INIT('h80)
	) name316 (
		_w140_,
		_w345_,
		_w349_,
		_w350_
	);
	LUT3 #(
		.INIT('h40)
	) name317 (
		_w152_,
		_w279_,
		_w350_,
		_w351_
	);
	LUT4 #(
		.INIT('h4000)
	) name318 (
		_w152_,
		_w279_,
		_w341_,
		_w350_,
		_w352_
	);
	LUT2 #(
		.INIT('h8)
	) name319 (
		_w122_,
		_w93_,
		_w353_
	);
	LUT2 #(
		.INIT('h8)
	) name320 (
		_w122_,
		_w44_,
		_w354_
	);
	LUT2 #(
		.INIT('h8)
	) name321 (
		_w122_,
		_w50_,
		_w355_
	);
	LUT3 #(
		.INIT('h57)
	) name322 (
		_w122_,
		_w50_,
		_w44_,
		_w356_
	);
	LUT4 #(
		.INIT('h5557)
	) name323 (
		_w122_,
		_w50_,
		_w93_,
		_w44_,
		_w357_
	);
	LUT2 #(
		.INIT('h8)
	) name324 (
		_w122_,
		_w56_,
		_w358_
	);
	LUT2 #(
		.INIT('h8)
	) name325 (
		_w38_,
		_w259_,
		_w359_
	);
	LUT2 #(
		.INIT('h8)
	) name326 (
		_w122_,
		_w46_,
		_w360_
	);
	LUT4 #(
		.INIT('h153f)
	) name327 (
		_w38_,
		_w122_,
		_w46_,
		_w259_,
		_w361_
	);
	LUT2 #(
		.INIT('h8)
	) name328 (
		_w110_,
		_w259_,
		_w362_
	);
	LUT2 #(
		.INIT('h8)
	) name329 (
		_w67_,
		_w259_,
		_w363_
	);
	LUT3 #(
		.INIT('h1f)
	) name330 (
		_w110_,
		_w67_,
		_w259_,
		_w364_
	);
	LUT2 #(
		.INIT('h8)
	) name331 (
		_w47_,
		_w259_,
		_w365_
	);
	LUT2 #(
		.INIT('h8)
	) name332 (
		_w65_,
		_w259_,
		_w366_
	);
	LUT3 #(
		.INIT('h1f)
	) name333 (
		_w47_,
		_w65_,
		_w259_,
		_w367_
	);
	LUT4 #(
		.INIT('h4000)
	) name334 (
		_w358_,
		_w361_,
		_w364_,
		_w367_,
		_w368_
	);
	LUT2 #(
		.INIT('h8)
	) name335 (
		_w122_,
		_w41_,
		_w369_
	);
	LUT3 #(
		.INIT('h37)
	) name336 (
		_w38_,
		_w122_,
		_w41_,
		_w370_
	);
	LUT4 #(
		.INIT('h3337)
	) name337 (
		_w38_,
		_w122_,
		_w41_,
		_w65_,
		_w371_
	);
	LUT4 #(
		.INIT('h8000)
	) name338 (
		_w123_,
		_w126_,
		_w149_,
		_w371_,
		_w372_
	);
	LUT3 #(
		.INIT('h80)
	) name339 (
		_w357_,
		_w368_,
		_w372_,
		_w373_
	);
	LUT2 #(
		.INIT('h8)
	) name340 (
		_w352_,
		_w373_,
		_w374_
	);
	LUT2 #(
		.INIT('h9)
	) name341 (
		\a[29] ,
		\a[30] ,
		_w375_
	);
	LUT3 #(
		.INIT('h80)
	) name342 (
		\a[29] ,
		\a[30] ,
		\a[31] ,
		_w376_
	);
	LUT3 #(
		.INIT('h60)
	) name343 (
		\a[29] ,
		\a[30] ,
		\a[31] ,
		_w377_
	);
	LUT4 #(
		.INIT('h0100)
	) name344 (
		\a[27] ,
		\a[28] ,
		\a[29] ,
		\a[30] ,
		_w378_
	);
	LUT2 #(
		.INIT('h8)
	) name345 (
		_w67_,
		_w378_,
		_w379_
	);
	LUT2 #(
		.INIT('h8)
	) name346 (
		_w38_,
		_w378_,
		_w380_
	);
	LUT3 #(
		.INIT('h1f)
	) name347 (
		_w38_,
		_w67_,
		_w378_,
		_w381_
	);
	LUT2 #(
		.INIT('h8)
	) name348 (
		_w52_,
		_w378_,
		_w382_
	);
	LUT2 #(
		.INIT('h8)
	) name349 (
		_w47_,
		_w378_,
		_w383_
	);
	LUT3 #(
		.INIT('h1f)
	) name350 (
		_w52_,
		_w47_,
		_w378_,
		_w384_
	);
	LUT2 #(
		.INIT('h8)
	) name351 (
		_w59_,
		_w378_,
		_w385_
	);
	LUT2 #(
		.INIT('h8)
	) name352 (
		_w41_,
		_w378_,
		_w386_
	);
	LUT3 #(
		.INIT('h1f)
	) name353 (
		_w59_,
		_w41_,
		_w378_,
		_w387_
	);
	LUT3 #(
		.INIT('h80)
	) name354 (
		_w384_,
		_w387_,
		_w381_,
		_w388_
	);
	LUT2 #(
		.INIT('h8)
	) name355 (
		_w50_,
		_w378_,
		_w389_
	);
	LUT2 #(
		.INIT('h8)
	) name356 (
		_w46_,
		_w378_,
		_w390_
	);
	LUT3 #(
		.INIT('h1f)
	) name357 (
		_w50_,
		_w46_,
		_w378_,
		_w391_
	);
	LUT2 #(
		.INIT('h8)
	) name358 (
		_w110_,
		_w378_,
		_w392_
	);
	LUT2 #(
		.INIT('h8)
	) name359 (
		_w85_,
		_w378_,
		_w393_
	);
	LUT3 #(
		.INIT('h1f)
	) name360 (
		_w85_,
		_w110_,
		_w378_,
		_w394_
	);
	LUT2 #(
		.INIT('h8)
	) name361 (
		_w391_,
		_w394_,
		_w395_
	);
	LUT2 #(
		.INIT('h8)
	) name362 (
		_w55_,
		_w378_,
		_w396_
	);
	LUT2 #(
		.INIT('h8)
	) name363 (
		_w65_,
		_w378_,
		_w397_
	);
	LUT2 #(
		.INIT('h8)
	) name364 (
		_w56_,
		_w378_,
		_w398_
	);
	LUT4 #(
		.INIT('h01ff)
	) name365 (
		_w55_,
		_w56_,
		_w65_,
		_w378_,
		_w399_
	);
	LUT2 #(
		.INIT('h8)
	) name366 (
		_w106_,
		_w46_,
		_w400_
	);
	LUT4 #(
		.INIT('h135f)
	) name367 (
		_w106_,
		_w44_,
		_w46_,
		_w378_,
		_w401_
	);
	LUT2 #(
		.INIT('h8)
	) name368 (
		_w93_,
		_w378_,
		_w402_
	);
	LUT3 #(
		.INIT('h1f)
	) name369 (
		_w90_,
		_w93_,
		_w378_,
		_w403_
	);
	LUT3 #(
		.INIT('h80)
	) name370 (
		_w401_,
		_w403_,
		_w399_,
		_w404_
	);
	LUT3 #(
		.INIT('h80)
	) name371 (
		_w395_,
		_w388_,
		_w404_,
		_w405_
	);
	LUT2 #(
		.INIT('h8)
	) name372 (
		_w106_,
		_w93_,
		_w406_
	);
	LUT2 #(
		.INIT('h8)
	) name373 (
		_w106_,
		_w41_,
		_w407_
	);
	LUT3 #(
		.INIT('h57)
	) name374 (
		_w106_,
		_w41_,
		_w93_,
		_w408_
	);
	LUT2 #(
		.INIT('h8)
	) name375 (
		_w106_,
		_w44_,
		_w409_
	);
	LUT2 #(
		.INIT('h8)
	) name376 (
		_w106_,
		_w56_,
		_w410_
	);
	LUT3 #(
		.INIT('h57)
	) name377 (
		_w106_,
		_w56_,
		_w44_,
		_w411_
	);
	LUT2 #(
		.INIT('h8)
	) name378 (
		_w106_,
		_w90_,
		_w412_
	);
	LUT2 #(
		.INIT('h8)
	) name379 (
		_w106_,
		_w50_,
		_w413_
	);
	LUT3 #(
		.INIT('h57)
	) name380 (
		_w106_,
		_w90_,
		_w50_,
		_w414_
	);
	LUT3 #(
		.INIT('h80)
	) name381 (
		_w408_,
		_w411_,
		_w414_,
		_w415_
	);
	LUT4 #(
		.INIT('h8000)
	) name382 (
		_w395_,
		_w388_,
		_w404_,
		_w415_,
		_w416_
	);
	LUT3 #(
		.INIT('h80)
	) name383 (
		_w131_,
		_w132_,
		_w144_,
		_w417_
	);
	LUT2 #(
		.INIT('h8)
	) name384 (
		_w416_,
		_w417_,
		_w418_
	);
	LUT4 #(
		.INIT('h0200)
	) name385 (
		\a[27] ,
		\a[28] ,
		\a[29] ,
		\a[30] ,
		_w419_
	);
	LUT2 #(
		.INIT('h8)
	) name386 (
		_w65_,
		_w419_,
		_w420_
	);
	LUT4 #(
		.INIT('h135f)
	) name387 (
		_w55_,
		_w65_,
		_w259_,
		_w419_,
		_w421_
	);
	LUT4 #(
		.INIT('h8000)
	) name388 (
		_w357_,
		_w368_,
		_w372_,
		_w421_,
		_w422_
	);
	LUT3 #(
		.INIT('h80)
	) name389 (
		_w121_,
		_w418_,
		_w422_,
		_w423_
	);
	LUT2 #(
		.INIT('h8)
	) name390 (
		_w59_,
		_w419_,
		_w424_
	);
	LUT2 #(
		.INIT('h8)
	) name391 (
		_w46_,
		_w419_,
		_w425_
	);
	LUT2 #(
		.INIT('h8)
	) name392 (
		_w93_,
		_w419_,
		_w426_
	);
	LUT3 #(
		.INIT('h1f)
	) name393 (
		_w93_,
		_w46_,
		_w419_,
		_w427_
	);
	LUT4 #(
		.INIT('h01ff)
	) name394 (
		_w59_,
		_w93_,
		_w46_,
		_w419_,
		_w428_
	);
	LUT2 #(
		.INIT('h8)
	) name395 (
		_w44_,
		_w419_,
		_w429_
	);
	LUT4 #(
		.INIT('h0400)
	) name396 (
		\a[27] ,
		\a[28] ,
		\a[29] ,
		\a[30] ,
		_w430_
	);
	LUT2 #(
		.INIT('h8)
	) name397 (
		_w47_,
		_w430_,
		_w431_
	);
	LUT2 #(
		.INIT('h8)
	) name398 (
		_w50_,
		_w419_,
		_w432_
	);
	LUT4 #(
		.INIT('h153f)
	) name399 (
		_w47_,
		_w50_,
		_w419_,
		_w430_,
		_w433_
	);
	LUT3 #(
		.INIT('h20)
	) name400 (
		_w428_,
		_w429_,
		_w433_,
		_w434_
	);
	LUT2 #(
		.INIT('h8)
	) name401 (
		_w56_,
		_w419_,
		_w435_
	);
	LUT2 #(
		.INIT('h8)
	) name402 (
		_w38_,
		_w419_,
		_w436_
	);
	LUT2 #(
		.INIT('h8)
	) name403 (
		_w67_,
		_w419_,
		_w437_
	);
	LUT4 #(
		.INIT('h01ff)
	) name404 (
		_w38_,
		_w67_,
		_w56_,
		_w419_,
		_w438_
	);
	LUT2 #(
		.INIT('h8)
	) name405 (
		_w85_,
		_w419_,
		_w439_
	);
	LUT2 #(
		.INIT('h8)
	) name406 (
		_w41_,
		_w419_,
		_w440_
	);
	LUT2 #(
		.INIT('h8)
	) name407 (
		_w65_,
		_w430_,
		_w441_
	);
	LUT4 #(
		.INIT('h135f)
	) name408 (
		_w41_,
		_w65_,
		_w419_,
		_w430_,
		_w442_
	);
	LUT2 #(
		.INIT('h8)
	) name409 (
		_w90_,
		_w419_,
		_w443_
	);
	LUT2 #(
		.INIT('h8)
	) name410 (
		_w55_,
		_w419_,
		_w444_
	);
	LUT2 #(
		.INIT('h8)
	) name411 (
		_w52_,
		_w419_,
		_w445_
	);
	LUT3 #(
		.INIT('h1f)
	) name412 (
		_w55_,
		_w52_,
		_w419_,
		_w446_
	);
	LUT4 #(
		.INIT('h01ff)
	) name413 (
		_w55_,
		_w52_,
		_w90_,
		_w419_,
		_w447_
	);
	LUT4 #(
		.INIT('h4000)
	) name414 (
		_w439_,
		_w442_,
		_w447_,
		_w438_,
		_w448_
	);
	LUT2 #(
		.INIT('h8)
	) name415 (
		_w434_,
		_w448_,
		_w449_
	);
	LUT2 #(
		.INIT('h8)
	) name416 (
		_w56_,
		_w430_,
		_w450_
	);
	LUT2 #(
		.INIT('h8)
	) name417 (
		_w55_,
		_w430_,
		_w451_
	);
	LUT2 #(
		.INIT('h8)
	) name418 (
		_w59_,
		_w430_,
		_w452_
	);
	LUT4 #(
		.INIT('h01ff)
	) name419 (
		_w55_,
		_w59_,
		_w56_,
		_w430_,
		_w453_
	);
	LUT2 #(
		.INIT('h8)
	) name420 (
		_w50_,
		_w430_,
		_w454_
	);
	LUT2 #(
		.INIT('h8)
	) name421 (
		_w52_,
		_w430_,
		_w455_
	);
	LUT3 #(
		.INIT('h1f)
	) name422 (
		_w52_,
		_w50_,
		_w430_,
		_w456_
	);
	LUT2 #(
		.INIT('h8)
	) name423 (
		_w47_,
		_w236_,
		_w457_
	);
	LUT2 #(
		.INIT('h8)
	) name424 (
		_w41_,
		_w430_,
		_w458_
	);
	LUT4 #(
		.INIT('h135f)
	) name425 (
		_w47_,
		_w41_,
		_w236_,
		_w430_,
		_w459_
	);
	LUT3 #(
		.INIT('h80)
	) name426 (
		_w456_,
		_w459_,
		_w453_,
		_w460_
	);
	LUT2 #(
		.INIT('h8)
	) name427 (
		_w93_,
		_w430_,
		_w461_
	);
	LUT2 #(
		.INIT('h8)
	) name428 (
		_w46_,
		_w430_,
		_w462_
	);
	LUT2 #(
		.INIT('h8)
	) name429 (
		_w44_,
		_w430_,
		_w463_
	);
	LUT3 #(
		.INIT('h1f)
	) name430 (
		_w44_,
		_w46_,
		_w430_,
		_w464_
	);
	LUT4 #(
		.INIT('h01ff)
	) name431 (
		_w93_,
		_w44_,
		_w46_,
		_w430_,
		_w465_
	);
	LUT4 #(
		.INIT('h8000)
	) name432 (
		_w456_,
		_w459_,
		_w453_,
		_w465_,
		_w466_
	);
	LUT2 #(
		.INIT('h2)
	) name433 (
		_w297_,
		_w288_,
		_w467_
	);
	LUT2 #(
		.INIT('h8)
	) name434 (
		_w67_,
		_w430_,
		_w468_
	);
	LUT2 #(
		.INIT('h8)
	) name435 (
		_w38_,
		_w430_,
		_w469_
	);
	LUT3 #(
		.INIT('h1f)
	) name436 (
		_w38_,
		_w67_,
		_w430_,
		_w470_
	);
	LUT2 #(
		.INIT('h8)
	) name437 (
		_w110_,
		_w430_,
		_w471_
	);
	LUT4 #(
		.INIT('h135f)
	) name438 (
		_w85_,
		_w110_,
		_w236_,
		_w430_,
		_w472_
	);
	LUT2 #(
		.INIT('h8)
	) name439 (
		_w110_,
		_w419_,
		_w473_
	);
	LUT4 #(
		.INIT('h153f)
	) name440 (
		_w110_,
		_w44_,
		_w236_,
		_w419_,
		_w474_
	);
	LUT3 #(
		.INIT('h80)
	) name441 (
		_w472_,
		_w474_,
		_w470_,
		_w475_
	);
	LUT2 #(
		.INIT('h8)
	) name442 (
		_w65_,
		_w236_,
		_w476_
	);
	LUT2 #(
		.INIT('h8)
	) name443 (
		_w90_,
		_w430_,
		_w477_
	);
	LUT2 #(
		.INIT('h8)
	) name444 (
		_w47_,
		_w419_,
		_w478_
	);
	LUT4 #(
		.INIT('h153f)
	) name445 (
		_w90_,
		_w47_,
		_w419_,
		_w430_,
		_w479_
	);
	LUT3 #(
		.INIT('h1f)
	) name446 (
		_w38_,
		_w67_,
		_w236_,
		_w480_
	);
	LUT2 #(
		.INIT('h8)
	) name447 (
		_w110_,
		_w236_,
		_w481_
	);
	LUT2 #(
		.INIT('h8)
	) name448 (
		_w85_,
		_w430_,
		_w482_
	);
	LUT4 #(
		.INIT('h153f)
	) name449 (
		_w85_,
		_w110_,
		_w236_,
		_w430_,
		_w483_
	);
	LUT4 #(
		.INIT('h4000)
	) name450 (
		_w476_,
		_w479_,
		_w480_,
		_w483_,
		_w484_
	);
	LUT4 #(
		.INIT('h8000)
	) name451 (
		_w466_,
		_w467_,
		_w475_,
		_w484_,
		_w485_
	);
	LUT2 #(
		.INIT('h8)
	) name452 (
		_w449_,
		_w485_,
		_w486_
	);
	LUT4 #(
		.INIT('h8000)
	) name453 (
		_w234_,
		_w200_,
		_w256_,
		_w175_,
		_w487_
	);
	LUT3 #(
		.INIT('h37)
	) name454 (
		_w67_,
		_w43_,
		_w65_,
		_w488_
	);
	LUT2 #(
		.INIT('h4)
	) name455 (
		_w317_,
		_w488_,
		_w489_
	);
	LUT3 #(
		.INIT('h1f)
	) name456 (
		_w38_,
		_w110_,
		_w43_,
		_w490_
	);
	LUT4 #(
		.INIT('h153f)
	) name457 (
		_w110_,
		_w47_,
		_w43_,
		_w176_,
		_w491_
	);
	LUT3 #(
		.INIT('h57)
	) name458 (
		_w41_,
		_w72_,
		_w259_,
		_w492_
	);
	LUT4 #(
		.INIT('h8000)
	) name459 (
		_w262_,
		_w490_,
		_w491_,
		_w492_,
		_w493_
	);
	LUT2 #(
		.INIT('h4)
	) name460 (
		_w264_,
		_w348_,
		_w494_
	);
	LUT4 #(
		.INIT('h135f)
	) name461 (
		_w110_,
		_w56_,
		_w72_,
		_w259_,
		_w495_
	);
	LUT4 #(
		.INIT('h153f)
	) name462 (
		_w55_,
		_w72_,
		_w44_,
		_w176_,
		_w496_
	);
	LUT3 #(
		.INIT('h1f)
	) name463 (
		_w38_,
		_w67_,
		_w176_,
		_w497_
	);
	LUT3 #(
		.INIT('h80)
	) name464 (
		_w496_,
		_w497_,
		_w495_,
		_w498_
	);
	LUT4 #(
		.INIT('h8000)
	) name465 (
		_w489_,
		_w493_,
		_w494_,
		_w498_,
		_w499_
	);
	LUT2 #(
		.INIT('h2)
	) name466 (
		_w123_,
		_w60_,
		_w500_
	);
	LUT4 #(
		.INIT('h135f)
	) name467 (
		_w52_,
		_w41_,
		_w43_,
		_w166_,
		_w501_
	);
	LUT3 #(
		.INIT('h1f)
	) name468 (
		_w56_,
		_w50_,
		_w43_,
		_w502_
	);
	LUT4 #(
		.INIT('h135f)
	) name469 (
		_w43_,
		_w93_,
		_w44_,
		_w166_,
		_w503_
	);
	LUT4 #(
		.INIT('h8000)
	) name470 (
		_w105_,
		_w503_,
		_w501_,
		_w502_,
		_w504_
	);
	LUT2 #(
		.INIT('h8)
	) name471 (
		_w500_,
		_w504_,
		_w505_
	);
	LUT4 #(
		.INIT('h131f)
	) name472 (
		_w55_,
		_w85_,
		_w43_,
		_w176_,
		_w506_
	);
	LUT3 #(
		.INIT('h80)
	) name473 (
		_w336_,
		_w340_,
		_w506_,
		_w507_
	);
	LUT3 #(
		.INIT('h80)
	) name474 (
		_w500_,
		_w504_,
		_w507_,
		_w508_
	);
	LUT3 #(
		.INIT('h80)
	) name475 (
		_w100_,
		_w499_,
		_w508_,
		_w509_
	);
	LUT3 #(
		.INIT('h80)
	) name476 (
		_w486_,
		_w487_,
		_w509_,
		_w510_
	);
	LUT2 #(
		.INIT('h1)
	) name477 (
		_w423_,
		_w510_,
		_w511_
	);
	LUT4 #(
		.INIT('h153f)
	) name478 (
		_w110_,
		_w41_,
		_w176_,
		_w430_,
		_w512_
	);
	LUT4 #(
		.INIT('h135f)
	) name479 (
		_w59_,
		_w78_,
		_w39_,
		_w65_,
		_w513_
	);
	LUT4 #(
		.INIT('h153f)
	) name480 (
		_w38_,
		_w59_,
		_w259_,
		_w430_,
		_w514_
	);
	LUT3 #(
		.INIT('h80)
	) name481 (
		_w513_,
		_w514_,
		_w512_,
		_w515_
	);
	LUT3 #(
		.INIT('h1f)
	) name482 (
		_w52_,
		_w67_,
		_w39_,
		_w516_
	);
	LUT4 #(
		.INIT('h135f)
	) name483 (
		_w90_,
		_w56_,
		_w72_,
		_w39_,
		_w517_
	);
	LUT4 #(
		.INIT('h0777)
	) name484 (
		_w38_,
		_w72_,
		_w39_,
		_w50_,
		_w518_
	);
	LUT4 #(
		.INIT('h135f)
	) name485 (
		_w52_,
		_w46_,
		_w259_,
		_w176_,
		_w519_
	);
	LUT4 #(
		.INIT('h8000)
	) name486 (
		_w518_,
		_w519_,
		_w516_,
		_w517_,
		_w520_
	);
	LUT3 #(
		.INIT('h57)
	) name487 (
		_w72_,
		_w93_,
		_w44_,
		_w521_
	);
	LUT4 #(
		.INIT('h135f)
	) name488 (
		_w85_,
		_w72_,
		_w39_,
		_w50_,
		_w522_
	);
	LUT4 #(
		.INIT('h135f)
	) name489 (
		_w41_,
		_w44_,
		_w158_,
		_w176_,
		_w523_
	);
	LUT3 #(
		.INIT('h1f)
	) name490 (
		_w110_,
		_w65_,
		_w236_,
		_w524_
	);
	LUT4 #(
		.INIT('h8000)
	) name491 (
		_w521_,
		_w522_,
		_w523_,
		_w524_,
		_w525_
	);
	LUT3 #(
		.INIT('h80)
	) name492 (
		_w515_,
		_w520_,
		_w525_,
		_w526_
	);
	LUT4 #(
		.INIT('h0777)
	) name493 (
		_w59_,
		_w72_,
		_w93_,
		_w176_,
		_w527_
	);
	LUT4 #(
		.INIT('h135f)
	) name494 (
		_w85_,
		_w59_,
		_w259_,
		_w176_,
		_w528_
	);
	LUT3 #(
		.INIT('h40)
	) name495 (
		_w482_,
		_w527_,
		_w528_,
		_w529_
	);
	LUT4 #(
		.INIT('h153f)
	) name496 (
		_w52_,
		_w78_,
		_w47_,
		_w72_,
		_w530_
	);
	LUT4 #(
		.INIT('h153f)
	) name497 (
		_w67_,
		_w44_,
		_w259_,
		_w430_,
		_w531_
	);
	LUT3 #(
		.INIT('h80)
	) name498 (
		_w87_,
		_w530_,
		_w531_,
		_w532_
	);
	LUT4 #(
		.INIT('h135f)
	) name499 (
		_w39_,
		_w50_,
		_w93_,
		_w176_,
		_w533_
	);
	LUT4 #(
		.INIT('h135f)
	) name500 (
		_w110_,
		_w56_,
		_w72_,
		_w176_,
		_w534_
	);
	LUT4 #(
		.INIT('h153f)
	) name501 (
		_w90_,
		_w39_,
		_w44_,
		_w430_,
		_w535_
	);
	LUT4 #(
		.INIT('h8000)
	) name502 (
		_w42_,
		_w533_,
		_w534_,
		_w535_,
		_w536_
	);
	LUT3 #(
		.INIT('h80)
	) name503 (
		_w532_,
		_w529_,
		_w536_,
		_w537_
	);
	LUT3 #(
		.INIT('h57)
	) name504 (
		_w90_,
		_w158_,
		_w176_,
		_w538_
	);
	LUT3 #(
		.INIT('h1f)
	) name505 (
		_w55_,
		_w90_,
		_w39_,
		_w539_
	);
	LUT2 #(
		.INIT('h8)
	) name506 (
		_w538_,
		_w539_,
		_w540_
	);
	LUT4 #(
		.INIT('h135f)
	) name507 (
		_w67_,
		_w56_,
		_w72_,
		_w158_,
		_w541_
	);
	LUT4 #(
		.INIT('h0800)
	) name508 (
		_w302_,
		_w305_,
		_w335_,
		_w541_,
		_w542_
	);
	LUT3 #(
		.INIT('h80)
	) name509 (
		_w466_,
		_w540_,
		_w542_,
		_w543_
	);
	LUT3 #(
		.INIT('h80)
	) name510 (
		_w526_,
		_w537_,
		_w543_,
		_w544_
	);
	LUT4 #(
		.INIT('h135f)
	) name511 (
		_w122_,
		_w106_,
		_w90_,
		_w65_,
		_w545_
	);
	LUT4 #(
		.INIT('h0777)
	) name512 (
		_w122_,
		_w56_,
		_w39_,
		_w46_,
		_w546_
	);
	LUT4 #(
		.INIT('h8000)
	) name513 (
		_w89_,
		_w357_,
		_w545_,
		_w546_,
		_w547_
	);
	LUT2 #(
		.INIT('h8)
	) name514 (
		_w467_,
		_w547_,
		_w548_
	);
	LUT2 #(
		.INIT('h4)
	) name515 (
		_w79_,
		_w348_,
		_w549_
	);
	LUT4 #(
		.INIT('h0777)
	) name516 (
		_w122_,
		_w59_,
		_w41_,
		_w43_,
		_w550_
	);
	LUT4 #(
		.INIT('h153f)
	) name517 (
		_w56_,
		_w47_,
		_w72_,
		_w259_,
		_w551_
	);
	LUT4 #(
		.INIT('h4000)
	) name518 (
		_w64_,
		_w66_,
		_w550_,
		_w551_,
		_w552_
	);
	LUT3 #(
		.INIT('h1f)
	) name519 (
		_w110_,
		_w47_,
		_w419_,
		_w553_
	);
	LUT3 #(
		.INIT('h57)
	) name520 (
		_w122_,
		_w47_,
		_w41_,
		_w554_
	);
	LUT4 #(
		.INIT('h153f)
	) name521 (
		_w85_,
		_w110_,
		_w39_,
		_w236_,
		_w555_
	);
	LUT4 #(
		.INIT('h8000)
	) name522 (
		_w480_,
		_w553_,
		_w554_,
		_w555_,
		_w556_
	);
	LUT4 #(
		.INIT('h8000)
	) name523 (
		_w145_,
		_w549_,
		_w556_,
		_w552_,
		_w557_
	);
	LUT3 #(
		.INIT('h80)
	) name524 (
		_w449_,
		_w548_,
		_w557_,
		_w558_
	);
	LUT2 #(
		.INIT('h8)
	) name525 (
		_w544_,
		_w558_,
		_w559_
	);
	LUT4 #(
		.INIT('h135f)
	) name526 (
		_w38_,
		_w46_,
		_w201_,
		_w158_,
		_w560_
	);
	LUT2 #(
		.INIT('h4)
	) name527 (
		_w337_,
		_w560_,
		_w561_
	);
	LUT4 #(
		.INIT('h135f)
	) name528 (
		_w106_,
		_w44_,
		_w46_,
		_w419_,
		_w562_
	);
	LUT4 #(
		.INIT('h153f)
	) name529 (
		_w110_,
		_w67_,
		_w72_,
		_w201_,
		_w563_
	);
	LUT4 #(
		.INIT('h135f)
	) name530 (
		_w106_,
		_w50_,
		_w44_,
		_w201_,
		_w564_
	);
	LUT4 #(
		.INIT('h4000)
	) name531 (
		_w251_,
		_w562_,
		_w563_,
		_w564_,
		_w565_
	);
	LUT4 #(
		.INIT('h153f)
	) name532 (
		_w85_,
		_w50_,
		_w158_,
		_w259_,
		_w566_
	);
	LUT4 #(
		.INIT('h135f)
	) name533 (
		_w106_,
		_w110_,
		_w56_,
		_w430_,
		_w567_
	);
	LUT3 #(
		.INIT('h40)
	) name534 (
		_w426_,
		_w567_,
		_w566_,
		_w568_
	);
	LUT3 #(
		.INIT('h80)
	) name535 (
		_w561_,
		_w565_,
		_w568_,
		_w569_
	);
	LUT4 #(
		.INIT('h113f)
	) name536 (
		_w85_,
		_w90_,
		_w259_,
		_w419_,
		_w570_
	);
	LUT3 #(
		.INIT('h1f)
	) name537 (
		_w52_,
		_w59_,
		_w201_,
		_w571_
	);
	LUT4 #(
		.INIT('h8000)
	) name538 (
		_w130_,
		_w81_,
		_w287_,
		_w571_,
		_w572_
	);
	LUT2 #(
		.INIT('h8)
	) name539 (
		_w570_,
		_w572_,
		_w573_
	);
	LUT4 #(
		.INIT('h153f)
	) name540 (
		_w56_,
		_w44_,
		_w201_,
		_w158_,
		_w574_
	);
	LUT4 #(
		.INIT('h0777)
	) name541 (
		_w122_,
		_w90_,
		_w41_,
		_w236_,
		_w575_
	);
	LUT3 #(
		.INIT('h80)
	) name542 (
		_w438_,
		_w574_,
		_w575_,
		_w576_
	);
	LUT3 #(
		.INIT('h1f)
	) name543 (
		_w93_,
		_w46_,
		_w236_,
		_w577_
	);
	LUT3 #(
		.INIT('h57)
	) name544 (
		_w65_,
		_w378_,
		_w430_,
		_w578_
	);
	LUT3 #(
		.INIT('h37)
	) name545 (
		_w43_,
		_w46_,
		_w201_,
		_w579_
	);
	LUT4 #(
		.INIT('h0777)
	) name546 (
		_w122_,
		_w59_,
		_w65_,
		_w201_,
		_w580_
	);
	LUT4 #(
		.INIT('h8000)
	) name547 (
		_w579_,
		_w580_,
		_w577_,
		_w578_,
		_w581_
	);
	LUT4 #(
		.INIT('h153f)
	) name548 (
		_w55_,
		_w65_,
		_w184_,
		_w419_,
		_w582_
	);
	LUT4 #(
		.INIT('h135f)
	) name549 (
		_w106_,
		_w41_,
		_w50_,
		_w201_,
		_w583_
	);
	LUT4 #(
		.INIT('h0777)
	) name550 (
		_w106_,
		_w90_,
		_w41_,
		_w43_,
		_w584_
	);
	LUT4 #(
		.INIT('h8000)
	) name551 (
		_w538_,
		_w582_,
		_w583_,
		_w584_,
		_w585_
	);
	LUT3 #(
		.INIT('h80)
	) name552 (
		_w581_,
		_w576_,
		_w585_,
		_w586_
	);
	LUT3 #(
		.INIT('h80)
	) name553 (
		_w569_,
		_w573_,
		_w586_,
		_w587_
	);
	LUT2 #(
		.INIT('h2)
	) name554 (
		_w132_,
		_w432_,
		_w588_
	);
	LUT4 #(
		.INIT('h153f)
	) name555 (
		_w59_,
		_w67_,
		_w201_,
		_w176_,
		_w589_
	);
	LUT4 #(
		.INIT('h153f)
	) name556 (
		_w55_,
		_w110_,
		_w184_,
		_w201_,
		_w590_
	);
	LUT3 #(
		.INIT('h80)
	) name557 (
		_w408_,
		_w589_,
		_w590_,
		_w591_
	);
	LUT2 #(
		.INIT('h8)
	) name558 (
		_w588_,
		_w591_,
		_w592_
	);
	LUT4 #(
		.INIT('h135f)
	) name559 (
		_w56_,
		_w93_,
		_w201_,
		_w176_,
		_w593_
	);
	LUT4 #(
		.INIT('h0777)
	) name560 (
		_w38_,
		_w72_,
		_w46_,
		_w419_,
		_w594_
	);
	LUT4 #(
		.INIT('h0777)
	) name561 (
		_w106_,
		_w52_,
		_w72_,
		_w65_,
		_w595_
	);
	LUT4 #(
		.INIT('h4000)
	) name562 (
		_w431_,
		_w594_,
		_w595_,
		_w593_,
		_w596_
	);
	LUT4 #(
		.INIT('h153f)
	) name563 (
		_w52_,
		_w41_,
		_w158_,
		_w419_,
		_w597_
	);
	LUT4 #(
		.INIT('h135f)
	) name564 (
		_w39_,
		_w93_,
		_w65_,
		_w201_,
		_w598_
	);
	LUT2 #(
		.INIT('h2)
	) name565 (
		_w254_,
		_w440_,
		_w599_
	);
	LUT4 #(
		.INIT('h2000)
	) name566 (
		_w254_,
		_w440_,
		_w597_,
		_w598_,
		_w600_
	);
	LUT4 #(
		.INIT('h035f)
	) name567 (
		_w122_,
		_w93_,
		_w44_,
		_w158_,
		_w601_
	);
	LUT4 #(
		.INIT('h135f)
	) name568 (
		_w110_,
		_w47_,
		_w72_,
		_w39_,
		_w602_
	);
	LUT2 #(
		.INIT('h8)
	) name569 (
		_w601_,
		_w602_,
		_w603_
	);
	LUT4 #(
		.INIT('h135f)
	) name570 (
		_w52_,
		_w59_,
		_w259_,
		_w419_,
		_w604_
	);
	LUT4 #(
		.INIT('h135f)
	) name571 (
		_w78_,
		_w56_,
		_w46_,
		_w236_,
		_w605_
	);
	LUT4 #(
		.INIT('h4000)
	) name572 (
		_w111_,
		_w231_,
		_w604_,
		_w605_,
		_w606_
	);
	LUT4 #(
		.INIT('h8000)
	) name573 (
		_w603_,
		_w606_,
		_w596_,
		_w600_,
		_w607_
	);
	LUT2 #(
		.INIT('h8)
	) name574 (
		_w592_,
		_w607_,
		_w608_
	);
	LUT4 #(
		.INIT('h0777)
	) name575 (
		_w38_,
		_w122_,
		_w47_,
		_w259_,
		_w609_
	);
	LUT4 #(
		.INIT('h153f)
	) name576 (
		_w38_,
		_w85_,
		_w39_,
		_w184_,
		_w610_
	);
	LUT4 #(
		.INIT('h0777)
	) name577 (
		_w56_,
		_w72_,
		_w65_,
		_w259_,
		_w611_
	);
	LUT3 #(
		.INIT('h80)
	) name578 (
		_w610_,
		_w611_,
		_w609_,
		_w612_
	);
	LUT3 #(
		.INIT('h1f)
	) name579 (
		_w85_,
		_w110_,
		_w78_,
		_w613_
	);
	LUT2 #(
		.INIT('h4)
	) name580 (
		_w360_,
		_w613_,
		_w614_
	);
	LUT4 #(
		.INIT('h135f)
	) name581 (
		_w72_,
		_w44_,
		_w46_,
		_w236_,
		_w615_
	);
	LUT4 #(
		.INIT('h8000)
	) name582 (
		_w125_,
		_w150_,
		_w553_,
		_w615_,
		_w616_
	);
	LUT3 #(
		.INIT('h80)
	) name583 (
		_w614_,
		_w612_,
		_w616_,
		_w617_
	);
	LUT4 #(
		.INIT('h01ff)
	) name584 (
		_w55_,
		_w59_,
		_w67_,
		_w39_,
		_w618_
	);
	LUT4 #(
		.INIT('h135f)
	) name585 (
		_w38_,
		_w47_,
		_w39_,
		_w378_,
		_w619_
	);
	LUT4 #(
		.INIT('h135f)
	) name586 (
		_w55_,
		_w52_,
		_w78_,
		_w39_,
		_w620_
	);
	LUT4 #(
		.INIT('h135f)
	) name587 (
		_w52_,
		_w67_,
		_w78_,
		_w184_,
		_w621_
	);
	LUT4 #(
		.INIT('h8000)
	) name588 (
		_w620_,
		_w621_,
		_w619_,
		_w618_,
		_w622_
	);
	LUT3 #(
		.INIT('h80)
	) name589 (
		_w489_,
		_w493_,
		_w622_,
		_w623_
	);
	LUT2 #(
		.INIT('h8)
	) name590 (
		_w617_,
		_w623_,
		_w624_
	);
	LUT3 #(
		.INIT('h80)
	) name591 (
		_w587_,
		_w608_,
		_w624_,
		_w625_
	);
	LUT2 #(
		.INIT('h1)
	) name592 (
		_w559_,
		_w625_,
		_w626_
	);
	LUT4 #(
		.INIT('h153f)
	) name593 (
		_w122_,
		_w106_,
		_w52_,
		_w59_,
		_w627_
	);
	LUT2 #(
		.INIT('h4)
	) name594 (
		_w210_,
		_w627_,
		_w628_
	);
	LUT4 #(
		.INIT('h153f)
	) name595 (
		_w52_,
		_w67_,
		_w78_,
		_w43_,
		_w629_
	);
	LUT4 #(
		.INIT('h153f)
	) name596 (
		_w52_,
		_w41_,
		_w184_,
		_w430_,
		_w630_
	);
	LUT4 #(
		.INIT('h153f)
	) name597 (
		_w90_,
		_w41_,
		_w259_,
		_w419_,
		_w631_
	);
	LUT3 #(
		.INIT('h80)
	) name598 (
		_w630_,
		_w629_,
		_w631_,
		_w632_
	);
	LUT2 #(
		.INIT('h8)
	) name599 (
		_w628_,
		_w632_,
		_w633_
	);
	LUT4 #(
		.INIT('h135f)
	) name600 (
		_w52_,
		_w90_,
		_w184_,
		_w430_,
		_w634_
	);
	LUT4 #(
		.INIT('h0777)
	) name601 (
		_w106_,
		_w85_,
		_w67_,
		_w378_,
		_w635_
	);
	LUT4 #(
		.INIT('h153f)
	) name602 (
		_w55_,
		_w90_,
		_w43_,
		_w378_,
		_w636_
	);
	LUT4 #(
		.INIT('h0777)
	) name603 (
		_w38_,
		_w106_,
		_w85_,
		_w184_,
		_w637_
	);
	LUT4 #(
		.INIT('h8000)
	) name604 (
		_w634_,
		_w635_,
		_w636_,
		_w637_,
		_w638_
	);
	LUT4 #(
		.INIT('h0777)
	) name605 (
		_w122_,
		_w65_,
		_w44_,
		_w430_,
		_w639_
	);
	LUT2 #(
		.INIT('h4)
	) name606 (
		_w102_,
		_w639_,
		_w640_
	);
	LUT4 #(
		.INIT('h135f)
	) name607 (
		_w59_,
		_w56_,
		_w72_,
		_w184_,
		_w641_
	);
	LUT4 #(
		.INIT('h4000)
	) name608 (
		_w102_,
		_w589_,
		_w641_,
		_w639_,
		_w642_
	);
	LUT4 #(
		.INIT('h153f)
	) name609 (
		_w38_,
		_w85_,
		_w259_,
		_w378_,
		_w643_
	);
	LUT3 #(
		.INIT('h40)
	) name610 (
		_w424_,
		_w611_,
		_w643_,
		_w644_
	);
	LUT4 #(
		.INIT('h135f)
	) name611 (
		_w110_,
		_w50_,
		_w201_,
		_w236_,
		_w645_
	);
	LUT3 #(
		.INIT('h40)
	) name612 (
		_w452_,
		_w605_,
		_w645_,
		_w646_
	);
	LUT4 #(
		.INIT('h8000)
	) name613 (
		_w644_,
		_w646_,
		_w638_,
		_w642_,
		_w647_
	);
	LUT2 #(
		.INIT('h8)
	) name614 (
		_w633_,
		_w647_,
		_w648_
	);
	LUT3 #(
		.INIT('h37)
	) name615 (
		_w106_,
		_w59_,
		_w378_,
		_w649_
	);
	LUT4 #(
		.INIT('h153f)
	) name616 (
		_w52_,
		_w59_,
		_w184_,
		_w378_,
		_w650_
	);
	LUT4 #(
		.INIT('h135f)
	) name617 (
		_w38_,
		_w85_,
		_w78_,
		_w419_,
		_w651_
	);
	LUT4 #(
		.INIT('h135f)
	) name618 (
		_w65_,
		_w44_,
		_w201_,
		_w158_,
		_w652_
	);
	LUT4 #(
		.INIT('h8000)
	) name619 (
		_w649_,
		_w650_,
		_w651_,
		_w652_,
		_w653_
	);
	LUT4 #(
		.INIT('h0800)
	) name620 (
		_w81_,
		_w213_,
		_w221_,
		_w262_,
		_w654_
	);
	LUT3 #(
		.INIT('h80)
	) name621 (
		_w242_,
		_w653_,
		_w654_,
		_w655_
	);
	LUT4 #(
		.INIT('h153f)
	) name622 (
		_w56_,
		_w47_,
		_w201_,
		_w430_,
		_w656_
	);
	LUT4 #(
		.INIT('h135f)
	) name623 (
		_w122_,
		_w93_,
		_w46_,
		_w184_,
		_w657_
	);
	LUT4 #(
		.INIT('h4000)
	) name624 (
		_w461_,
		_w446_,
		_w656_,
		_w657_,
		_w658_
	);
	LUT4 #(
		.INIT('h0777)
	) name625 (
		_w106_,
		_w55_,
		_w72_,
		_w65_,
		_w659_
	);
	LUT3 #(
		.INIT('h57)
	) name626 (
		_w110_,
		_w78_,
		_w378_,
		_w660_
	);
	LUT4 #(
		.INIT('h2000)
	) name627 (
		_w116_,
		_w339_,
		_w659_,
		_w660_,
		_w661_
	);
	LUT4 #(
		.INIT('h135f)
	) name628 (
		_w38_,
		_w85_,
		_w419_,
		_w378_,
		_w662_
	);
	LUT4 #(
		.INIT('h153f)
	) name629 (
		_w85_,
		_w67_,
		_w419_,
		_w430_,
		_w663_
	);
	LUT4 #(
		.INIT('h4000)
	) name630 (
		_w454_,
		_w538_,
		_w662_,
		_w663_,
		_w664_
	);
	LUT4 #(
		.INIT('h8000)
	) name631 (
		_w500_,
		_w658_,
		_w661_,
		_w664_,
		_w665_
	);
	LUT4 #(
		.INIT('h8000)
	) name632 (
		_w633_,
		_w647_,
		_w655_,
		_w665_,
		_w666_
	);
	LUT4 #(
		.INIT('h135f)
	) name633 (
		_w39_,
		_w43_,
		_w93_,
		_w65_,
		_w667_
	);
	LUT4 #(
		.INIT('h135f)
	) name634 (
		_w43_,
		_w65_,
		_w46_,
		_w166_,
		_w668_
	);
	LUT4 #(
		.INIT('h8000)
	) name635 (
		_w305_,
		_w364_,
		_w668_,
		_w667_,
		_w669_
	);
	LUT4 #(
		.INIT('h135f)
	) name636 (
		_w52_,
		_w56_,
		_w72_,
		_w158_,
		_w670_
	);
	LUT4 #(
		.INIT('h153f)
	) name637 (
		_w41_,
		_w39_,
		_w65_,
		_w158_,
		_w671_
	);
	LUT4 #(
		.INIT('h4000)
	) name638 (
		_w355_,
		_w553_,
		_w670_,
		_w671_,
		_w672_
	);
	LUT4 #(
		.INIT('h153f)
	) name639 (
		_w38_,
		_w110_,
		_w166_,
		_w176_,
		_w673_
	);
	LUT3 #(
		.INIT('h40)
	) name640 (
		_w124_,
		_w584_,
		_w673_,
		_w674_
	);
	LUT4 #(
		.INIT('h135f)
	) name641 (
		_w122_,
		_w50_,
		_w93_,
		_w259_,
		_w675_
	);
	LUT4 #(
		.INIT('h153f)
	) name642 (
		_w78_,
		_w41_,
		_w72_,
		_w44_,
		_w676_
	);
	LUT4 #(
		.INIT('h0777)
	) name643 (
		_w110_,
		_w39_,
		_w44_,
		_w236_,
		_w677_
	);
	LUT4 #(
		.INIT('h135f)
	) name644 (
		_w67_,
		_w44_,
		_w166_,
		_w259_,
		_w678_
	);
	LUT4 #(
		.INIT('h8000)
	) name645 (
		_w675_,
		_w676_,
		_w677_,
		_w678_,
		_w679_
	);
	LUT4 #(
		.INIT('h8000)
	) name646 (
		_w674_,
		_w679_,
		_w669_,
		_w672_,
		_w680_
	);
	LUT4 #(
		.INIT('h0777)
	) name647 (
		_w78_,
		_w90_,
		_w56_,
		_w39_,
		_w681_
	);
	LUT4 #(
		.INIT('h153f)
	) name648 (
		_w56_,
		_w39_,
		_w50_,
		_w176_,
		_w682_
	);
	LUT4 #(
		.INIT('h135f)
	) name649 (
		_w106_,
		_w67_,
		_w44_,
		_w176_,
		_w683_
	);
	LUT4 #(
		.INIT('h8000)
	) name650 (
		_w88_,
		_w681_,
		_w682_,
		_w683_,
		_w684_
	);
	LUT4 #(
		.INIT('h153f)
	) name651 (
		_w122_,
		_w59_,
		_w78_,
		_w90_,
		_w685_
	);
	LUT4 #(
		.INIT('h135f)
	) name652 (
		_w38_,
		_w41_,
		_w166_,
		_w176_,
		_w686_
	);
	LUT4 #(
		.INIT('h135f)
	) name653 (
		_w39_,
		_w93_,
		_w44_,
		_w158_,
		_w687_
	);
	LUT4 #(
		.INIT('h8000)
	) name654 (
		_w470_,
		_w687_,
		_w685_,
		_w686_,
		_w688_
	);
	LUT4 #(
		.INIT('h153f)
	) name655 (
		_w55_,
		_w47_,
		_w39_,
		_w166_,
		_w689_
	);
	LUT4 #(
		.INIT('h0777)
	) name656 (
		_w122_,
		_w67_,
		_w47_,
		_w166_,
		_w690_
	);
	LUT4 #(
		.INIT('h1000)
	) name657 (
		_w185_,
		_w451_,
		_w689_,
		_w690_,
		_w691_
	);
	LUT2 #(
		.INIT('h8)
	) name658 (
		_w688_,
		_w691_,
		_w692_
	);
	LUT3 #(
		.INIT('h80)
	) name659 (
		_w684_,
		_w688_,
		_w691_,
		_w693_
	);
	LUT2 #(
		.INIT('h8)
	) name660 (
		_w680_,
		_w693_,
		_w694_
	);
	LUT2 #(
		.INIT('h8)
	) name661 (
		_w666_,
		_w694_,
		_w695_
	);
	LUT3 #(
		.INIT('h1f)
	) name662 (
		_w67_,
		_w90_,
		_w72_,
		_w696_
	);
	LUT4 #(
		.INIT('h135f)
	) name663 (
		_w106_,
		_w78_,
		_w56_,
		_w46_,
		_w697_
	);
	LUT4 #(
		.INIT('h135f)
	) name664 (
		_w55_,
		_w47_,
		_w72_,
		_w236_,
		_w698_
	);
	LUT4 #(
		.INIT('h4000)
	) name665 (
		_w476_,
		_w696_,
		_w697_,
		_w698_,
		_w699_
	);
	LUT3 #(
		.INIT('h1f)
	) name666 (
		_w110_,
		_w44_,
		_w259_,
		_w700_
	);
	LUT4 #(
		.INIT('h135f)
	) name667 (
		_w122_,
		_w59_,
		_w44_,
		_w430_,
		_w701_
	);
	LUT4 #(
		.INIT('h135f)
	) name668 (
		_w85_,
		_w46_,
		_w166_,
		_w158_,
		_w702_
	);
	LUT4 #(
		.INIT('h8000)
	) name669 (
		_w663_,
		_w702_,
		_w700_,
		_w701_,
		_w703_
	);
	LUT4 #(
		.INIT('h135f)
	) name670 (
		_w52_,
		_w41_,
		_w72_,
		_w430_,
		_w704_
	);
	LUT4 #(
		.INIT('h153f)
	) name671 (
		_w106_,
		_w41_,
		_w72_,
		_w65_,
		_w705_
	);
	LUT4 #(
		.INIT('h153f)
	) name672 (
		_w90_,
		_w39_,
		_w65_,
		_w184_,
		_w706_
	);
	LUT3 #(
		.INIT('h57)
	) name673 (
		_w67_,
		_w78_,
		_w378_,
		_w707_
	);
	LUT4 #(
		.INIT('h8000)
	) name674 (
		_w704_,
		_w706_,
		_w707_,
		_w705_,
		_w708_
	);
	LUT3 #(
		.INIT('h80)
	) name675 (
		_w703_,
		_w699_,
		_w708_,
		_w709_
	);
	LUT4 #(
		.INIT('h153f)
	) name676 (
		_w52_,
		_w93_,
		_w158_,
		_w430_,
		_w710_
	);
	LUT4 #(
		.INIT('h135f)
	) name677 (
		_w85_,
		_w46_,
		_w184_,
		_w430_,
		_w711_
	);
	LUT3 #(
		.INIT('h40)
	) name678 (
		_w230_,
		_w711_,
		_w710_,
		_w712_
	);
	LUT3 #(
		.INIT('h1f)
	) name679 (
		_w93_,
		_w44_,
		_w184_,
		_w713_
	);
	LUT4 #(
		.INIT('h153f)
	) name680 (
		_w110_,
		_w78_,
		_w50_,
		_w43_,
		_w714_
	);
	LUT4 #(
		.INIT('h1000)
	) name681 (
		_w206_,
		_w413_,
		_w713_,
		_w714_,
		_w715_
	);
	LUT2 #(
		.INIT('h8)
	) name682 (
		_w712_,
		_w715_,
		_w716_
	);
	LUT4 #(
		.INIT('h0777)
	) name683 (
		_w78_,
		_w90_,
		_w93_,
		_w236_,
		_w717_
	);
	LUT4 #(
		.INIT('h135f)
	) name684 (
		_w41_,
		_w50_,
		_w419_,
		_w378_,
		_w718_
	);
	LUT2 #(
		.INIT('h8)
	) name685 (
		_w717_,
		_w718_,
		_w719_
	);
	LUT4 #(
		.INIT('h153f)
	) name686 (
		_w90_,
		_w44_,
		_w419_,
		_w378_,
		_w720_
	);
	LUT4 #(
		.INIT('h135f)
	) name687 (
		_w55_,
		_w59_,
		_w43_,
		_w184_,
		_w721_
	);
	LUT3 #(
		.INIT('h1f)
	) name688 (
		_w90_,
		_w44_,
		_w166_,
		_w722_
	);
	LUT4 #(
		.INIT('h4000)
	) name689 (
		_w436_,
		_w720_,
		_w721_,
		_w722_,
		_w723_
	);
	LUT4 #(
		.INIT('h8000)
	) name690 (
		_w712_,
		_w715_,
		_w719_,
		_w723_,
		_w724_
	);
	LUT3 #(
		.INIT('h80)
	) name691 (
		_w328_,
		_w709_,
		_w724_,
		_w725_
	);
	LUT4 #(
		.INIT('h0777)
	) name692 (
		_w56_,
		_w72_,
		_w50_,
		_w158_,
		_w726_
	);
	LUT2 #(
		.INIT('h4)
	) name693 (
		_w451_,
		_w726_,
		_w727_
	);
	LUT4 #(
		.INIT('h153f)
	) name694 (
		_w52_,
		_w43_,
		_w46_,
		_w166_,
		_w728_
	);
	LUT4 #(
		.INIT('h2000)
	) name695 (
		_w252_,
		_w402_,
		_w514_,
		_w728_,
		_w729_
	);
	LUT2 #(
		.INIT('h8)
	) name696 (
		_w727_,
		_w729_,
		_w730_
	);
	LUT4 #(
		.INIT('h135f)
	) name697 (
		_w122_,
		_w52_,
		_w110_,
		_w259_,
		_w731_
	);
	LUT4 #(
		.INIT('h135f)
	) name698 (
		_w52_,
		_w46_,
		_w184_,
		_w236_,
		_w732_
	);
	LUT3 #(
		.INIT('h40)
	) name699 (
		_w282_,
		_w731_,
		_w732_,
		_w733_
	);
	LUT4 #(
		.INIT('h135f)
	) name700 (
		_w110_,
		_w90_,
		_w72_,
		_w39_,
		_w734_
	);
	LUT4 #(
		.INIT('h135f)
	) name701 (
		_w122_,
		_w59_,
		_w56_,
		_w176_,
		_w735_
	);
	LUT3 #(
		.INIT('h40)
	) name702 (
		_w392_,
		_w734_,
		_w735_,
		_w736_
	);
	LUT3 #(
		.INIT('h37)
	) name703 (
		_w39_,
		_w44_,
		_w378_,
		_w737_
	);
	LUT4 #(
		.INIT('h153f)
	) name704 (
		_w59_,
		_w56_,
		_w201_,
		_w166_,
		_w738_
	);
	LUT4 #(
		.INIT('h153f)
	) name705 (
		_w55_,
		_w39_,
		_w50_,
		_w184_,
		_w739_
	);
	LUT3 #(
		.INIT('h80)
	) name706 (
		_w738_,
		_w739_,
		_w737_,
		_w740_
	);
	LUT3 #(
		.INIT('h80)
	) name707 (
		_w736_,
		_w733_,
		_w740_,
		_w741_
	);
	LUT4 #(
		.INIT('h135f)
	) name708 (
		_w55_,
		_w41_,
		_w39_,
		_w236_,
		_w742_
	);
	LUT3 #(
		.INIT('h37)
	) name709 (
		_w78_,
		_w93_,
		_w259_,
		_w743_
	);
	LUT4 #(
		.INIT('h153f)
	) name710 (
		_w47_,
		_w44_,
		_w176_,
		_w419_,
		_w744_
	);
	LUT3 #(
		.INIT('h80)
	) name711 (
		_w743_,
		_w744_,
		_w742_,
		_w745_
	);
	LUT4 #(
		.INIT('h135f)
	) name712 (
		_w52_,
		_w56_,
		_w201_,
		_w166_,
		_w746_
	);
	LUT4 #(
		.INIT('h0777)
	) name713 (
		_w78_,
		_w41_,
		_w46_,
		_w176_,
		_w747_
	);
	LUT4 #(
		.INIT('h1000)
	) name714 (
		_w276_,
		_w432_,
		_w746_,
		_w747_,
		_w748_
	);
	LUT2 #(
		.INIT('h8)
	) name715 (
		_w745_,
		_w748_,
		_w749_
	);
	LUT4 #(
		.INIT('h0777)
	) name716 (
		_w55_,
		_w78_,
		_w44_,
		_w158_,
		_w750_
	);
	LUT2 #(
		.INIT('h8)
	) name717 (
		_w496_,
		_w750_,
		_w751_
	);
	LUT4 #(
		.INIT('h131f)
	) name718 (
		_w52_,
		_w50_,
		_w43_,
		_w166_,
		_w752_
	);
	LUT4 #(
		.INIT('h153f)
	) name719 (
		_w59_,
		_w110_,
		_w78_,
		_w201_,
		_w753_
	);
	LUT3 #(
		.INIT('h40)
	) name720 (
		_w426_,
		_w752_,
		_w753_,
		_w754_
	);
	LUT4 #(
		.INIT('h135f)
	) name721 (
		_w110_,
		_w56_,
		_w236_,
		_w419_,
		_w755_
	);
	LUT4 #(
		.INIT('h0200)
	) name722 (
		_w361_,
		_w406_,
		_w468_,
		_w755_,
		_w756_
	);
	LUT4 #(
		.INIT('h135f)
	) name723 (
		_w122_,
		_w110_,
		_w50_,
		_w419_,
		_w757_
	);
	LUT4 #(
		.INIT('h0777)
	) name724 (
		_w59_,
		_w78_,
		_w44_,
		_w201_,
		_w758_
	);
	LUT4 #(
		.INIT('h153f)
	) name725 (
		_w38_,
		_w50_,
		_w184_,
		_w378_,
		_w759_
	);
	LUT4 #(
		.INIT('h153f)
	) name726 (
		_w50_,
		_w93_,
		_w201_,
		_w236_,
		_w760_
	);
	LUT4 #(
		.INIT('h8000)
	) name727 (
		_w757_,
		_w759_,
		_w760_,
		_w758_,
		_w761_
	);
	LUT4 #(
		.INIT('h8000)
	) name728 (
		_w756_,
		_w751_,
		_w761_,
		_w754_,
		_w762_
	);
	LUT2 #(
		.INIT('h8)
	) name729 (
		_w749_,
		_w762_,
		_w763_
	);
	LUT4 #(
		.INIT('h8000)
	) name730 (
		_w730_,
		_w741_,
		_w749_,
		_w762_,
		_w764_
	);
	LUT2 #(
		.INIT('h8)
	) name731 (
		_w725_,
		_w764_,
		_w765_
	);
	LUT4 #(
		.INIT('h0777)
	) name732 (
		_w666_,
		_w694_,
		_w725_,
		_w764_,
		_w766_
	);
	LUT4 #(
		.INIT('h135f)
	) name733 (
		_w85_,
		_w50_,
		_w166_,
		_w176_,
		_w767_
	);
	LUT4 #(
		.INIT('h135f)
	) name734 (
		_w67_,
		_w46_,
		_w259_,
		_w176_,
		_w768_
	);
	LUT4 #(
		.INIT('h135f)
	) name735 (
		_w122_,
		_w106_,
		_w85_,
		_w47_,
		_w769_
	);
	LUT4 #(
		.INIT('h153f)
	) name736 (
		_w59_,
		_w39_,
		_w93_,
		_w201_,
		_w770_
	);
	LUT4 #(
		.INIT('h8000)
	) name737 (
		_w767_,
		_w768_,
		_w769_,
		_w770_,
		_w771_
	);
	LUT4 #(
		.INIT('h153f)
	) name738 (
		_w55_,
		_w85_,
		_w184_,
		_w378_,
		_w772_
	);
	LUT2 #(
		.INIT('h8)
	) name739 (
		_w731_,
		_w772_,
		_w773_
	);
	LUT3 #(
		.INIT('h57)
	) name740 (
		_w85_,
		_w43_,
		_w201_,
		_w774_
	);
	LUT4 #(
		.INIT('h153f)
	) name741 (
		_w90_,
		_w41_,
		_w378_,
		_w430_,
		_w775_
	);
	LUT4 #(
		.INIT('h153f)
	) name742 (
		_w55_,
		_w65_,
		_w166_,
		_w176_,
		_w776_
	);
	LUT4 #(
		.INIT('h0777)
	) name743 (
		_w106_,
		_w110_,
		_w44_,
		_w430_,
		_w777_
	);
	LUT4 #(
		.INIT('h8000)
	) name744 (
		_w776_,
		_w777_,
		_w774_,
		_w775_,
		_w778_
	);
	LUT3 #(
		.INIT('h80)
	) name745 (
		_w773_,
		_w771_,
		_w778_,
		_w779_
	);
	LUT4 #(
		.INIT('h135f)
	) name746 (
		_w56_,
		_w46_,
		_w184_,
		_w419_,
		_w780_
	);
	LUT4 #(
		.INIT('h0777)
	) name747 (
		_w52_,
		_w78_,
		_w41_,
		_w176_,
		_w781_
	);
	LUT3 #(
		.INIT('h80)
	) name748 (
		_w265_,
		_w781_,
		_w780_,
		_w782_
	);
	LUT3 #(
		.INIT('h57)
	) name749 (
		_w90_,
		_w72_,
		_w158_,
		_w783_
	);
	LUT4 #(
		.INIT('h153f)
	) name750 (
		_w55_,
		_w67_,
		_w39_,
		_w43_,
		_w784_
	);
	LUT3 #(
		.INIT('h57)
	) name751 (
		_w47_,
		_w43_,
		_w201_,
		_w785_
	);
	LUT4 #(
		.INIT('h4000)
	) name752 (
		_w152_,
		_w783_,
		_w784_,
		_w785_,
		_w786_
	);
	LUT4 #(
		.INIT('h131f)
	) name753 (
		_w41_,
		_w44_,
		_w158_,
		_w378_,
		_w787_
	);
	LUT4 #(
		.INIT('h153f)
	) name754 (
		_w90_,
		_w43_,
		_w44_,
		_w378_,
		_w788_
	);
	LUT4 #(
		.INIT('h153f)
	) name755 (
		_w38_,
		_w55_,
		_w184_,
		_w236_,
		_w789_
	);
	LUT3 #(
		.INIT('h37)
	) name756 (
		_w85_,
		_w72_,
		_w46_,
		_w790_
	);
	LUT4 #(
		.INIT('h8000)
	) name757 (
		_w582_,
		_w788_,
		_w789_,
		_w790_,
		_w791_
	);
	LUT4 #(
		.INIT('h8000)
	) name758 (
		_w782_,
		_w786_,
		_w787_,
		_w791_,
		_w792_
	);
	LUT4 #(
		.INIT('h153f)
	) name759 (
		_w38_,
		_w55_,
		_w72_,
		_w430_,
		_w793_
	);
	LUT4 #(
		.INIT('h153f)
	) name760 (
		_w47_,
		_w65_,
		_w236_,
		_w419_,
		_w794_
	);
	LUT4 #(
		.INIT('h0777)
	) name761 (
		_w122_,
		_w55_,
		_w44_,
		_w176_,
		_w795_
	);
	LUT4 #(
		.INIT('h4000)
	) name762 (
		_w353_,
		_w793_,
		_w794_,
		_w795_,
		_w796_
	);
	LUT4 #(
		.INIT('h153f)
	) name763 (
		_w90_,
		_w47_,
		_w166_,
		_w259_,
		_w797_
	);
	LUT4 #(
		.INIT('h153f)
	) name764 (
		_w47_,
		_w46_,
		_w184_,
		_w158_,
		_w798_
	);
	LUT4 #(
		.INIT('h2000)
	) name765 (
		_w132_,
		_w429_,
		_w797_,
		_w798_,
		_w799_
	);
	LUT2 #(
		.INIT('h8)
	) name766 (
		_w796_,
		_w799_,
		_w800_
	);
	LUT3 #(
		.INIT('h80)
	) name767 (
		_w779_,
		_w792_,
		_w800_,
		_w801_
	);
	LUT4 #(
		.INIT('h153f)
	) name768 (
		_w110_,
		_w43_,
		_w93_,
		_w158_,
		_w802_
	);
	LUT3 #(
		.INIT('h1f)
	) name769 (
		_w122_,
		_w78_,
		_w50_,
		_w803_
	);
	LUT4 #(
		.INIT('h135f)
	) name770 (
		_w52_,
		_w41_,
		_w201_,
		_w430_,
		_w804_
	);
	LUT3 #(
		.INIT('h80)
	) name771 (
		_w803_,
		_w804_,
		_w802_,
		_w805_
	);
	LUT3 #(
		.INIT('h57)
	) name772 (
		_w110_,
		_w72_,
		_w259_,
		_w806_
	);
	LUT4 #(
		.INIT('h135f)
	) name773 (
		_w52_,
		_w90_,
		_w39_,
		_w201_,
		_w807_
	);
	LUT4 #(
		.INIT('h135f)
	) name774 (
		_w59_,
		_w67_,
		_w166_,
		_w158_,
		_w808_
	);
	LUT4 #(
		.INIT('h153f)
	) name775 (
		_w110_,
		_w46_,
		_w166_,
		_w419_,
		_w809_
	);
	LUT4 #(
		.INIT('h8000)
	) name776 (
		_w806_,
		_w807_,
		_w808_,
		_w809_,
		_w810_
	);
	LUT4 #(
		.INIT('h135f)
	) name777 (
		_w55_,
		_w93_,
		_w236_,
		_w158_,
		_w811_
	);
	LUT4 #(
		.INIT('h4000)
	) name778 (
		_w79_,
		_w348_,
		_w583_,
		_w811_,
		_w812_
	);
	LUT3 #(
		.INIT('h80)
	) name779 (
		_w805_,
		_w810_,
		_w812_,
		_w813_
	);
	LUT4 #(
		.INIT('h153f)
	) name780 (
		_w56_,
		_w44_,
		_w166_,
		_w259_,
		_w814_
	);
	LUT2 #(
		.INIT('h4)
	) name781 (
		_w334_,
		_w814_,
		_w815_
	);
	LUT4 #(
		.INIT('h0777)
	) name782 (
		_w122_,
		_w56_,
		_w50_,
		_w419_,
		_w816_
	);
	LUT4 #(
		.INIT('h0777)
	) name783 (
		_w106_,
		_w55_,
		_w65_,
		_w430_,
		_w817_
	);
	LUT3 #(
		.INIT('h1f)
	) name784 (
		_w39_,
		_w43_,
		_w46_,
		_w818_
	);
	LUT3 #(
		.INIT('h80)
	) name785 (
		_w817_,
		_w816_,
		_w818_,
		_w819_
	);
	LUT4 #(
		.INIT('h135f)
	) name786 (
		_w110_,
		_w46_,
		_w201_,
		_w430_,
		_w820_
	);
	LUT4 #(
		.INIT('h135f)
	) name787 (
		_w38_,
		_w55_,
		_w39_,
		_w430_,
		_w821_
	);
	LUT2 #(
		.INIT('h8)
	) name788 (
		_w820_,
		_w821_,
		_w822_
	);
	LUT3 #(
		.INIT('h1f)
	) name789 (
		_w50_,
		_w93_,
		_w236_,
		_w823_
	);
	LUT4 #(
		.INIT('h153f)
	) name790 (
		_w110_,
		_w90_,
		_w166_,
		_w378_,
		_w824_
	);
	LUT4 #(
		.INIT('h0777)
	) name791 (
		_w38_,
		_w122_,
		_w46_,
		_w259_,
		_w825_
	);
	LUT4 #(
		.INIT('h4000)
	) name792 (
		_w314_,
		_w823_,
		_w824_,
		_w825_,
		_w826_
	);
	LUT4 #(
		.INIT('h8000)
	) name793 (
		_w822_,
		_w815_,
		_w819_,
		_w826_,
		_w827_
	);
	LUT4 #(
		.INIT('h0777)
	) name794 (
		_w72_,
		_w50_,
		_w46_,
		_w201_,
		_w828_
	);
	LUT4 #(
		.INIT('h135f)
	) name795 (
		_w106_,
		_w56_,
		_w46_,
		_w378_,
		_w829_
	);
	LUT4 #(
		.INIT('h0777)
	) name796 (
		_w59_,
		_w78_,
		_w41_,
		_w43_,
		_w830_
	);
	LUT4 #(
		.INIT('h4000)
	) name797 (
		_w244_,
		_w828_,
		_w829_,
		_w830_,
		_w831_
	);
	LUT4 #(
		.INIT('h0777)
	) name798 (
		_w110_,
		_w78_,
		_w44_,
		_w259_,
		_w832_
	);
	LUT2 #(
		.INIT('h4)
	) name799 (
		_w439_,
		_w832_,
		_w833_
	);
	LUT4 #(
		.INIT('h153f)
	) name800 (
		_w85_,
		_w65_,
		_w158_,
		_w259_,
		_w834_
	);
	LUT4 #(
		.INIT('h153f)
	) name801 (
		_w106_,
		_w55_,
		_w78_,
		_w41_,
		_w835_
	);
	LUT4 #(
		.INIT('h4000)
	) name802 (
		_w439_,
		_w832_,
		_w834_,
		_w835_,
		_w836_
	);
	LUT2 #(
		.INIT('h8)
	) name803 (
		_w831_,
		_w836_,
		_w837_
	);
	LUT3 #(
		.INIT('h37)
	) name804 (
		_w122_,
		_w59_,
		_w259_,
		_w838_
	);
	LUT4 #(
		.INIT('h153f)
	) name805 (
		_w59_,
		_w47_,
		_w39_,
		_w43_,
		_w839_
	);
	LUT3 #(
		.INIT('h37)
	) name806 (
		_w56_,
		_w72_,
		_w65_,
		_w840_
	);
	LUT4 #(
		.INIT('h4000)
	) name807 (
		_w445_,
		_w839_,
		_w840_,
		_w838_,
		_w841_
	);
	LUT4 #(
		.INIT('h135f)
	) name808 (
		_w67_,
		_w50_,
		_w43_,
		_w158_,
		_w842_
	);
	LUT4 #(
		.INIT('h153f)
	) name809 (
		_w67_,
		_w56_,
		_w158_,
		_w430_,
		_w843_
	);
	LUT4 #(
		.INIT('h135f)
	) name810 (
		_w90_,
		_w47_,
		_w39_,
		_w259_,
		_w844_
	);
	LUT4 #(
		.INIT('h8000)
	) name811 (
		_w650_,
		_w842_,
		_w843_,
		_w844_,
		_w845_
	);
	LUT4 #(
		.INIT('h135f)
	) name812 (
		_w122_,
		_w52_,
		_w47_,
		_w184_,
		_w846_
	);
	LUT4 #(
		.INIT('h135f)
	) name813 (
		_w41_,
		_w44_,
		_w184_,
		_w236_,
		_w847_
	);
	LUT4 #(
		.INIT('h153f)
	) name814 (
		_w52_,
		_w41_,
		_w39_,
		_w166_,
		_w848_
	);
	LUT4 #(
		.INIT('h4000)
	) name815 (
		_w359_,
		_w846_,
		_w847_,
		_w848_,
		_w849_
	);
	LUT3 #(
		.INIT('h80)
	) name816 (
		_w841_,
		_w845_,
		_w849_,
		_w850_
	);
	LUT4 #(
		.INIT('h8000)
	) name817 (
		_w813_,
		_w827_,
		_w837_,
		_w850_,
		_w851_
	);
	LUT2 #(
		.INIT('h8)
	) name818 (
		_w801_,
		_w851_,
		_w852_
	);
	LUT4 #(
		.INIT('h153f)
	) name819 (
		_w55_,
		_w85_,
		_w72_,
		_w43_,
		_w853_
	);
	LUT4 #(
		.INIT('h8000)
	) name820 (
		_w68_,
		_w391_,
		_w394_,
		_w853_,
		_w854_
	);
	LUT4 #(
		.INIT('h153f)
	) name821 (
		_w85_,
		_w78_,
		_w46_,
		_w236_,
		_w855_
	);
	LUT4 #(
		.INIT('h153f)
	) name822 (
		_w90_,
		_w56_,
		_w378_,
		_w430_,
		_w856_
	);
	LUT4 #(
		.INIT('h135f)
	) name823 (
		_w55_,
		_w47_,
		_w158_,
		_w259_,
		_w857_
	);
	LUT4 #(
		.INIT('h4000)
	) name824 (
		_w412_,
		_w855_,
		_w856_,
		_w857_,
		_w858_
	);
	LUT2 #(
		.INIT('h8)
	) name825 (
		_w854_,
		_w858_,
		_w859_
	);
	LUT4 #(
		.INIT('h153f)
	) name826 (
		_w56_,
		_w44_,
		_w236_,
		_w259_,
		_w860_
	);
	LUT4 #(
		.INIT('h153f)
	) name827 (
		_w38_,
		_w67_,
		_w166_,
		_w430_,
		_w861_
	);
	LUT3 #(
		.INIT('h80)
	) name828 (
		_w281_,
		_w861_,
		_w860_,
		_w862_
	);
	LUT4 #(
		.INIT('h135f)
	) name829 (
		_w44_,
		_w46_,
		_w184_,
		_w419_,
		_w863_
	);
	LUT4 #(
		.INIT('h153f)
	) name830 (
		_w50_,
		_w43_,
		_w93_,
		_w201_,
		_w864_
	);
	LUT4 #(
		.INIT('h135f)
	) name831 (
		_w106_,
		_w52_,
		_w47_,
		_w72_,
		_w865_
	);
	LUT3 #(
		.INIT('h80)
	) name832 (
		_w864_,
		_w865_,
		_w863_,
		_w866_
	);
	LUT4 #(
		.INIT('h135f)
	) name833 (
		_w52_,
		_w41_,
		_w184_,
		_w430_,
		_w867_
	);
	LUT4 #(
		.INIT('h0777)
	) name834 (
		_w78_,
		_w41_,
		_w65_,
		_w158_,
		_w868_
	);
	LUT4 #(
		.INIT('h8000)
	) name835 (
		_w216_,
		_w768_,
		_w867_,
		_w868_,
		_w869_
	);
	LUT3 #(
		.INIT('h80)
	) name836 (
		_w862_,
		_w866_,
		_w869_,
		_w870_
	);
	LUT2 #(
		.INIT('h8)
	) name837 (
		_w859_,
		_w870_,
		_w871_
	);
	LUT4 #(
		.INIT('h135f)
	) name838 (
		_w38_,
		_w90_,
		_w201_,
		_w176_,
		_w872_
	);
	LUT4 #(
		.INIT('h153f)
	) name839 (
		_w93_,
		_w65_,
		_w378_,
		_w430_,
		_w873_
	);
	LUT4 #(
		.INIT('h0777)
	) name840 (
		_w38_,
		_w106_,
		_w56_,
		_w39_,
		_w874_
	);
	LUT4 #(
		.INIT('h4000)
	) name841 (
		_w429_,
		_w873_,
		_w874_,
		_w872_,
		_w875_
	);
	LUT4 #(
		.INIT('h135f)
	) name842 (
		_w122_,
		_w59_,
		_w50_,
		_w419_,
		_w876_
	);
	LUT4 #(
		.INIT('h0777)
	) name843 (
		_w106_,
		_w67_,
		_w44_,
		_w158_,
		_w877_
	);
	LUT4 #(
		.INIT('h153f)
	) name844 (
		_w56_,
		_w46_,
		_w166_,
		_w176_,
		_w878_
	);
	LUT2 #(
		.INIT('h8)
	) name845 (
		_w877_,
		_w878_,
		_w879_
	);
	LUT4 #(
		.INIT('h4000)
	) name846 (
		_w107_,
		_w876_,
		_w877_,
		_w878_,
		_w880_
	);
	LUT2 #(
		.INIT('h8)
	) name847 (
		_w875_,
		_w880_,
		_w881_
	);
	LUT4 #(
		.INIT('h153f)
	) name848 (
		_w52_,
		_w93_,
		_w166_,
		_w158_,
		_w882_
	);
	LUT2 #(
		.INIT('h4)
	) name849 (
		_w468_,
		_w882_,
		_w883_
	);
	LUT3 #(
		.INIT('h37)
	) name850 (
		_w78_,
		_w50_,
		_w158_,
		_w884_
	);
	LUT4 #(
		.INIT('h135f)
	) name851 (
		_w55_,
		_w52_,
		_w419_,
		_w430_,
		_w885_
	);
	LUT4 #(
		.INIT('h135f)
	) name852 (
		_w56_,
		_w47_,
		_w184_,
		_w158_,
		_w886_
	);
	LUT4 #(
		.INIT('h135f)
	) name853 (
		_w38_,
		_w85_,
		_w72_,
		_w39_,
		_w887_
	);
	LUT4 #(
		.INIT('h8000)
	) name854 (
		_w886_,
		_w887_,
		_w884_,
		_w885_,
		_w888_
	);
	LUT4 #(
		.INIT('h0777)
	) name855 (
		_w122_,
		_w85_,
		_w44_,
		_w201_,
		_w889_
	);
	LUT4 #(
		.INIT('h135f)
	) name856 (
		_w85_,
		_w67_,
		_w43_,
		_w176_,
		_w890_
	);
	LUT3 #(
		.INIT('h40)
	) name857 (
		_w362_,
		_w890_,
		_w889_,
		_w891_
	);
	LUT3 #(
		.INIT('h37)
	) name858 (
		_w78_,
		_w47_,
		_w430_,
		_w892_
	);
	LUT4 #(
		.INIT('h135f)
	) name859 (
		_w85_,
		_w52_,
		_w78_,
		_w176_,
		_w893_
	);
	LUT3 #(
		.INIT('h57)
	) name860 (
		_w67_,
		_w43_,
		_w378_,
		_w894_
	);
	LUT4 #(
		.INIT('h135f)
	) name861 (
		_w78_,
		_w90_,
		_w44_,
		_w378_,
		_w895_
	);
	LUT4 #(
		.INIT('h8000)
	) name862 (
		_w892_,
		_w893_,
		_w894_,
		_w895_,
		_w896_
	);
	LUT4 #(
		.INIT('h8000)
	) name863 (
		_w883_,
		_w891_,
		_w896_,
		_w888_,
		_w897_
	);
	LUT3 #(
		.INIT('h02)
	) name864 (
		_w245_,
		_w457_,
		_w437_,
		_w898_
	);
	LUT4 #(
		.INIT('h135f)
	) name865 (
		_w106_,
		_w110_,
		_w93_,
		_w176_,
		_w899_
	);
	LUT3 #(
		.INIT('h1f)
	) name866 (
		_w90_,
		_w46_,
		_w158_,
		_w900_
	);
	LUT4 #(
		.INIT('h153f)
	) name867 (
		_w52_,
		_w41_,
		_w39_,
		_w43_,
		_w901_
	);
	LUT4 #(
		.INIT('h135f)
	) name868 (
		_w41_,
		_w50_,
		_w184_,
		_w166_,
		_w902_
	);
	LUT4 #(
		.INIT('h8000)
	) name869 (
		_w899_,
		_w900_,
		_w901_,
		_w902_,
		_w903_
	);
	LUT4 #(
		.INIT('h0737)
	) name870 (
		_w38_,
		_w122_,
		_w41_,
		_w259_,
		_w904_
	);
	LUT4 #(
		.INIT('h135f)
	) name871 (
		_w55_,
		_w110_,
		_w72_,
		_w43_,
		_w905_
	);
	LUT4 #(
		.INIT('h153f)
	) name872 (
		_w52_,
		_w67_,
		_w201_,
		_w166_,
		_w906_
	);
	LUT3 #(
		.INIT('h80)
	) name873 (
		_w905_,
		_w906_,
		_w904_,
		_w907_
	);
	LUT4 #(
		.INIT('h135f)
	) name874 (
		_w38_,
		_w106_,
		_w78_,
		_w50_,
		_w908_
	);
	LUT4 #(
		.INIT('h0777)
	) name875 (
		_w56_,
		_w43_,
		_w93_,
		_w419_,
		_w909_
	);
	LUT4 #(
		.INIT('h135f)
	) name876 (
		_w38_,
		_w55_,
		_w43_,
		_w378_,
		_w910_
	);
	LUT3 #(
		.INIT('h80)
	) name877 (
		_w909_,
		_w908_,
		_w910_,
		_w911_
	);
	LUT4 #(
		.INIT('h8000)
	) name878 (
		_w898_,
		_w907_,
		_w911_,
		_w903_,
		_w912_
	);
	LUT4 #(
		.INIT('h0777)
	) name879 (
		_w106_,
		_w52_,
		_w59_,
		_w72_,
		_w913_
	);
	LUT4 #(
		.INIT('h135f)
	) name880 (
		_w47_,
		_w50_,
		_w184_,
		_w176_,
		_w914_
	);
	LUT2 #(
		.INIT('h8)
	) name881 (
		_w913_,
		_w914_,
		_w915_
	);
	LUT4 #(
		.INIT('h153f)
	) name882 (
		_w90_,
		_w47_,
		_w39_,
		_w184_,
		_w916_
	);
	LUT4 #(
		.INIT('h135f)
	) name883 (
		_w122_,
		_w110_,
		_w47_,
		_w39_,
		_w917_
	);
	LUT4 #(
		.INIT('h135f)
	) name884 (
		_w122_,
		_w47_,
		_w65_,
		_w419_,
		_w918_
	);
	LUT4 #(
		.INIT('h135f)
	) name885 (
		_w38_,
		_w46_,
		_w158_,
		_w259_,
		_w919_
	);
	LUT4 #(
		.INIT('h8000)
	) name886 (
		_w916_,
		_w918_,
		_w919_,
		_w917_,
		_w920_
	);
	LUT4 #(
		.INIT('h153f)
	) name887 (
		_w110_,
		_w41_,
		_w43_,
		_w166_,
		_w921_
	);
	LUT2 #(
		.INIT('h8)
	) name888 (
		_w252_,
		_w921_,
		_w922_
	);
	LUT4 #(
		.INIT('h135f)
	) name889 (
		_w106_,
		_w85_,
		_w41_,
		_w166_,
		_w923_
	);
	LUT3 #(
		.INIT('h57)
	) name890 (
		_w52_,
		_w78_,
		_w236_,
		_w924_
	);
	LUT4 #(
		.INIT('h4000)
	) name891 (
		_w454_,
		_w789_,
		_w924_,
		_w923_,
		_w925_
	);
	LUT4 #(
		.INIT('h8000)
	) name892 (
		_w915_,
		_w920_,
		_w922_,
		_w925_,
		_w926_
	);
	LUT4 #(
		.INIT('h8000)
	) name893 (
		_w881_,
		_w897_,
		_w912_,
		_w926_,
		_w927_
	);
	LUT2 #(
		.INIT('h8)
	) name894 (
		_w871_,
		_w927_,
		_w928_
	);
	LUT4 #(
		.INIT('h0777)
	) name895 (
		_w801_,
		_w851_,
		_w871_,
		_w927_,
		_w929_
	);
	LUT4 #(
		.INIT('h153f)
	) name896 (
		_w110_,
		_w65_,
		_w201_,
		_w430_,
		_w930_
	);
	LUT4 #(
		.INIT('h135f)
	) name897 (
		_w67_,
		_w50_,
		_w378_,
		_w430_,
		_w931_
	);
	LUT4 #(
		.INIT('h8000)
	) name898 (
		_w95_,
		_w342_,
		_w931_,
		_w930_,
		_w932_
	);
	LUT4 #(
		.INIT('h153f)
	) name899 (
		_w52_,
		_w110_,
		_w166_,
		_w378_,
		_w933_
	);
	LUT3 #(
		.INIT('h80)
	) name900 (
		_w403_,
		_w783_,
		_w933_,
		_w934_
	);
	LUT4 #(
		.INIT('h135f)
	) name901 (
		_w122_,
		_w55_,
		_w85_,
		_w72_,
		_w935_
	);
	LUT4 #(
		.INIT('h0777)
	) name902 (
		_w106_,
		_w59_,
		_w65_,
		_w158_,
		_w936_
	);
	LUT4 #(
		.INIT('h153f)
	) name903 (
		_w55_,
		_w56_,
		_w72_,
		_w201_,
		_w937_
	);
	LUT3 #(
		.INIT('h80)
	) name904 (
		_w936_,
		_w937_,
		_w935_,
		_w938_
	);
	LUT3 #(
		.INIT('h80)
	) name905 (
		_w934_,
		_w932_,
		_w938_,
		_w939_
	);
	LUT4 #(
		.INIT('h0777)
	) name906 (
		_w90_,
		_w39_,
		_w46_,
		_w259_,
		_w940_
	);
	LUT4 #(
		.INIT('h0777)
	) name907 (
		_w38_,
		_w72_,
		_w46_,
		_w166_,
		_w941_
	);
	LUT4 #(
		.INIT('h153f)
	) name908 (
		_w55_,
		_w52_,
		_w166_,
		_w419_,
		_w942_
	);
	LUT3 #(
		.INIT('h80)
	) name909 (
		_w941_,
		_w942_,
		_w940_,
		_w943_
	);
	LUT4 #(
		.INIT('h153f)
	) name910 (
		_w38_,
		_w67_,
		_w39_,
		_w166_,
		_w944_
	);
	LUT4 #(
		.INIT('h135f)
	) name911 (
		_w55_,
		_w59_,
		_w236_,
		_w378_,
		_w945_
	);
	LUT4 #(
		.INIT('h153f)
	) name912 (
		_w65_,
		_w46_,
		_w158_,
		_w419_,
		_w946_
	);
	LUT4 #(
		.INIT('h8000)
	) name913 (
		_w312_,
		_w945_,
		_w944_,
		_w946_,
		_w947_
	);
	LUT4 #(
		.INIT('h0777)
	) name914 (
		_w106_,
		_w55_,
		_w46_,
		_w430_,
		_w948_
	);
	LUT4 #(
		.INIT('h153f)
	) name915 (
		_w122_,
		_w41_,
		_w39_,
		_w65_,
		_w949_
	);
	LUT4 #(
		.INIT('h153f)
	) name916 (
		_w38_,
		_w56_,
		_w184_,
		_w158_,
		_w950_
	);
	LUT4 #(
		.INIT('h135f)
	) name917 (
		_w85_,
		_w59_,
		_w158_,
		_w176_,
		_w951_
	);
	LUT4 #(
		.INIT('h8000)
	) name918 (
		_w948_,
		_w949_,
		_w950_,
		_w951_,
		_w952_
	);
	LUT4 #(
		.INIT('h135f)
	) name919 (
		_w122_,
		_w85_,
		_w67_,
		_w43_,
		_w953_
	);
	LUT4 #(
		.INIT('h1000)
	) name920 (
		_w118_,
		_w223_,
		_w663_,
		_w953_,
		_w954_
	);
	LUT4 #(
		.INIT('h8000)
	) name921 (
		_w943_,
		_w947_,
		_w952_,
		_w954_,
		_w955_
	);
	LUT4 #(
		.INIT('h135f)
	) name922 (
		_w72_,
		_w93_,
		_w65_,
		_w158_,
		_w956_
	);
	LUT4 #(
		.INIT('h0777)
	) name923 (
		_w122_,
		_w47_,
		_w44_,
		_w378_,
		_w957_
	);
	LUT4 #(
		.INIT('h0777)
	) name924 (
		_w106_,
		_w90_,
		_w50_,
		_w176_,
		_w958_
	);
	LUT4 #(
		.INIT('h8000)
	) name925 (
		_w662_,
		_w956_,
		_w957_,
		_w958_,
		_w959_
	);
	LUT4 #(
		.INIT('h0777)
	) name926 (
		_w122_,
		_w52_,
		_w47_,
		_w201_,
		_w960_
	);
	LUT4 #(
		.INIT('h1000)
	) name927 (
		_w275_,
		_w455_,
		_w706_,
		_w960_,
		_w961_
	);
	LUT4 #(
		.INIT('h153f)
	) name928 (
		_w55_,
		_w39_,
		_w93_,
		_w259_,
		_w962_
	);
	LUT4 #(
		.INIT('h153f)
	) name929 (
		_w67_,
		_w47_,
		_w43_,
		_w201_,
		_w963_
	);
	LUT4 #(
		.INIT('h153f)
	) name930 (
		_w47_,
		_w72_,
		_w46_,
		_w184_,
		_w964_
	);
	LUT3 #(
		.INIT('h80)
	) name931 (
		_w963_,
		_w964_,
		_w962_,
		_w965_
	);
	LUT4 #(
		.INIT('h0777)
	) name932 (
		_w85_,
		_w39_,
		_w46_,
		_w378_,
		_w966_
	);
	LUT4 #(
		.INIT('h8000)
	) name933 (
		_w772_,
		_w892_,
		_w857_,
		_w966_,
		_w967_
	);
	LUT4 #(
		.INIT('h8000)
	) name934 (
		_w965_,
		_w967_,
		_w959_,
		_w961_,
		_w968_
	);
	LUT4 #(
		.INIT('h135f)
	) name935 (
		_w52_,
		_w56_,
		_w419_,
		_w378_,
		_w969_
	);
	LUT2 #(
		.INIT('h4)
	) name936 (
		_w202_,
		_w969_,
		_w970_
	);
	LUT4 #(
		.INIT('h0777)
	) name937 (
		_w106_,
		_w56_,
		_w50_,
		_w378_,
		_w971_
	);
	LUT3 #(
		.INIT('h37)
	) name938 (
		_w106_,
		_w41_,
		_w378_,
		_w972_
	);
	LUT4 #(
		.INIT('h4000)
	) name939 (
		_w186_,
		_w675_,
		_w971_,
		_w972_,
		_w973_
	);
	LUT4 #(
		.INIT('h135f)
	) name940 (
		_w78_,
		_w41_,
		_w44_,
		_w201_,
		_w974_
	);
	LUT4 #(
		.INIT('h153f)
	) name941 (
		_w41_,
		_w43_,
		_w44_,
		_w430_,
		_w975_
	);
	LUT4 #(
		.INIT('h135f)
	) name942 (
		_w59_,
		_w110_,
		_w236_,
		_w158_,
		_w976_
	);
	LUT3 #(
		.INIT('h80)
	) name943 (
		_w975_,
		_w976_,
		_w974_,
		_w977_
	);
	LUT4 #(
		.INIT('h153f)
	) name944 (
		_w55_,
		_w43_,
		_w65_,
		_w184_,
		_w978_
	);
	LUT4 #(
		.INIT('h153f)
	) name945 (
		_w56_,
		_w47_,
		_w72_,
		_w43_,
		_w979_
	);
	LUT4 #(
		.INIT('h0777)
	) name946 (
		_w106_,
		_w47_,
		_w46_,
		_w184_,
		_w980_
	);
	LUT4 #(
		.INIT('h8000)
	) name947 (
		_w924_,
		_w978_,
		_w979_,
		_w980_,
		_w981_
	);
	LUT4 #(
		.INIT('h8000)
	) name948 (
		_w970_,
		_w977_,
		_w981_,
		_w973_,
		_w982_
	);
	LUT4 #(
		.INIT('h8000)
	) name949 (
		_w968_,
		_w982_,
		_w939_,
		_w955_,
		_w983_
	);
	LUT2 #(
		.INIT('h8)
	) name950 (
		_w763_,
		_w983_,
		_w984_
	);
	LUT4 #(
		.INIT('h153f)
	) name951 (
		_w106_,
		_w50_,
		_w43_,
		_w44_,
		_w985_
	);
	LUT4 #(
		.INIT('h0777)
	) name952 (
		_w106_,
		_w52_,
		_w44_,
		_w259_,
		_w986_
	);
	LUT3 #(
		.INIT('h40)
	) name953 (
		_w268_,
		_w986_,
		_w985_,
		_w987_
	);
	LUT4 #(
		.INIT('h135f)
	) name954 (
		_w90_,
		_w44_,
		_w259_,
		_w430_,
		_w988_
	);
	LUT2 #(
		.INIT('h4)
	) name955 (
		_w468_,
		_w988_,
		_w989_
	);
	LUT4 #(
		.INIT('h0777)
	) name956 (
		_w41_,
		_w39_,
		_w65_,
		_w259_,
		_w990_
	);
	LUT3 #(
		.INIT('h57)
	) name957 (
		_w38_,
		_w78_,
		_w419_,
		_w991_
	);
	LUT4 #(
		.INIT('h135f)
	) name958 (
		_w67_,
		_w44_,
		_w184_,
		_w419_,
		_w992_
	);
	LUT4 #(
		.INIT('h8000)
	) name959 (
		_w807_,
		_w990_,
		_w991_,
		_w992_,
		_w993_
	);
	LUT3 #(
		.INIT('h80)
	) name960 (
		_w987_,
		_w989_,
		_w993_,
		_w994_
	);
	LUT4 #(
		.INIT('h153f)
	) name961 (
		_w55_,
		_w56_,
		_w176_,
		_w430_,
		_w995_
	);
	LUT2 #(
		.INIT('h8)
	) name962 (
		_w116_,
		_w995_,
		_w996_
	);
	LUT4 #(
		.INIT('h135f)
	) name963 (
		_w122_,
		_w50_,
		_w44_,
		_w184_,
		_w997_
	);
	LUT4 #(
		.INIT('h135f)
	) name964 (
		_w38_,
		_w106_,
		_w39_,
		_w93_,
		_w998_
	);
	LUT4 #(
		.INIT('h8000)
	) name965 (
		_w846_,
		_w847_,
		_w997_,
		_w998_,
		_w999_
	);
	LUT2 #(
		.INIT('h8)
	) name966 (
		_w996_,
		_w999_,
		_w1000_
	);
	LUT4 #(
		.INIT('h153f)
	) name967 (
		_w47_,
		_w43_,
		_w65_,
		_w184_,
		_w1001_
	);
	LUT4 #(
		.INIT('h4000)
	) name968 (
		_w369_,
		_w609_,
		_w636_,
		_w1001_,
		_w1002_
	);
	LUT4 #(
		.INIT('h0777)
	) name969 (
		_w106_,
		_w110_,
		_w72_,
		_w65_,
		_w1003_
	);
	LUT4 #(
		.INIT('h135f)
	) name970 (
		_w85_,
		_w59_,
		_w78_,
		_w166_,
		_w1004_
	);
	LUT3 #(
		.INIT('h80)
	) name971 (
		_w820_,
		_w1004_,
		_w1003_,
		_w1005_
	);
	LUT4 #(
		.INIT('h0777)
	) name972 (
		_w38_,
		_w106_,
		_w59_,
		_w158_,
		_w1006_
	);
	LUT4 #(
		.INIT('h0800)
	) name973 (
		_w252_,
		_w496_,
		_w445_,
		_w1006_,
		_w1007_
	);
	LUT3 #(
		.INIT('h80)
	) name974 (
		_w1002_,
		_w1005_,
		_w1007_,
		_w1008_
	);
	LUT3 #(
		.INIT('h80)
	) name975 (
		_w994_,
		_w1000_,
		_w1008_,
		_w1009_
	);
	LUT4 #(
		.INIT('h0777)
	) name976 (
		_w122_,
		_w52_,
		_w90_,
		_w72_,
		_w1010_
	);
	LUT2 #(
		.INIT('h8)
	) name977 (
		_w126_,
		_w1010_,
		_w1011_
	);
	LUT4 #(
		.INIT('h135f)
	) name978 (
		_w106_,
		_w85_,
		_w59_,
		_w166_,
		_w1012_
	);
	LUT4 #(
		.INIT('h153f)
	) name979 (
		_w90_,
		_w46_,
		_w184_,
		_w419_,
		_w1013_
	);
	LUT4 #(
		.INIT('h135f)
	) name980 (
		_w38_,
		_w67_,
		_w236_,
		_w378_,
		_w1014_
	);
	LUT4 #(
		.INIT('h8000)
	) name981 (
		_w950_,
		_w1012_,
		_w1013_,
		_w1014_,
		_w1015_
	);
	LUT4 #(
		.INIT('h153f)
	) name982 (
		_w59_,
		_w78_,
		_w46_,
		_w201_,
		_w1016_
	);
	LUT4 #(
		.INIT('h8000)
	) name983 (
		_w48_,
		_w828_,
		_w906_,
		_w1016_,
		_w1017_
	);
	LUT3 #(
		.INIT('h80)
	) name984 (
		_w1011_,
		_w1015_,
		_w1017_,
		_w1018_
	);
	LUT4 #(
		.INIT('h153f)
	) name985 (
		_w90_,
		_w93_,
		_w184_,
		_w166_,
		_w1019_
	);
	LUT3 #(
		.INIT('h40)
	) name986 (
		_w285_,
		_w555_,
		_w1019_,
		_w1020_
	);
	LUT3 #(
		.INIT('h1f)
	) name987 (
		_w110_,
		_w90_,
		_w184_,
		_w1021_
	);
	LUT2 #(
		.INIT('h4)
	) name988 (
		_w437_,
		_w1021_,
		_w1022_
	);
	LUT4 #(
		.INIT('h153f)
	) name989 (
		_w85_,
		_w41_,
		_w236_,
		_w259_,
		_w1023_
	);
	LUT4 #(
		.INIT('h0800)
	) name990 (
		_w68_,
		_w70_,
		_w353_,
		_w1023_,
		_w1024_
	);
	LUT4 #(
		.INIT('h8000)
	) name991 (
		_w540_,
		_w1022_,
		_w1020_,
		_w1024_,
		_w1025_
	);
	LUT4 #(
		.INIT('h0777)
	) name992 (
		_w85_,
		_w39_,
		_w65_,
		_w430_,
		_w1026_
	);
	LUT4 #(
		.INIT('h135f)
	) name993 (
		_w55_,
		_w65_,
		_w184_,
		_w378_,
		_w1027_
	);
	LUT2 #(
		.INIT('h8)
	) name994 (
		_w1026_,
		_w1027_,
		_w1028_
	);
	LUT4 #(
		.INIT('h135f)
	) name995 (
		_w59_,
		_w41_,
		_w39_,
		_w259_,
		_w1029_
	);
	LUT2 #(
		.INIT('h4)
	) name996 (
		_w400_,
		_w1029_,
		_w1030_
	);
	LUT4 #(
		.INIT('h0400)
	) name997 (
		_w325_,
		_w361_,
		_w400_,
		_w1029_,
		_w1031_
	);
	LUT3 #(
		.INIT('h10)
	) name998 (
		_w147_,
		_w182_,
		_w806_,
		_w1032_
	);
	LUT3 #(
		.INIT('h57)
	) name999 (
		_w93_,
		_w158_,
		_w176_,
		_w1033_
	);
	LUT4 #(
		.INIT('h4000)
	) name1000 (
		_w380_,
		_w781_,
		_w865_,
		_w1033_,
		_w1034_
	);
	LUT4 #(
		.INIT('h8000)
	) name1001 (
		_w1032_,
		_w1028_,
		_w1034_,
		_w1031_,
		_w1035_
	);
	LUT4 #(
		.INIT('h153f)
	) name1002 (
		_w52_,
		_w59_,
		_w184_,
		_w201_,
		_w1036_
	);
	LUT4 #(
		.INIT('h135f)
	) name1003 (
		_w47_,
		_w46_,
		_w236_,
		_w166_,
		_w1037_
	);
	LUT4 #(
		.INIT('h8000)
	) name1004 (
		_w582_,
		_w656_,
		_w1036_,
		_w1037_,
		_w1038_
	);
	LUT3 #(
		.INIT('h1f)
	) name1005 (
		_w38_,
		_w44_,
		_w184_,
		_w1039_
	);
	LUT3 #(
		.INIT('h37)
	) name1006 (
		_w38_,
		_w72_,
		_w46_,
		_w1040_
	);
	LUT4 #(
		.INIT('h153f)
	) name1007 (
		_w85_,
		_w67_,
		_w158_,
		_w430_,
		_w1041_
	);
	LUT4 #(
		.INIT('h4000)
	) name1008 (
		_w271_,
		_w1039_,
		_w1040_,
		_w1041_,
		_w1042_
	);
	LUT4 #(
		.INIT('h135f)
	) name1009 (
		_w52_,
		_w56_,
		_w259_,
		_w419_,
		_w1043_
	);
	LUT2 #(
		.INIT('h4)
	) name1010 (
		_w294_,
		_w1043_,
		_w1044_
	);
	LUT4 #(
		.INIT('h153f)
	) name1011 (
		_w59_,
		_w41_,
		_w166_,
		_w259_,
		_w1045_
	);
	LUT4 #(
		.INIT('h135f)
	) name1012 (
		_w106_,
		_w85_,
		_w56_,
		_w184_,
		_w1046_
	);
	LUT4 #(
		.INIT('h153f)
	) name1013 (
		_w52_,
		_w93_,
		_w259_,
		_w176_,
		_w1047_
	);
	LUT3 #(
		.INIT('h80)
	) name1014 (
		_w1046_,
		_w1047_,
		_w1045_,
		_w1048_
	);
	LUT4 #(
		.INIT('h8000)
	) name1015 (
		_w1038_,
		_w1042_,
		_w1044_,
		_w1048_,
		_w1049_
	);
	LUT4 #(
		.INIT('h8000)
	) name1016 (
		_w1018_,
		_w1025_,
		_w1035_,
		_w1049_,
		_w1050_
	);
	LUT2 #(
		.INIT('h8)
	) name1017 (
		_w1009_,
		_w1050_,
		_w1051_
	);
	LUT4 #(
		.INIT('h0777)
	) name1018 (
		_w763_,
		_w983_,
		_w1009_,
		_w1050_,
		_w1052_
	);
	LUT4 #(
		.INIT('h153f)
	) name1019 (
		_w55_,
		_w110_,
		_w184_,
		_w236_,
		_w1053_
	);
	LUT2 #(
		.INIT('h4)
	) name1020 (
		_w354_,
		_w1053_,
		_w1054_
	);
	LUT4 #(
		.INIT('h135f)
	) name1021 (
		_w106_,
		_w41_,
		_w46_,
		_w184_,
		_w1055_
	);
	LUT4 #(
		.INIT('h8000)
	) name1022 (
		_w148_,
		_w681_,
		_w1003_,
		_w1055_,
		_w1056_
	);
	LUT2 #(
		.INIT('h8)
	) name1023 (
		_w1054_,
		_w1056_,
		_w1057_
	);
	LUT4 #(
		.INIT('h135f)
	) name1024 (
		_w47_,
		_w44_,
		_w184_,
		_w419_,
		_w1058_
	);
	LUT4 #(
		.INIT('h135f)
	) name1025 (
		_w106_,
		_w55_,
		_w67_,
		_w166_,
		_w1059_
	);
	LUT4 #(
		.INIT('h135f)
	) name1026 (
		_w52_,
		_w44_,
		_w378_,
		_w430_,
		_w1060_
	);
	LUT4 #(
		.INIT('h135f)
	) name1027 (
		_w122_,
		_w67_,
		_w41_,
		_w43_,
		_w1061_
	);
	LUT4 #(
		.INIT('h8000)
	) name1028 (
		_w1058_,
		_w1060_,
		_w1061_,
		_w1059_,
		_w1062_
	);
	LUT4 #(
		.INIT('h135f)
	) name1029 (
		_w85_,
		_w110_,
		_w72_,
		_w39_,
		_w1063_
	);
	LUT4 #(
		.INIT('h153f)
	) name1030 (
		_w44_,
		_w46_,
		_w236_,
		_w259_,
		_w1064_
	);
	LUT3 #(
		.INIT('h40)
	) name1031 (
		_w393_,
		_w1063_,
		_w1064_,
		_w1065_
	);
	LUT4 #(
		.INIT('h135f)
	) name1032 (
		_w85_,
		_w44_,
		_w201_,
		_w176_,
		_w1066_
	);
	LUT4 #(
		.INIT('h153f)
	) name1033 (
		_w110_,
		_w72_,
		_w93_,
		_w430_,
		_w1067_
	);
	LUT3 #(
		.INIT('h57)
	) name1034 (
		_w110_,
		_w78_,
		_w259_,
		_w1068_
	);
	LUT3 #(
		.INIT('h80)
	) name1035 (
		_w1067_,
		_w1068_,
		_w1066_,
		_w1069_
	);
	LUT3 #(
		.INIT('h80)
	) name1036 (
		_w1065_,
		_w1062_,
		_w1069_,
		_w1070_
	);
	LUT2 #(
		.INIT('h8)
	) name1037 (
		_w1057_,
		_w1070_,
		_w1071_
	);
	LUT4 #(
		.INIT('h135f)
	) name1038 (
		_w39_,
		_w93_,
		_w44_,
		_w419_,
		_w1072_
	);
	LUT2 #(
		.INIT('h4)
	) name1039 (
		_w444_,
		_w1072_,
		_w1073_
	);
	LUT4 #(
		.INIT('h0777)
	) name1040 (
		_w78_,
		_w41_,
		_w46_,
		_w184_,
		_w1074_
	);
	LUT4 #(
		.INIT('h0777)
	) name1041 (
		_w41_,
		_w72_,
		_w43_,
		_w46_,
		_w1075_
	);
	LUT3 #(
		.INIT('h80)
	) name1042 (
		_w381_,
		_w1075_,
		_w1074_,
		_w1076_
	);
	LUT2 #(
		.INIT('h8)
	) name1043 (
		_w1073_,
		_w1076_,
		_w1077_
	);
	LUT4 #(
		.INIT('h153f)
	) name1044 (
		_w50_,
		_w65_,
		_w184_,
		_w236_,
		_w1078_
	);
	LUT4 #(
		.INIT('h153f)
	) name1045 (
		_w47_,
		_w93_,
		_w166_,
		_w378_,
		_w1079_
	);
	LUT4 #(
		.INIT('h135f)
	) name1046 (
		_w38_,
		_w65_,
		_w201_,
		_w166_,
		_w1080_
	);
	LUT3 #(
		.INIT('h80)
	) name1047 (
		_w1079_,
		_w1080_,
		_w1078_,
		_w1081_
	);
	LUT4 #(
		.INIT('h153f)
	) name1048 (
		_w38_,
		_w52_,
		_w236_,
		_w158_,
		_w1082_
	);
	LUT4 #(
		.INIT('h8000)
	) name1049 (
		_w479_,
		_w604_,
		_w566_,
		_w1082_,
		_w1083_
	);
	LUT4 #(
		.INIT('h153f)
	) name1050 (
		_w56_,
		_w39_,
		_w46_,
		_w166_,
		_w1084_
	);
	LUT4 #(
		.INIT('h2000)
	) name1051 (
		_w204_,
		_w457_,
		_w908_,
		_w1084_,
		_w1085_
	);
	LUT3 #(
		.INIT('h80)
	) name1052 (
		_w1081_,
		_w1083_,
		_w1085_,
		_w1086_
	);
	LUT4 #(
		.INIT('h153f)
	) name1053 (
		_w52_,
		_w56_,
		_w72_,
		_w201_,
		_w1087_
	);
	LUT4 #(
		.INIT('h153f)
	) name1054 (
		_w50_,
		_w93_,
		_w176_,
		_w430_,
		_w1088_
	);
	LUT4 #(
		.INIT('h0777)
	) name1055 (
		_w55_,
		_w78_,
		_w50_,
		_w201_,
		_w1089_
	);
	LUT4 #(
		.INIT('h8000)
	) name1056 (
		_w802_,
		_w1089_,
		_w1087_,
		_w1088_,
		_w1090_
	);
	LUT4 #(
		.INIT('h153f)
	) name1057 (
		_w110_,
		_w67_,
		_w78_,
		_w236_,
		_w1091_
	);
	LUT4 #(
		.INIT('h135f)
	) name1058 (
		_w38_,
		_w59_,
		_w166_,
		_w378_,
		_w1092_
	);
	LUT4 #(
		.INIT('h8000)
	) name1059 (
		_w843_,
		_w940_,
		_w1091_,
		_w1092_,
		_w1093_
	);
	LUT4 #(
		.INIT('h135f)
	) name1060 (
		_w90_,
		_w46_,
		_w166_,
		_w158_,
		_w1094_
	);
	LUT4 #(
		.INIT('h2000)
	) name1061 (
		_w54_,
		_w177_,
		_w809_,
		_w1094_,
		_w1095_
	);
	LUT3 #(
		.INIT('h80)
	) name1062 (
		_w1090_,
		_w1093_,
		_w1095_,
		_w1096_
	);
	LUT4 #(
		.INIT('h0777)
	) name1063 (
		_w122_,
		_w59_,
		_w56_,
		_w236_,
		_w1097_
	);
	LUT2 #(
		.INIT('h4)
	) name1064 (
		_w310_,
		_w1097_,
		_w1098_
	);
	LUT4 #(
		.INIT('h153f)
	) name1065 (
		_w52_,
		_w59_,
		_w78_,
		_w419_,
		_w1099_
	);
	LUT4 #(
		.INIT('h4000)
	) name1066 (
		_w295_,
		_w408_,
		_w951_,
		_w1099_,
		_w1100_
	);
	LUT4 #(
		.INIT('h8000)
	) name1067 (
		_w782_,
		_w786_,
		_w1098_,
		_w1100_,
		_w1101_
	);
	LUT4 #(
		.INIT('h8000)
	) name1068 (
		_w1077_,
		_w1086_,
		_w1096_,
		_w1101_,
		_w1102_
	);
	LUT2 #(
		.INIT('h8)
	) name1069 (
		_w1071_,
		_w1102_,
		_w1103_
	);
	LUT4 #(
		.INIT('h135f)
	) name1070 (
		_w39_,
		_w43_,
		_w65_,
		_w44_,
		_w1104_
	);
	LUT3 #(
		.INIT('h40)
	) name1071 (
		_w325_,
		_w361_,
		_w1104_,
		_w1105_
	);
	LUT4 #(
		.INIT('h135f)
	) name1072 (
		_w67_,
		_w44_,
		_w184_,
		_w236_,
		_w1106_
	);
	LUT3 #(
		.INIT('h40)
	) name1073 (
		_w363_,
		_w931_,
		_w1106_,
		_w1107_
	);
	LUT4 #(
		.INIT('h0777)
	) name1074 (
		_w122_,
		_w85_,
		_w90_,
		_w259_,
		_w1108_
	);
	LUT4 #(
		.INIT('h153f)
	) name1075 (
		_w38_,
		_w43_,
		_w93_,
		_w430_,
		_w1109_
	);
	LUT3 #(
		.INIT('h80)
	) name1076 (
		_w302_,
		_w1108_,
		_w1109_,
		_w1110_
	);
	LUT3 #(
		.INIT('h80)
	) name1077 (
		_w1107_,
		_w1110_,
		_w1105_,
		_w1111_
	);
	LUT4 #(
		.INIT('h0777)
	) name1078 (
		_w38_,
		_w122_,
		_w93_,
		_w176_,
		_w1112_
	);
	LUT4 #(
		.INIT('h135f)
	) name1079 (
		_w122_,
		_w55_,
		_w59_,
		_w166_,
		_w1113_
	);
	LUT3 #(
		.INIT('h37)
	) name1080 (
		_w106_,
		_w55_,
		_w72_,
		_w1114_
	);
	LUT4 #(
		.INIT('h8000)
	) name1081 (
		_w42_,
		_w1112_,
		_w1113_,
		_w1114_,
		_w1115_
	);
	LUT4 #(
		.INIT('h135f)
	) name1082 (
		_w110_,
		_w72_,
		_w39_,
		_w44_,
		_w1116_
	);
	LUT2 #(
		.INIT('h4)
	) name1083 (
		_w276_,
		_w1116_,
		_w1117_
	);
	LUT3 #(
		.INIT('h1f)
	) name1084 (
		_w90_,
		_w46_,
		_w184_,
		_w1118_
	);
	LUT4 #(
		.INIT('h153f)
	) name1085 (
		_w55_,
		_w52_,
		_w236_,
		_w378_,
		_w1119_
	);
	LUT4 #(
		.INIT('h4000)
	) name1086 (
		_w276_,
		_w1116_,
		_w1118_,
		_w1119_,
		_w1120_
	);
	LUT2 #(
		.INIT('h8)
	) name1087 (
		_w1115_,
		_w1120_,
		_w1121_
	);
	LUT4 #(
		.INIT('h153f)
	) name1088 (
		_w85_,
		_w93_,
		_w201_,
		_w158_,
		_w1122_
	);
	LUT2 #(
		.INIT('h4)
	) name1089 (
		_w451_,
		_w1122_,
		_w1123_
	);
	LUT4 #(
		.INIT('h135f)
	) name1090 (
		_w52_,
		_w59_,
		_w184_,
		_w201_,
		_w1124_
	);
	LUT4 #(
		.INIT('h153f)
	) name1091 (
		_w90_,
		_w41_,
		_w176_,
		_w378_,
		_w1125_
	);
	LUT4 #(
		.INIT('h0777)
	) name1092 (
		_w122_,
		_w90_,
		_w41_,
		_w43_,
		_w1126_
	);
	LUT4 #(
		.INIT('h153f)
	) name1093 (
		_w47_,
		_w50_,
		_w184_,
		_w259_,
		_w1127_
	);
	LUT4 #(
		.INIT('h8000)
	) name1094 (
		_w1124_,
		_w1126_,
		_w1127_,
		_w1125_,
		_w1128_
	);
	LUT2 #(
		.INIT('h8)
	) name1095 (
		_w1123_,
		_w1128_,
		_w1129_
	);
	LUT4 #(
		.INIT('h135f)
	) name1096 (
		_w78_,
		_w47_,
		_w50_,
		_w158_,
		_w1130_
	);
	LUT3 #(
		.INIT('h37)
	) name1097 (
		_w59_,
		_w78_,
		_w93_,
		_w1131_
	);
	LUT4 #(
		.INIT('h135f)
	) name1098 (
		_w106_,
		_w65_,
		_w44_,
		_w166_,
		_w1132_
	);
	LUT4 #(
		.INIT('h8000)
	) name1099 (
		_w978_,
		_w1131_,
		_w1132_,
		_w1130_,
		_w1133_
	);
	LUT4 #(
		.INIT('h0200)
	) name1100 (
		_w81_,
		_w193_,
		_w314_,
		_w823_,
		_w1134_
	);
	LUT4 #(
		.INIT('h8000)
	) name1101 (
		_w1123_,
		_w1128_,
		_w1133_,
		_w1134_,
		_w1135_
	);
	LUT3 #(
		.INIT('h80)
	) name1102 (
		_w1121_,
		_w1111_,
		_w1135_,
		_w1136_
	);
	LUT4 #(
		.INIT('h135f)
	) name1103 (
		_w93_,
		_w44_,
		_w419_,
		_w378_,
		_w1137_
	);
	LUT3 #(
		.INIT('h1f)
	) name1104 (
		_w110_,
		_w44_,
		_w201_,
		_w1138_
	);
	LUT4 #(
		.INIT('h135f)
	) name1105 (
		_w85_,
		_w110_,
		_w43_,
		_w158_,
		_w1139_
	);
	LUT3 #(
		.INIT('h80)
	) name1106 (
		_w1138_,
		_w1139_,
		_w1137_,
		_w1140_
	);
	LUT4 #(
		.INIT('h135f)
	) name1107 (
		_w56_,
		_w41_,
		_w39_,
		_w236_,
		_w1141_
	);
	LUT2 #(
		.INIT('h4)
	) name1108 (
		_w383_,
		_w1141_,
		_w1142_
	);
	LUT4 #(
		.INIT('h135f)
	) name1109 (
		_w85_,
		_w59_,
		_w72_,
		_w419_,
		_w1143_
	);
	LUT4 #(
		.INIT('h153f)
	) name1110 (
		_w106_,
		_w52_,
		_w78_,
		_w46_,
		_w1144_
	);
	LUT4 #(
		.INIT('h4000)
	) name1111 (
		_w64_,
		_w678_,
		_w1143_,
		_w1144_,
		_w1145_
	);
	LUT3 #(
		.INIT('h80)
	) name1112 (
		_w1142_,
		_w1140_,
		_w1145_,
		_w1146_
	);
	LUT4 #(
		.INIT('h135f)
	) name1113 (
		_w122_,
		_w55_,
		_w44_,
		_w259_,
		_w1147_
	);
	LUT4 #(
		.INIT('h135f)
	) name1114 (
		_w52_,
		_w59_,
		_w259_,
		_w176_,
		_w1148_
	);
	LUT2 #(
		.INIT('h8)
	) name1115 (
		_w1147_,
		_w1148_,
		_w1149_
	);
	LUT4 #(
		.INIT('h153f)
	) name1116 (
		_w38_,
		_w39_,
		_w44_,
		_w236_,
		_w1150_
	);
	LUT4 #(
		.INIT('h135f)
	) name1117 (
		_w38_,
		_w65_,
		_w419_,
		_w378_,
		_w1151_
	);
	LUT4 #(
		.INIT('h4000)
	) name1118 (
		_w412_,
		_w855_,
		_w1150_,
		_w1151_,
		_w1152_
	);
	LUT4 #(
		.INIT('h153f)
	) name1119 (
		_w52_,
		_w65_,
		_w201_,
		_w158_,
		_w1153_
	);
	LUT4 #(
		.INIT('h135f)
	) name1120 (
		_w56_,
		_w50_,
		_w236_,
		_w259_,
		_w1154_
	);
	LUT3 #(
		.INIT('h80)
	) name1121 (
		_w115_,
		_w1154_,
		_w1153_,
		_w1155_
	);
	LUT3 #(
		.INIT('h1f)
	) name1122 (
		_w90_,
		_w41_,
		_w166_,
		_w1156_
	);
	LUT3 #(
		.INIT('h1f)
	) name1123 (
		_w85_,
		_w52_,
		_w419_,
		_w1157_
	);
	LUT4 #(
		.INIT('h153f)
	) name1124 (
		_w90_,
		_w46_,
		_w158_,
		_w419_,
		_w1158_
	);
	LUT4 #(
		.INIT('h8000)
	) name1125 (
		_w1004_,
		_w1156_,
		_w1157_,
		_w1158_,
		_w1159_
	);
	LUT4 #(
		.INIT('h8000)
	) name1126 (
		_w1149_,
		_w1155_,
		_w1159_,
		_w1152_,
		_w1160_
	);
	LUT3 #(
		.INIT('h57)
	) name1127 (
		_w59_,
		_w43_,
		_w259_,
		_w1161_
	);
	LUT4 #(
		.INIT('h135f)
	) name1128 (
		_w106_,
		_w110_,
		_w93_,
		_w378_,
		_w1162_
	);
	LUT2 #(
		.INIT('h8)
	) name1129 (
		_w1161_,
		_w1162_,
		_w1163_
	);
	LUT4 #(
		.INIT('h135f)
	) name1130 (
		_w52_,
		_w56_,
		_w72_,
		_w176_,
		_w1164_
	);
	LUT4 #(
		.INIT('h153f)
	) name1131 (
		_w106_,
		_w90_,
		_w43_,
		_w65_,
		_w1165_
	);
	LUT4 #(
		.INIT('h135f)
	) name1132 (
		_w47_,
		_w50_,
		_w201_,
		_w158_,
		_w1166_
	);
	LUT4 #(
		.INIT('h8000)
	) name1133 (
		_w757_,
		_w1164_,
		_w1165_,
		_w1166_,
		_w1167_
	);
	LUT4 #(
		.INIT('h153f)
	) name1134 (
		_w65_,
		_w46_,
		_w201_,
		_w430_,
		_w1168_
	);
	LUT4 #(
		.INIT('h153f)
	) name1135 (
		_w52_,
		_w65_,
		_w236_,
		_w378_,
		_w1169_
	);
	LUT3 #(
		.INIT('h40)
	) name1136 (
		_w477_,
		_w1169_,
		_w1168_,
		_w1170_
	);
	LUT3 #(
		.INIT('h40)
	) name1137 (
		_w435_,
		_w937_,
		_w1067_,
		_w1171_
	);
	LUT4 #(
		.INIT('h8000)
	) name1138 (
		_w1170_,
		_w1171_,
		_w1163_,
		_w1167_,
		_w1172_
	);
	LUT4 #(
		.INIT('h0777)
	) name1139 (
		_w55_,
		_w43_,
		_w46_,
		_w236_,
		_w1173_
	);
	LUT4 #(
		.INIT('h153f)
	) name1140 (
		_w122_,
		_w55_,
		_w39_,
		_w93_,
		_w1174_
	);
	LUT4 #(
		.INIT('h8000)
	) name1141 (
		_w1036_,
		_w1084_,
		_w1173_,
		_w1174_,
		_w1175_
	);
	LUT4 #(
		.INIT('h153f)
	) name1142 (
		_w85_,
		_w41_,
		_w72_,
		_w39_,
		_w1176_
	);
	LUT4 #(
		.INIT('h135f)
	) name1143 (
		_w106_,
		_w52_,
		_w110_,
		_w176_,
		_w1177_
	);
	LUT4 #(
		.INIT('h8000)
	) name1144 (
		_w713_,
		_w816_,
		_w1176_,
		_w1177_,
		_w1178_
	);
	LUT4 #(
		.INIT('h153f)
	) name1145 (
		_w90_,
		_w72_,
		_w65_,
		_w158_,
		_w1179_
	);
	LUT4 #(
		.INIT('h153f)
	) name1146 (
		_w38_,
		_w90_,
		_w72_,
		_w184_,
		_w1180_
	);
	LUT4 #(
		.INIT('h0777)
	) name1147 (
		_w38_,
		_w106_,
		_w41_,
		_w158_,
		_w1181_
	);
	LUT4 #(
		.INIT('h135f)
	) name1148 (
		_w65_,
		_w46_,
		_w419_,
		_w378_,
		_w1182_
	);
	LUT4 #(
		.INIT('h8000)
	) name1149 (
		_w1179_,
		_w1180_,
		_w1181_,
		_w1182_,
		_w1183_
	);
	LUT4 #(
		.INIT('h153f)
	) name1150 (
		_w110_,
		_w78_,
		_w44_,
		_w236_,
		_w1184_
	);
	LUT4 #(
		.INIT('h4000)
	) name1151 (
		_w161_,
		_w639_,
		_w711_,
		_w1184_,
		_w1185_
	);
	LUT4 #(
		.INIT('h8000)
	) name1152 (
		_w1175_,
		_w1178_,
		_w1183_,
		_w1185_,
		_w1186_
	);
	LUT4 #(
		.INIT('h8000)
	) name1153 (
		_w1146_,
		_w1160_,
		_w1172_,
		_w1186_,
		_w1187_
	);
	LUT2 #(
		.INIT('h8)
	) name1154 (
		_w1136_,
		_w1187_,
		_w1188_
	);
	LUT4 #(
		.INIT('h0777)
	) name1155 (
		_w1071_,
		_w1102_,
		_w1136_,
		_w1187_,
		_w1189_
	);
	LUT4 #(
		.INIT('h135f)
	) name1156 (
		_w52_,
		_w90_,
		_w72_,
		_w259_,
		_w1190_
	);
	LUT4 #(
		.INIT('h0777)
	) name1157 (
		_w41_,
		_w43_,
		_w44_,
		_w430_,
		_w1191_
	);
	LUT4 #(
		.INIT('h135f)
	) name1158 (
		_w56_,
		_w46_,
		_w201_,
		_w259_,
		_w1192_
	);
	LUT4 #(
		.INIT('h8000)
	) name1159 (
		_w1012_,
		_w1190_,
		_w1191_,
		_w1192_,
		_w1193_
	);
	LUT4 #(
		.INIT('h2000)
	) name1160 (
		_w95_,
		_w295_,
		_w882_,
		_w913_,
		_w1194_
	);
	LUT3 #(
		.INIT('h80)
	) name1161 (
		_w1170_,
		_w1193_,
		_w1194_,
		_w1195_
	);
	LUT4 #(
		.INIT('h135f)
	) name1162 (
		_w41_,
		_w93_,
		_w176_,
		_w378_,
		_w1196_
	);
	LUT4 #(
		.INIT('h4000)
	) name1163 (
		_w363_,
		_w931_,
		_w1106_,
		_w1196_,
		_w1197_
	);
	LUT4 #(
		.INIT('h153f)
	) name1164 (
		_w55_,
		_w41_,
		_w72_,
		_w259_,
		_w1198_
	);
	LUT2 #(
		.INIT('h8)
	) name1165 (
		_w1037_,
		_w1198_,
		_w1199_
	);
	LUT3 #(
		.INIT('h20)
	) name1166 (
		_w126_,
		_w182_,
		_w806_,
		_w1200_
	);
	LUT4 #(
		.INIT('h8000)
	) name1167 (
		_w561_,
		_w565_,
		_w1199_,
		_w1200_,
		_w1201_
	);
	LUT3 #(
		.INIT('h80)
	) name1168 (
		_w1197_,
		_w1195_,
		_w1201_,
		_w1202_
	);
	LUT4 #(
		.INIT('h0777)
	) name1169 (
		_w59_,
		_w78_,
		_w47_,
		_w72_,
		_w1203_
	);
	LUT4 #(
		.INIT('h135f)
	) name1170 (
		_w41_,
		_w65_,
		_w184_,
		_w419_,
		_w1204_
	);
	LUT4 #(
		.INIT('h135f)
	) name1171 (
		_w67_,
		_w56_,
		_w158_,
		_w419_,
		_w1205_
	);
	LUT4 #(
		.INIT('h135f)
	) name1172 (
		_w67_,
		_w56_,
		_w166_,
		_w378_,
		_w1206_
	);
	LUT4 #(
		.INIT('h8000)
	) name1173 (
		_w1205_,
		_w1206_,
		_w1203_,
		_w1204_,
		_w1207_
	);
	LUT3 #(
		.INIT('h1f)
	) name1174 (
		_w85_,
		_w67_,
		_w176_,
		_w1208_
	);
	LUT4 #(
		.INIT('h135f)
	) name1175 (
		_w106_,
		_w67_,
		_w50_,
		_w430_,
		_w1209_
	);
	LUT2 #(
		.INIT('h8)
	) name1176 (
		_w1208_,
		_w1209_,
		_w1210_
	);
	LUT4 #(
		.INIT('h135f)
	) name1177 (
		_w106_,
		_w55_,
		_w65_,
		_w419_,
		_w1211_
	);
	LUT4 #(
		.INIT('h1000)
	) name1178 (
		_w294_,
		_w276_,
		_w746_,
		_w1211_,
		_w1212_
	);
	LUT3 #(
		.INIT('h80)
	) name1179 (
		_w1210_,
		_w1207_,
		_w1212_,
		_w1213_
	);
	LUT4 #(
		.INIT('h135f)
	) name1180 (
		_w106_,
		_w55_,
		_w85_,
		_w78_,
		_w1214_
	);
	LUT4 #(
		.INIT('h153f)
	) name1181 (
		_w52_,
		_w93_,
		_w184_,
		_w430_,
		_w1215_
	);
	LUT4 #(
		.INIT('h135f)
	) name1182 (
		_w55_,
		_w47_,
		_w236_,
		_w158_,
		_w1216_
	);
	LUT4 #(
		.INIT('h8000)
	) name1183 (
		_w594_,
		_w1215_,
		_w1216_,
		_w1214_,
		_w1217_
	);
	LUT4 #(
		.INIT('h153f)
	) name1184 (
		_w110_,
		_w43_,
		_w46_,
		_w166_,
		_w1218_
	);
	LUT3 #(
		.INIT('h40)
	) name1185 (
		_w393_,
		_w611_,
		_w1218_,
		_w1219_
	);
	LUT4 #(
		.INIT('h135f)
	) name1186 (
		_w72_,
		_w65_,
		_w44_,
		_w184_,
		_w1220_
	);
	LUT4 #(
		.INIT('h0777)
	) name1187 (
		_w52_,
		_w78_,
		_w41_,
		_w378_,
		_w1221_
	);
	LUT4 #(
		.INIT('h135f)
	) name1188 (
		_w47_,
		_w41_,
		_w43_,
		_w430_,
		_w1222_
	);
	LUT4 #(
		.INIT('h8000)
	) name1189 (
		_w770_,
		_w1221_,
		_w1222_,
		_w1220_,
		_w1223_
	);
	LUT3 #(
		.INIT('h80)
	) name1190 (
		_w1219_,
		_w1217_,
		_w1223_,
		_w1224_
	);
	LUT2 #(
		.INIT('h4)
	) name1191 (
		_w61_,
		_w370_,
		_w1225_
	);
	LUT4 #(
		.INIT('h0777)
	) name1192 (
		_w122_,
		_w50_,
		_w65_,
		_w176_,
		_w1226_
	);
	LUT3 #(
		.INIT('h40)
	) name1193 (
		_w186_,
		_w971_,
		_w1226_,
		_w1227_
	);
	LUT2 #(
		.INIT('h8)
	) name1194 (
		_w1225_,
		_w1227_,
		_w1228_
	);
	LUT4 #(
		.INIT('h135f)
	) name1195 (
		_w85_,
		_w90_,
		_w158_,
		_w378_,
		_w1229_
	);
	LUT4 #(
		.INIT('h4000)
	) name1196 (
		_w469_,
		_w597_,
		_w598_,
		_w1229_,
		_w1230_
	);
	LUT4 #(
		.INIT('h4000)
	) name1197 (
		_w339_,
		_w660_,
		_w997_,
		_w998_,
		_w1231_
	);
	LUT4 #(
		.INIT('h8000)
	) name1198 (
		_w1225_,
		_w1227_,
		_w1230_,
		_w1231_,
		_w1232_
	);
	LUT3 #(
		.INIT('h80)
	) name1199 (
		_w1213_,
		_w1224_,
		_w1232_,
		_w1233_
	);
	LUT2 #(
		.INIT('h8)
	) name1200 (
		_w1202_,
		_w1233_,
		_w1234_
	);
	LUT4 #(
		.INIT('h135f)
	) name1201 (
		_w38_,
		_w90_,
		_w166_,
		_w176_,
		_w1235_
	);
	LUT2 #(
		.INIT('h4)
	) name1202 (
		_w324_,
		_w1235_,
		_w1236_
	);
	LUT4 #(
		.INIT('h135f)
	) name1203 (
		_w85_,
		_w50_,
		_w43_,
		_w166_,
		_w1237_
	);
	LUT4 #(
		.INIT('h153f)
	) name1204 (
		_w38_,
		_w78_,
		_w65_,
		_w259_,
		_w1238_
	);
	LUT4 #(
		.INIT('h135f)
	) name1205 (
		_w55_,
		_w56_,
		_w201_,
		_w259_,
		_w1239_
	);
	LUT4 #(
		.INIT('h4000)
	) name1206 (
		_w365_,
		_w1238_,
		_w1237_,
		_w1239_,
		_w1240_
	);
	LUT2 #(
		.INIT('h8)
	) name1207 (
		_w1236_,
		_w1240_,
		_w1241_
	);
	LUT4 #(
		.INIT('h0777)
	) name1208 (
		_w67_,
		_w78_,
		_w72_,
		_w93_,
		_w1242_
	);
	LUT4 #(
		.INIT('h153f)
	) name1209 (
		_w38_,
		_w55_,
		_w184_,
		_w430_,
		_w1243_
	);
	LUT4 #(
		.INIT('h4000)
	) name1210 (
		_w247_,
		_w964_,
		_w1242_,
		_w1243_,
		_w1244_
	);
	LUT4 #(
		.INIT('h135f)
	) name1211 (
		_w52_,
		_w90_,
		_w158_,
		_w430_,
		_w1245_
	);
	LUT4 #(
		.INIT('h1000)
	) name1212 (
		_w74_,
		_w203_,
		_w1014_,
		_w1245_,
		_w1246_
	);
	LUT4 #(
		.INIT('h135f)
	) name1213 (
		_w52_,
		_w46_,
		_w201_,
		_w430_,
		_w1247_
	);
	LUT4 #(
		.INIT('h153f)
	) name1214 (
		_w85_,
		_w52_,
		_w39_,
		_w176_,
		_w1248_
	);
	LUT3 #(
		.INIT('h80)
	) name1215 (
		_w975_,
		_w1248_,
		_w1247_,
		_w1249_
	);
	LUT3 #(
		.INIT('h37)
	) name1216 (
		_w78_,
		_w41_,
		_w43_,
		_w1250_
	);
	LUT4 #(
		.INIT('h8000)
	) name1217 (
		_w305_,
		_w384_,
		_w893_,
		_w1250_,
		_w1251_
	);
	LUT4 #(
		.INIT('h8000)
	) name1218 (
		_w1249_,
		_w1251_,
		_w1244_,
		_w1246_,
		_w1252_
	);
	LUT2 #(
		.INIT('h8)
	) name1219 (
		_w1241_,
		_w1252_,
		_w1253_
	);
	LUT3 #(
		.INIT('h57)
	) name1220 (
		_w67_,
		_w236_,
		_w176_,
		_w1254_
	);
	LUT4 #(
		.INIT('h135f)
	) name1221 (
		_w65_,
		_w44_,
		_w176_,
		_w430_,
		_w1255_
	);
	LUT2 #(
		.INIT('h8)
	) name1222 (
		_w1254_,
		_w1255_,
		_w1256_
	);
	LUT4 #(
		.INIT('h0777)
	) name1223 (
		_w56_,
		_w39_,
		_w65_,
		_w184_,
		_w1257_
	);
	LUT4 #(
		.INIT('h0777)
	) name1224 (
		_w59_,
		_w39_,
		_w43_,
		_w46_,
		_w1258_
	);
	LUT4 #(
		.INIT('h153f)
	) name1225 (
		_w90_,
		_w47_,
		_w39_,
		_w201_,
		_w1259_
	);
	LUT3 #(
		.INIT('h80)
	) name1226 (
		_w1257_,
		_w1258_,
		_w1259_,
		_w1260_
	);
	LUT2 #(
		.INIT('h8)
	) name1227 (
		_w1256_,
		_w1260_,
		_w1261_
	);
	LUT4 #(
		.INIT('h0777)
	) name1228 (
		_w122_,
		_w50_,
		_w44_,
		_w419_,
		_w1262_
	);
	LUT3 #(
		.INIT('h40)
	) name1229 (
		_w471_,
		_w601_,
		_w1262_,
		_w1263_
	);
	LUT4 #(
		.INIT('h1000)
	) name1230 (
		_w271_,
		_w439_,
		_w832_,
		_w1039_,
		_w1264_
	);
	LUT4 #(
		.INIT('h135f)
	) name1231 (
		_w110_,
		_w41_,
		_w236_,
		_w378_,
		_w1265_
	);
	LUT4 #(
		.INIT('h135f)
	) name1232 (
		_w106_,
		_w59_,
		_w47_,
		_w166_,
		_w1266_
	);
	LUT3 #(
		.INIT('h40)
	) name1233 (
		_w325_,
		_w1265_,
		_w1266_,
		_w1267_
	);
	LUT4 #(
		.INIT('h153f)
	) name1234 (
		_w59_,
		_w47_,
		_w72_,
		_w158_,
		_w1268_
	);
	LUT3 #(
		.INIT('h57)
	) name1235 (
		_w50_,
		_w236_,
		_w176_,
		_w1269_
	);
	LUT4 #(
		.INIT('h8000)
	) name1236 (
		_w924_,
		_w909_,
		_w1269_,
		_w1268_,
		_w1270_
	);
	LUT4 #(
		.INIT('h8000)
	) name1237 (
		_w1267_,
		_w1270_,
		_w1263_,
		_w1264_,
		_w1271_
	);
	LUT2 #(
		.INIT('h8)
	) name1238 (
		_w1261_,
		_w1271_,
		_w1272_
	);
	LUT4 #(
		.INIT('h153f)
	) name1239 (
		_w38_,
		_w110_,
		_w166_,
		_w158_,
		_w1273_
	);
	LUT4 #(
		.INIT('h135f)
	) name1240 (
		_w78_,
		_w56_,
		_w44_,
		_w201_,
		_w1274_
	);
	LUT4 #(
		.INIT('h153f)
	) name1241 (
		_w85_,
		_w52_,
		_w419_,
		_w430_,
		_w1275_
	);
	LUT4 #(
		.INIT('h0777)
	) name1242 (
		_w122_,
		_w55_,
		_w56_,
		_w430_,
		_w1276_
	);
	LUT4 #(
		.INIT('h8000)
	) name1243 (
		_w1273_,
		_w1275_,
		_w1276_,
		_w1274_,
		_w1277_
	);
	LUT3 #(
		.INIT('h37)
	) name1244 (
		_w39_,
		_w65_,
		_w378_,
		_w1278_
	);
	LUT4 #(
		.INIT('h4000)
	) name1245 (
		_w380_,
		_w806_,
		_w794_,
		_w1278_,
		_w1279_
	);
	LUT4 #(
		.INIT('h153f)
	) name1246 (
		_w55_,
		_w90_,
		_w259_,
		_w176_,
		_w1280_
	);
	LUT4 #(
		.INIT('h135f)
	) name1247 (
		_w106_,
		_w93_,
		_w44_,
		_w176_,
		_w1281_
	);
	LUT3 #(
		.INIT('h80)
	) name1248 (
		_w1198_,
		_w1281_,
		_w1280_,
		_w1282_
	);
	LUT3 #(
		.INIT('h80)
	) name1249 (
		_w1279_,
		_w1277_,
		_w1282_,
		_w1283_
	);
	LUT4 #(
		.INIT('h153f)
	) name1250 (
		_w38_,
		_w52_,
		_w72_,
		_w43_,
		_w1284_
	);
	LUT4 #(
		.INIT('h0777)
	) name1251 (
		_w122_,
		_w56_,
		_w93_,
		_w184_,
		_w1285_
	);
	LUT2 #(
		.INIT('h8)
	) name1252 (
		_w1284_,
		_w1285_,
		_w1286_
	);
	LUT4 #(
		.INIT('h135f)
	) name1253 (
		_w78_,
		_w47_,
		_w93_,
		_w201_,
		_w1287_
	);
	LUT4 #(
		.INIT('h135f)
	) name1254 (
		_w59_,
		_w47_,
		_w72_,
		_w430_,
		_w1288_
	);
	LUT3 #(
		.INIT('h80)
	) name1255 (
		_w132_,
		_w1288_,
		_w1287_,
		_w1289_
	);
	LUT2 #(
		.INIT('h4)
	) name1256 (
		_w273_,
		_w348_,
		_w1290_
	);
	LUT4 #(
		.INIT('h135f)
	) name1257 (
		_w85_,
		_w46_,
		_w166_,
		_w419_,
		_w1291_
	);
	LUT4 #(
		.INIT('h4000)
	) name1258 (
		_w454_,
		_w662_,
		_w1084_,
		_w1291_,
		_w1292_
	);
	LUT4 #(
		.INIT('h8000)
	) name1259 (
		_w1290_,
		_w1286_,
		_w1289_,
		_w1292_,
		_w1293_
	);
	LUT4 #(
		.INIT('h8000)
	) name1260 (
		_w1261_,
		_w1271_,
		_w1283_,
		_w1293_,
		_w1294_
	);
	LUT2 #(
		.INIT('h8)
	) name1261 (
		_w1253_,
		_w1294_,
		_w1295_
	);
	LUT4 #(
		.INIT('h0777)
	) name1262 (
		_w1202_,
		_w1233_,
		_w1253_,
		_w1294_,
		_w1296_
	);
	LUT4 #(
		.INIT('h0777)
	) name1263 (
		_w85_,
		_w78_,
		_w41_,
		_w419_,
		_w1297_
	);
	LUT4 #(
		.INIT('h153f)
	) name1264 (
		_w90_,
		_w72_,
		_w50_,
		_w201_,
		_w1298_
	);
	LUT3 #(
		.INIT('h57)
	) name1265 (
		_w44_,
		_w236_,
		_w166_,
		_w1299_
	);
	LUT3 #(
		.INIT('h80)
	) name1266 (
		_w1297_,
		_w1298_,
		_w1299_,
		_w1300_
	);
	LUT4 #(
		.INIT('h153f)
	) name1267 (
		_w38_,
		_w106_,
		_w65_,
		_w176_,
		_w1301_
	);
	LUT2 #(
		.INIT('h8)
	) name1268 (
		_w112_,
		_w1301_,
		_w1302_
	);
	LUT4 #(
		.INIT('h153f)
	) name1269 (
		_w47_,
		_w93_,
		_w236_,
		_w419_,
		_w1303_
	);
	LUT4 #(
		.INIT('h135f)
	) name1270 (
		_w67_,
		_w50_,
		_w158_,
		_w430_,
		_w1304_
	);
	LUT4 #(
		.INIT('h153f)
	) name1271 (
		_w56_,
		_w65_,
		_w236_,
		_w430_,
		_w1305_
	);
	LUT4 #(
		.INIT('h4000)
	) name1272 (
		_w60_,
		_w1303_,
		_w1304_,
		_w1305_,
		_w1306_
	);
	LUT3 #(
		.INIT('h80)
	) name1273 (
		_w1302_,
		_w1300_,
		_w1306_,
		_w1307_
	);
	LUT4 #(
		.INIT('h135f)
	) name1274 (
		_w41_,
		_w50_,
		_w201_,
		_w176_,
		_w1308_
	);
	LUT2 #(
		.INIT('h4)
	) name1275 (
		_w347_,
		_w1308_,
		_w1309_
	);
	LUT4 #(
		.INIT('h153f)
	) name1276 (
		_w67_,
		_w50_,
		_w43_,
		_w259_,
		_w1310_
	);
	LUT4 #(
		.INIT('h153f)
	) name1277 (
		_w38_,
		_w90_,
		_w39_,
		_w184_,
		_w1311_
	);
	LUT3 #(
		.INIT('h40)
	) name1278 (
		_w268_,
		_w1310_,
		_w1311_,
		_w1312_
	);
	LUT2 #(
		.INIT('h8)
	) name1279 (
		_w1309_,
		_w1312_,
		_w1313_
	);
	LUT4 #(
		.INIT('h135f)
	) name1280 (
		_w106_,
		_w41_,
		_w46_,
		_w166_,
		_w1314_
	);
	LUT4 #(
		.INIT('h8000)
	) name1281 (
		_w148_,
		_w66_,
		_w611_,
		_w1314_,
		_w1315_
	);
	LUT4 #(
		.INIT('h0777)
	) name1282 (
		_w122_,
		_w85_,
		_w72_,
		_w46_,
		_w1316_
	);
	LUT2 #(
		.INIT('h4)
	) name1283 (
		_w212_,
		_w1316_,
		_w1317_
	);
	LUT4 #(
		.INIT('h135f)
	) name1284 (
		_w122_,
		_w56_,
		_w46_,
		_w176_,
		_w1318_
	);
	LUT4 #(
		.INIT('h153f)
	) name1285 (
		_w85_,
		_w78_,
		_w50_,
		_w378_,
		_w1319_
	);
	LUT4 #(
		.INIT('h4000)
	) name1286 (
		_w212_,
		_w1316_,
		_w1318_,
		_w1319_,
		_w1320_
	);
	LUT4 #(
		.INIT('h0777)
	) name1287 (
		_w106_,
		_w67_,
		_w47_,
		_w176_,
		_w1321_
	);
	LUT3 #(
		.INIT('h80)
	) name1288 (
		_w384_,
		_w1184_,
		_w1321_,
		_w1322_
	);
	LUT3 #(
		.INIT('h80)
	) name1289 (
		_w634_,
		_w1182_,
		_w1190_,
		_w1323_
	);
	LUT4 #(
		.INIT('h8000)
	) name1290 (
		_w1322_,
		_w1323_,
		_w1315_,
		_w1320_,
		_w1324_
	);
	LUT3 #(
		.INIT('h80)
	) name1291 (
		_w1313_,
		_w1307_,
		_w1324_,
		_w1325_
	);
	LUT4 #(
		.INIT('h0777)
	) name1292 (
		_w122_,
		_w110_,
		_w90_,
		_w43_,
		_w1326_
	);
	LUT3 #(
		.INIT('h40)
	) name1293 (
		_w435_,
		_w1147_,
		_w1326_,
		_w1327_
	);
	LUT4 #(
		.INIT('h0777)
	) name1294 (
		_w38_,
		_w106_,
		_w85_,
		_w201_,
		_w1328_
	);
	LUT4 #(
		.INIT('h0777)
	) name1295 (
		_w106_,
		_w85_,
		_w65_,
		_w184_,
		_w1329_
	);
	LUT4 #(
		.INIT('h135f)
	) name1296 (
		_w47_,
		_w93_,
		_w236_,
		_w259_,
		_w1330_
	);
	LUT4 #(
		.INIT('h4000)
	) name1297 (
		_w308_,
		_w1328_,
		_w1329_,
		_w1330_,
		_w1331_
	);
	LUT4 #(
		.INIT('h0777)
	) name1298 (
		_w122_,
		_w52_,
		_w47_,
		_w166_,
		_w1332_
	);
	LUT4 #(
		.INIT('h153f)
	) name1299 (
		_w38_,
		_w78_,
		_w47_,
		_w43_,
		_w1333_
	);
	LUT4 #(
		.INIT('h135f)
	) name1300 (
		_w52_,
		_w59_,
		_w201_,
		_w158_,
		_w1334_
	);
	LUT3 #(
		.INIT('h80)
	) name1301 (
		_w1333_,
		_w1334_,
		_w1332_,
		_w1335_
	);
	LUT3 #(
		.INIT('h80)
	) name1302 (
		_w1331_,
		_w1327_,
		_w1335_,
		_w1336_
	);
	LUT4 #(
		.INIT('h135f)
	) name1303 (
		_w78_,
		_w43_,
		_w93_,
		_w44_,
		_w1337_
	);
	LUT2 #(
		.INIT('h4)
	) name1304 (
		_w276_,
		_w1337_,
		_w1338_
	);
	LUT4 #(
		.INIT('h135f)
	) name1305 (
		_w56_,
		_w44_,
		_w184_,
		_w201_,
		_w1339_
	);
	LUT4 #(
		.INIT('h153f)
	) name1306 (
		_w52_,
		_w59_,
		_w419_,
		_w430_,
		_w1340_
	);
	LUT3 #(
		.INIT('h57)
	) name1307 (
		_w93_,
		_w201_,
		_w430_,
		_w1341_
	);
	LUT4 #(
		.INIT('h153f)
	) name1308 (
		_w38_,
		_w56_,
		_w43_,
		_w236_,
		_w1342_
	);
	LUT4 #(
		.INIT('h8000)
	) name1309 (
		_w1341_,
		_w1342_,
		_w1339_,
		_w1340_,
		_w1343_
	);
	LUT2 #(
		.INIT('h8)
	) name1310 (
		_w496_,
		_w806_,
		_w1344_
	);
	LUT4 #(
		.INIT('h135f)
	) name1311 (
		_w41_,
		_w72_,
		_w39_,
		_w65_,
		_w1345_
	);
	LUT4 #(
		.INIT('h135f)
	) name1312 (
		_w85_,
		_w67_,
		_w176_,
		_w419_,
		_w1346_
	);
	LUT4 #(
		.INIT('h153f)
	) name1313 (
		_w85_,
		_w67_,
		_w39_,
		_w43_,
		_w1347_
	);
	LUT4 #(
		.INIT('h8000)
	) name1314 (
		_w969_,
		_w1347_,
		_w1345_,
		_w1346_,
		_w1348_
	);
	LUT4 #(
		.INIT('h8000)
	) name1315 (
		_w1344_,
		_w1338_,
		_w1343_,
		_w1348_,
		_w1349_
	);
	LUT4 #(
		.INIT('h0777)
	) name1316 (
		_w85_,
		_w72_,
		_w65_,
		_w201_,
		_w1350_
	);
	LUT4 #(
		.INIT('h135f)
	) name1317 (
		_w56_,
		_w47_,
		_w158_,
		_w430_,
		_w1351_
	);
	LUT4 #(
		.INIT('h135f)
	) name1318 (
		_w67_,
		_w46_,
		_w201_,
		_w176_,
		_w1352_
	);
	LUT4 #(
		.INIT('h8000)
	) name1319 (
		_w584_,
		_w1350_,
		_w1351_,
		_w1352_,
		_w1353_
	);
	LUT4 #(
		.INIT('h0777)
	) name1320 (
		_w78_,
		_w90_,
		_w47_,
		_w201_,
		_w1354_
	);
	LUT4 #(
		.INIT('h135f)
	) name1321 (
		_w93_,
		_w44_,
		_w176_,
		_w419_,
		_w1355_
	);
	LUT4 #(
		.INIT('h135f)
	) name1322 (
		_w85_,
		_w65_,
		_w166_,
		_w378_,
		_w1356_
	);
	LUT2 #(
		.INIT('h4)
	) name1323 (
		_w473_,
		_w1356_,
		_w1357_
	);
	LUT4 #(
		.INIT('h4000)
	) name1324 (
		_w473_,
		_w1354_,
		_w1355_,
		_w1356_,
		_w1358_
	);
	LUT4 #(
		.INIT('h0777)
	) name1325 (
		_w59_,
		_w72_,
		_w39_,
		_w50_,
		_w1359_
	);
	LUT4 #(
		.INIT('h135f)
	) name1326 (
		_w106_,
		_w55_,
		_w52_,
		_w430_,
		_w1360_
	);
	LUT3 #(
		.INIT('h80)
	) name1327 (
		_w1067_,
		_w1360_,
		_w1359_,
		_w1361_
	);
	LUT4 #(
		.INIT('h0777)
	) name1328 (
		_w55_,
		_w78_,
		_w47_,
		_w184_,
		_w1362_
	);
	LUT2 #(
		.INIT('h4)
	) name1329 (
		_w114_,
		_w1362_,
		_w1363_
	);
	LUT4 #(
		.INIT('h153f)
	) name1330 (
		_w38_,
		_w67_,
		_w184_,
		_w201_,
		_w1364_
	);
	LUT4 #(
		.INIT('h4000)
	) name1331 (
		_w114_,
		_w651_,
		_w1362_,
		_w1364_,
		_w1365_
	);
	LUT4 #(
		.INIT('h8000)
	) name1332 (
		_w1361_,
		_w1365_,
		_w1353_,
		_w1358_,
		_w1366_
	);
	LUT4 #(
		.INIT('h8000)
	) name1333 (
		_w1228_,
		_w1336_,
		_w1349_,
		_w1366_,
		_w1367_
	);
	LUT2 #(
		.INIT('h8)
	) name1334 (
		_w1325_,
		_w1367_,
		_w1368_
	);
	LUT2 #(
		.INIT('h4)
	) name1335 (
		_w468_,
		_w611_,
		_w1369_
	);
	LUT3 #(
		.INIT('h40)
	) name1336 (
		_w468_,
		_w611_,
		_w975_,
		_w1370_
	);
	LUT4 #(
		.INIT('h135f)
	) name1337 (
		_w38_,
		_w85_,
		_w176_,
		_w430_,
		_w1371_
	);
	LUT4 #(
		.INIT('h0777)
	) name1338 (
		_w106_,
		_w67_,
		_w56_,
		_w201_,
		_w1372_
	);
	LUT3 #(
		.INIT('h1f)
	) name1339 (
		_w41_,
		_w93_,
		_w378_,
		_w1373_
	);
	LUT3 #(
		.INIT('h1f)
	) name1340 (
		_w85_,
		_w90_,
		_w201_,
		_w1374_
	);
	LUT4 #(
		.INIT('h8000)
	) name1341 (
		_w1371_,
		_w1372_,
		_w1373_,
		_w1374_,
		_w1375_
	);
	LUT3 #(
		.INIT('h80)
	) name1342 (
		_w1110_,
		_w1370_,
		_w1375_,
		_w1376_
	);
	LUT4 #(
		.INIT('h0777)
	) name1343 (
		_w122_,
		_w59_,
		_w78_,
		_w41_,
		_w1377_
	);
	LUT2 #(
		.INIT('h4)
	) name1344 (
		_w276_,
		_w1377_,
		_w1378_
	);
	LUT4 #(
		.INIT('h8000)
	) name1345 (
		_w66_,
		_w456_,
		_w649_,
		_w1068_,
		_w1379_
	);
	LUT4 #(
		.INIT('h8000)
	) name1346 (
		_w1183_,
		_w1185_,
		_w1378_,
		_w1379_,
		_w1380_
	);
	LUT2 #(
		.INIT('h8)
	) name1347 (
		_w1376_,
		_w1380_,
		_w1381_
	);
	LUT4 #(
		.INIT('h153f)
	) name1348 (
		_w85_,
		_w52_,
		_w43_,
		_w236_,
		_w1382_
	);
	LUT4 #(
		.INIT('h1000)
	) name1349 (
		_w162_,
		_w365_,
		_w1237_,
		_w1382_,
		_w1383_
	);
	LUT4 #(
		.INIT('h135f)
	) name1350 (
		_w47_,
		_w41_,
		_w72_,
		_w259_,
		_w1384_
	);
	LUT4 #(
		.INIT('h153f)
	) name1351 (
		_w90_,
		_w93_,
		_w259_,
		_w176_,
		_w1385_
	);
	LUT4 #(
		.INIT('h135f)
	) name1352 (
		_w122_,
		_w55_,
		_w44_,
		_w166_,
		_w1386_
	);
	LUT4 #(
		.INIT('h4000)
	) name1353 (
		_w407_,
		_w1384_,
		_w1385_,
		_w1386_,
		_w1387_
	);
	LUT4 #(
		.INIT('h135f)
	) name1354 (
		_w85_,
		_w52_,
		_w176_,
		_w419_,
		_w1388_
	);
	LUT3 #(
		.INIT('h80)
	) name1355 (
		_w919_,
		_w1078_,
		_w1388_,
		_w1389_
	);
	LUT4 #(
		.INIT('h0777)
	) name1356 (
		_w78_,
		_w56_,
		_w39_,
		_w93_,
		_w1390_
	);
	LUT3 #(
		.INIT('h80)
	) name1357 (
		_w643_,
		_w894_,
		_w1390_,
		_w1391_
	);
	LUT4 #(
		.INIT('h8000)
	) name1358 (
		_w1389_,
		_w1391_,
		_w1383_,
		_w1387_,
		_w1392_
	);
	LUT4 #(
		.INIT('h0777)
	) name1359 (
		_w106_,
		_w85_,
		_w67_,
		_w39_,
		_w1393_
	);
	LUT2 #(
		.INIT('h4)
	) name1360 (
		_w215_,
		_w1393_,
		_w1394_
	);
	LUT3 #(
		.INIT('h57)
	) name1361 (
		_w110_,
		_w158_,
		_w176_,
		_w1395_
	);
	LUT3 #(
		.INIT('h80)
	) name1362 (
		_w495_,
		_w941_,
		_w1395_,
		_w1396_
	);
	LUT4 #(
		.INIT('h8000)
	) name1363 (
		_w1175_,
		_w1178_,
		_w1394_,
		_w1396_,
		_w1397_
	);
	LUT4 #(
		.INIT('h8000)
	) name1364 (
		_w1228_,
		_w1366_,
		_w1392_,
		_w1397_,
		_w1398_
	);
	LUT2 #(
		.INIT('h8)
	) name1365 (
		_w1381_,
		_w1398_,
		_w1399_
	);
	LUT4 #(
		.INIT('h0777)
	) name1366 (
		_w1325_,
		_w1367_,
		_w1381_,
		_w1398_,
		_w1400_
	);
	LUT4 #(
		.INIT('h153f)
	) name1367 (
		_w78_,
		_w41_,
		_w39_,
		_w46_,
		_w1401_
	);
	LUT4 #(
		.INIT('h153f)
	) name1368 (
		_w55_,
		_w41_,
		_w166_,
		_w259_,
		_w1402_
	);
	LUT4 #(
		.INIT('h135f)
	) name1369 (
		_w122_,
		_w106_,
		_w67_,
		_w65_,
		_w1403_
	);
	LUT4 #(
		.INIT('h8000)
	) name1370 (
		_w829_,
		_w1401_,
		_w1402_,
		_w1403_,
		_w1404_
	);
	LUT3 #(
		.INIT('h57)
	) name1371 (
		_w122_,
		_w55_,
		_w90_,
		_w1405_
	);
	LUT4 #(
		.INIT('h4000)
	) name1372 (
		_w64_,
		_w769_,
		_w1143_,
		_w1405_,
		_w1406_
	);
	LUT3 #(
		.INIT('h80)
	) name1373 (
		_w1117_,
		_w1404_,
		_w1406_,
		_w1407_
	);
	LUT4 #(
		.INIT('h153f)
	) name1374 (
		_w55_,
		_w90_,
		_w236_,
		_w158_,
		_w1408_
	);
	LUT4 #(
		.INIT('h1000)
	) name1375 (
		_w186_,
		_w435_,
		_w971_,
		_w1408_,
		_w1409_
	);
	LUT4 #(
		.INIT('h153f)
	) name1376 (
		_w59_,
		_w56_,
		_w201_,
		_w378_,
		_w1410_
	);
	LUT4 #(
		.INIT('h153f)
	) name1377 (
		_w90_,
		_w47_,
		_w236_,
		_w430_,
		_w1411_
	);
	LUT4 #(
		.INIT('h8000)
	) name1378 (
		_w68_,
		_w777_,
		_w1410_,
		_w1411_,
		_w1412_
	);
	LUT2 #(
		.INIT('h8)
	) name1379 (
		_w1409_,
		_w1412_,
		_w1413_
	);
	LUT4 #(
		.INIT('h153f)
	) name1380 (
		_w90_,
		_w50_,
		_w236_,
		_w166_,
		_w1414_
	);
	LUT4 #(
		.INIT('h135f)
	) name1381 (
		_w65_,
		_w44_,
		_w176_,
		_w419_,
		_w1415_
	);
	LUT4 #(
		.INIT('h153f)
	) name1382 (
		_w55_,
		_w78_,
		_w47_,
		_w430_,
		_w1416_
	);
	LUT3 #(
		.INIT('h80)
	) name1383 (
		_w1415_,
		_w1416_,
		_w1414_,
		_w1417_
	);
	LUT4 #(
		.INIT('h153f)
	) name1384 (
		_w52_,
		_w110_,
		_w72_,
		_w184_,
		_w1418_
	);
	LUT4 #(
		.INIT('h8000)
	) name1385 (
		_w198_,
		_w957_,
		_w1297_,
		_w1418_,
		_w1419_
	);
	LUT4 #(
		.INIT('h0777)
	) name1386 (
		_w122_,
		_w110_,
		_w41_,
		_w72_,
		_w1420_
	);
	LUT4 #(
		.INIT('h135f)
	) name1387 (
		_w56_,
		_w44_,
		_w259_,
		_w176_,
		_w1421_
	);
	LUT3 #(
		.INIT('h80)
	) name1388 (
		_w924_,
		_w1420_,
		_w1421_,
		_w1422_
	);
	LUT4 #(
		.INIT('h153f)
	) name1389 (
		_w38_,
		_w47_,
		_w72_,
		_w259_,
		_w1423_
	);
	LUT3 #(
		.INIT('h40)
	) name1390 (
		_w151_,
		_w710_,
		_w1423_,
		_w1424_
	);
	LUT4 #(
		.INIT('h8000)
	) name1391 (
		_w1422_,
		_w1424_,
		_w1417_,
		_w1419_,
		_w1425_
	);
	LUT3 #(
		.INIT('h80)
	) name1392 (
		_w1407_,
		_w1413_,
		_w1425_,
		_w1426_
	);
	LUT4 #(
		.INIT('h0777)
	) name1393 (
		_w67_,
		_w72_,
		_w65_,
		_w236_,
		_w1427_
	);
	LUT2 #(
		.INIT('h4)
	) name1394 (
		_w45_,
		_w1427_,
		_w1428_
	);
	LUT4 #(
		.INIT('h135f)
	) name1395 (
		_w55_,
		_w52_,
		_w39_,
		_w43_,
		_w1429_
	);
	LUT4 #(
		.INIT('h135f)
	) name1396 (
		_w55_,
		_w85_,
		_w184_,
		_w378_,
		_w1430_
	);
	LUT3 #(
		.INIT('h1f)
	) name1397 (
		_w55_,
		_w67_,
		_w419_,
		_w1431_
	);
	LUT4 #(
		.INIT('h4000)
	) name1398 (
		_w253_,
		_w1429_,
		_w1430_,
		_w1431_,
		_w1432_
	);
	LUT4 #(
		.INIT('h0777)
	) name1399 (
		_w106_,
		_w52_,
		_w67_,
		_w43_,
		_w1433_
	);
	LUT3 #(
		.INIT('h57)
	) name1400 (
		_w55_,
		_w43_,
		_w176_,
		_w1434_
	);
	LUT4 #(
		.INIT('h135f)
	) name1401 (
		_w85_,
		_w110_,
		_w236_,
		_w259_,
		_w1435_
	);
	LUT3 #(
		.INIT('h80)
	) name1402 (
		_w1434_,
		_w1435_,
		_w1433_,
		_w1436_
	);
	LUT4 #(
		.INIT('h135f)
	) name1403 (
		_w44_,
		_w46_,
		_w201_,
		_w419_,
		_w1437_
	);
	LUT4 #(
		.INIT('h0777)
	) name1404 (
		_w59_,
		_w78_,
		_w65_,
		_w166_,
		_w1438_
	);
	LUT4 #(
		.INIT('h153f)
	) name1405 (
		_w38_,
		_w41_,
		_w201_,
		_w430_,
		_w1439_
	);
	LUT3 #(
		.INIT('h80)
	) name1406 (
		_w1438_,
		_w1439_,
		_w1437_,
		_w1440_
	);
	LUT4 #(
		.INIT('h8000)
	) name1407 (
		_w1436_,
		_w1428_,
		_w1440_,
		_w1432_,
		_w1441_
	);
	LUT4 #(
		.INIT('h0777)
	) name1408 (
		_w38_,
		_w122_,
		_w67_,
		_w78_,
		_w1442_
	);
	LUT2 #(
		.INIT('h4)
	) name1409 (
		_w160_,
		_w1442_,
		_w1443_
	);
	LUT4 #(
		.INIT('h135f)
	) name1410 (
		_w85_,
		_w93_,
		_w184_,
		_w166_,
		_w1444_
	);
	LUT4 #(
		.INIT('h0777)
	) name1411 (
		_w106_,
		_w90_,
		_w46_,
		_w259_,
		_w1445_
	);
	LUT3 #(
		.INIT('h40)
	) name1412 (
		_w452_,
		_w1444_,
		_w1445_,
		_w1446_
	);
	LUT3 #(
		.INIT('h57)
	) name1413 (
		_w38_,
		_w106_,
		_w166_,
		_w1447_
	);
	LUT4 #(
		.INIT('h135f)
	) name1414 (
		_w78_,
		_w39_,
		_w50_,
		_w65_,
		_w1448_
	);
	LUT3 #(
		.INIT('h80)
	) name1415 (
		_w1362_,
		_w1448_,
		_w1447_,
		_w1449_
	);
	LUT4 #(
		.INIT('h135f)
	) name1416 (
		_w59_,
		_w93_,
		_w184_,
		_w176_,
		_w1450_
	);
	LUT4 #(
		.INIT('h153f)
	) name1417 (
		_w55_,
		_w50_,
		_w184_,
		_w236_,
		_w1451_
	);
	LUT4 #(
		.INIT('h1000)
	) name1418 (
		_w104_,
		_w339_,
		_w1450_,
		_w1451_,
		_w1452_
	);
	LUT4 #(
		.INIT('h8000)
	) name1419 (
		_w1443_,
		_w1446_,
		_w1449_,
		_w1452_,
		_w1453_
	);
	LUT2 #(
		.INIT('h8)
	) name1420 (
		_w1441_,
		_w1453_,
		_w1454_
	);
	LUT4 #(
		.INIT('h153f)
	) name1421 (
		_w38_,
		_w106_,
		_w59_,
		_w236_,
		_w1455_
	);
	LUT4 #(
		.INIT('h153f)
	) name1422 (
		_w122_,
		_w52_,
		_w39_,
		_w46_,
		_w1456_
	);
	LUT3 #(
		.INIT('h80)
	) name1423 (
		_w1113_,
		_w1456_,
		_w1455_,
		_w1457_
	);
	LUT4 #(
		.INIT('h113f)
	) name1424 (
		_w59_,
		_w50_,
		_w158_,
		_w176_,
		_w1458_
	);
	LUT4 #(
		.INIT('h153f)
	) name1425 (
		_w41_,
		_w72_,
		_w93_,
		_w184_,
		_w1459_
	);
	LUT4 #(
		.INIT('h135f)
	) name1426 (
		_w106_,
		_w110_,
		_w50_,
		_w236_,
		_w1460_
	);
	LUT4 #(
		.INIT('h4000)
	) name1427 (
		_w152_,
		_w783_,
		_w1459_,
		_w1460_,
		_w1461_
	);
	LUT3 #(
		.INIT('h80)
	) name1428 (
		_w1458_,
		_w1457_,
		_w1461_,
		_w1462_
	);
	LUT4 #(
		.INIT('h153f)
	) name1429 (
		_w110_,
		_w90_,
		_w184_,
		_w201_,
		_w1463_
	);
	LUT4 #(
		.INIT('h135f)
	) name1430 (
		_w85_,
		_w93_,
		_w158_,
		_w419_,
		_w1464_
	);
	LUT2 #(
		.INIT('h8)
	) name1431 (
		_w1463_,
		_w1464_,
		_w1465_
	);
	LUT4 #(
		.INIT('h135f)
	) name1432 (
		_w38_,
		_w59_,
		_w78_,
		_w259_,
		_w1466_
	);
	LUT3 #(
		.INIT('h80)
	) name1433 (
		_w408_,
		_w610_,
		_w1466_,
		_w1467_
	);
	LUT2 #(
		.INIT('h8)
	) name1434 (
		_w1465_,
		_w1467_,
		_w1468_
	);
	LUT4 #(
		.INIT('h135f)
	) name1435 (
		_w38_,
		_w56_,
		_w201_,
		_w176_,
		_w1469_
	);
	LUT4 #(
		.INIT('h135f)
	) name1436 (
		_w85_,
		_w65_,
		_w419_,
		_w430_,
		_w1470_
	);
	LUT4 #(
		.INIT('h2000)
	) name1437 (
		_w225_,
		_w354_,
		_w1470_,
		_w1469_,
		_w1471_
	);
	LUT4 #(
		.INIT('h153f)
	) name1438 (
		_w56_,
		_w41_,
		_w378_,
		_w430_,
		_w1472_
	);
	LUT4 #(
		.INIT('h0777)
	) name1439 (
		_w38_,
		_w43_,
		_w65_,
		_w419_,
		_w1473_
	);
	LUT4 #(
		.INIT('h135f)
	) name1440 (
		_w85_,
		_w56_,
		_w43_,
		_w166_,
		_w1474_
	);
	LUT4 #(
		.INIT('h135f)
	) name1441 (
		_w55_,
		_w93_,
		_w201_,
		_w378_,
		_w1475_
	);
	LUT4 #(
		.INIT('h8000)
	) name1442 (
		_w1472_,
		_w1473_,
		_w1474_,
		_w1475_,
		_w1476_
	);
	LUT4 #(
		.INIT('h8000)
	) name1443 (
		_w1155_,
		_w1369_,
		_w1476_,
		_w1471_,
		_w1477_
	);
	LUT3 #(
		.INIT('h80)
	) name1444 (
		_w1468_,
		_w1462_,
		_w1477_,
		_w1478_
	);
	LUT3 #(
		.INIT('h80)
	) name1445 (
		_w1454_,
		_w1426_,
		_w1478_,
		_w1479_
	);
	LUT4 #(
		.INIT('h135f)
	) name1446 (
		_w78_,
		_w41_,
		_w93_,
		_w166_,
		_w1480_
	);
	LUT4 #(
		.INIT('h135f)
	) name1447 (
		_w106_,
		_w93_,
		_w65_,
		_w166_,
		_w1481_
	);
	LUT3 #(
		.INIT('h80)
	) name1448 (
		_w1334_,
		_w1481_,
		_w1480_,
		_w1482_
	);
	LUT4 #(
		.INIT('h153f)
	) name1449 (
		_w47_,
		_w43_,
		_w93_,
		_w430_,
		_w1483_
	);
	LUT4 #(
		.INIT('h153f)
	) name1450 (
		_w106_,
		_w67_,
		_w78_,
		_w44_,
		_w1484_
	);
	LUT2 #(
		.INIT('h8)
	) name1451 (
		_w1483_,
		_w1484_,
		_w1485_
	);
	LUT4 #(
		.INIT('h153f)
	) name1452 (
		_w38_,
		_w110_,
		_w184_,
		_w158_,
		_w1486_
	);
	LUT4 #(
		.INIT('h4000)
	) name1453 (
		_w410_,
		_w1384_,
		_w1385_,
		_w1486_,
		_w1487_
	);
	LUT3 #(
		.INIT('h80)
	) name1454 (
		_w1485_,
		_w1482_,
		_w1487_,
		_w1488_
	);
	LUT3 #(
		.INIT('h40)
	) name1455 (
		_w308_,
		_w428_,
		_w1328_,
		_w1489_
	);
	LUT4 #(
		.INIT('h153f)
	) name1456 (
		_w52_,
		_w65_,
		_w166_,
		_w158_,
		_w1490_
	);
	LUT4 #(
		.INIT('h1000)
	) name1457 (
		_w114_,
		_w160_,
		_w1362_,
		_w1490_,
		_w1491_
	);
	LUT4 #(
		.INIT('h153f)
	) name1458 (
		_w90_,
		_w65_,
		_w236_,
		_w259_,
		_w1492_
	);
	LUT4 #(
		.INIT('h135f)
	) name1459 (
		_w55_,
		_w110_,
		_w72_,
		_w201_,
		_w1493_
	);
	LUT4 #(
		.INIT('h153f)
	) name1460 (
		_w55_,
		_w52_,
		_w72_,
		_w378_,
		_w1494_
	);
	LUT3 #(
		.INIT('h80)
	) name1461 (
		_w1493_,
		_w1494_,
		_w1492_,
		_w1495_
	);
	LUT4 #(
		.INIT('h153f)
	) name1462 (
		_w47_,
		_w39_,
		_w93_,
		_w166_,
		_w1496_
	);
	LUT4 #(
		.INIT('h153f)
	) name1463 (
		_w110_,
		_w78_,
		_w65_,
		_w158_,
		_w1497_
	);
	LUT4 #(
		.INIT('h8000)
	) name1464 (
		_w265_,
		_w1472_,
		_w1496_,
		_w1497_,
		_w1498_
	);
	LUT4 #(
		.INIT('h8000)
	) name1465 (
		_w1495_,
		_w1498_,
		_w1489_,
		_w1491_,
		_w1499_
	);
	LUT2 #(
		.INIT('h4)
	) name1466 (
		_w303_,
		_w370_,
		_w1500_
	);
	LUT3 #(
		.INIT('h80)
	) name1467 (
		_w1488_,
		_w1499_,
		_w1500_,
		_w1501_
	);
	LUT4 #(
		.INIT('h135f)
	) name1468 (
		_w110_,
		_w47_,
		_w39_,
		_w378_,
		_w1502_
	);
	LUT2 #(
		.INIT('h8)
	) name1469 (
		_w902_,
		_w1502_,
		_w1503_
	);
	LUT4 #(
		.INIT('h135f)
	) name1470 (
		_w122_,
		_w55_,
		_w65_,
		_w236_,
		_w1504_
	);
	LUT4 #(
		.INIT('h135f)
	) name1471 (
		_w122_,
		_w85_,
		_w56_,
		_w419_,
		_w1505_
	);
	LUT4 #(
		.INIT('h135f)
	) name1472 (
		_w38_,
		_w59_,
		_w43_,
		_w430_,
		_w1506_
	);
	LUT4 #(
		.INIT('h8000)
	) name1473 (
		_w1359_,
		_w1504_,
		_w1505_,
		_w1506_,
		_w1507_
	);
	LUT2 #(
		.INIT('h8)
	) name1474 (
		_w1503_,
		_w1507_,
		_w1508_
	);
	LUT3 #(
		.INIT('h80)
	) name1475 (
		_w579_,
		_w589_,
		_w894_,
		_w1509_
	);
	LUT4 #(
		.INIT('h153f)
	) name1476 (
		_w41_,
		_w44_,
		_w184_,
		_w419_,
		_w1510_
	);
	LUT4 #(
		.INIT('h153f)
	) name1477 (
		_w50_,
		_w44_,
		_w236_,
		_w378_,
		_w1511_
	);
	LUT4 #(
		.INIT('h4000)
	) name1478 (
		_w53_,
		_w262_,
		_w1510_,
		_w1511_,
		_w1512_
	);
	LUT4 #(
		.INIT('h135f)
	) name1479 (
		_w55_,
		_w93_,
		_w259_,
		_w378_,
		_w1513_
	);
	LUT4 #(
		.INIT('h135f)
	) name1480 (
		_w38_,
		_w59_,
		_w39_,
		_w378_,
		_w1514_
	);
	LUT4 #(
		.INIT('h153f)
	) name1481 (
		_w85_,
		_w59_,
		_w236_,
		_w176_,
		_w1515_
	);
	LUT3 #(
		.INIT('h80)
	) name1482 (
		_w1514_,
		_w1513_,
		_w1515_,
		_w1516_
	);
	LUT4 #(
		.INIT('h8000)
	) name1483 (
		_w1171_,
		_w1516_,
		_w1509_,
		_w1512_,
		_w1517_
	);
	LUT4 #(
		.INIT('h153f)
	) name1484 (
		_w65_,
		_w44_,
		_w201_,
		_w430_,
		_w1518_
	);
	LUT4 #(
		.INIT('h0777)
	) name1485 (
		_w78_,
		_w56_,
		_w43_,
		_w65_,
		_w1519_
	);
	LUT4 #(
		.INIT('h8000)
	) name1486 (
		_w777_,
		_w868_,
		_w1518_,
		_w1519_,
		_w1520_
	);
	LUT4 #(
		.INIT('h135f)
	) name1487 (
		_w122_,
		_w55_,
		_w90_,
		_w39_,
		_w1521_
	);
	LUT2 #(
		.INIT('h4)
	) name1488 (
		_w380_,
		_w1521_,
		_w1522_
	);
	LUT4 #(
		.INIT('h0777)
	) name1489 (
		_w78_,
		_w90_,
		_w41_,
		_w72_,
		_w1523_
	);
	LUT4 #(
		.INIT('h153f)
	) name1490 (
		_w59_,
		_w67_,
		_w184_,
		_w259_,
		_w1524_
	);
	LUT4 #(
		.INIT('h135f)
	) name1491 (
		_w38_,
		_w41_,
		_w184_,
		_w158_,
		_w1525_
	);
	LUT4 #(
		.INIT('h135f)
	) name1492 (
		_w38_,
		_w47_,
		_w236_,
		_w176_,
		_w1526_
	);
	LUT4 #(
		.INIT('h8000)
	) name1493 (
		_w1523_,
		_w1524_,
		_w1525_,
		_w1526_,
		_w1527_
	);
	LUT3 #(
		.INIT('h80)
	) name1494 (
		_w1522_,
		_w1520_,
		_w1527_,
		_w1528_
	);
	LUT4 #(
		.INIT('h135f)
	) name1495 (
		_w122_,
		_w106_,
		_w55_,
		_w50_,
		_w1529_
	);
	LUT4 #(
		.INIT('h0777)
	) name1496 (
		_w72_,
		_w65_,
		_w46_,
		_w158_,
		_w1530_
	);
	LUT3 #(
		.INIT('h80)
	) name1497 (
		_w1173_,
		_w1530_,
		_w1529_,
		_w1531_
	);
	LUT4 #(
		.INIT('h0777)
	) name1498 (
		_w59_,
		_w78_,
		_w93_,
		_w236_,
		_w1532_
	);
	LUT4 #(
		.INIT('h135f)
	) name1499 (
		_w56_,
		_w46_,
		_w158_,
		_w378_,
		_w1533_
	);
	LUT4 #(
		.INIT('h0777)
	) name1500 (
		_w122_,
		_w85_,
		_w56_,
		_w39_,
		_w1534_
	);
	LUT4 #(
		.INIT('h8000)
	) name1501 (
		_w886_,
		_w1534_,
		_w1532_,
		_w1533_,
		_w1535_
	);
	LUT2 #(
		.INIT('h8)
	) name1502 (
		_w1531_,
		_w1535_,
		_w1536_
	);
	LUT4 #(
		.INIT('h153f)
	) name1503 (
		_w85_,
		_w59_,
		_w201_,
		_w430_,
		_w1537_
	);
	LUT4 #(
		.INIT('h135f)
	) name1504 (
		_w56_,
		_w93_,
		_w201_,
		_w158_,
		_w1538_
	);
	LUT3 #(
		.INIT('h80)
	) name1505 (
		_w287_,
		_w1537_,
		_w1538_,
		_w1539_
	);
	LUT4 #(
		.INIT('h153f)
	) name1506 (
		_w110_,
		_w47_,
		_w43_,
		_w166_,
		_w1540_
	);
	LUT4 #(
		.INIT('h135f)
	) name1507 (
		_w90_,
		_w50_,
		_w184_,
		_w259_,
		_w1541_
	);
	LUT4 #(
		.INIT('h153f)
	) name1508 (
		_w85_,
		_w59_,
		_w43_,
		_w166_,
		_w1542_
	);
	LUT4 #(
		.INIT('h4000)
	) name1509 (
		_w360_,
		_w1540_,
		_w1541_,
		_w1542_,
		_w1543_
	);
	LUT4 #(
		.INIT('h8000)
	) name1510 (
		_w1531_,
		_w1535_,
		_w1539_,
		_w1543_,
		_w1544_
	);
	LUT4 #(
		.INIT('h8000)
	) name1511 (
		_w1508_,
		_w1517_,
		_w1528_,
		_w1544_,
		_w1545_
	);
	LUT2 #(
		.INIT('h8)
	) name1512 (
		_w1501_,
		_w1545_,
		_w1546_
	);
	LUT2 #(
		.INIT('h1)
	) name1513 (
		_w1479_,
		_w1546_,
		_w1547_
	);
	LUT2 #(
		.INIT('h4)
	) name1514 (
		_w267_,
		_w979_,
		_w1548_
	);
	LUT3 #(
		.INIT('h57)
	) name1515 (
		_w47_,
		_w39_,
		_w176_,
		_w1549_
	);
	LUT4 #(
		.INIT('h0777)
	) name1516 (
		_w55_,
		_w43_,
		_w44_,
		_w378_,
		_w1550_
	);
	LUT4 #(
		.INIT('h153f)
	) name1517 (
		_w47_,
		_w72_,
		_w44_,
		_w158_,
		_w1551_
	);
	LUT3 #(
		.INIT('h80)
	) name1518 (
		_w1550_,
		_w1551_,
		_w1549_,
		_w1552_
	);
	LUT3 #(
		.INIT('h80)
	) name1519 (
		_w1516_,
		_w1548_,
		_w1552_,
		_w1553_
	);
	LUT4 #(
		.INIT('h153f)
	) name1520 (
		_w90_,
		_w56_,
		_w184_,
		_w201_,
		_w1554_
	);
	LUT2 #(
		.INIT('h4)
	) name1521 (
		_w270_,
		_w1554_,
		_w1555_
	);
	LUT4 #(
		.INIT('h135f)
	) name1522 (
		_w72_,
		_w39_,
		_w50_,
		_w93_,
		_w1556_
	);
	LUT4 #(
		.INIT('h135f)
	) name1523 (
		_w67_,
		_w44_,
		_w236_,
		_w176_,
		_w1557_
	);
	LUT3 #(
		.INIT('h80)
	) name1524 (
		_w1192_,
		_w1557_,
		_w1556_,
		_w1558_
	);
	LUT2 #(
		.INIT('h8)
	) name1525 (
		_w1555_,
		_w1558_,
		_w1559_
	);
	LUT4 #(
		.INIT('h153f)
	) name1526 (
		_w52_,
		_w110_,
		_w72_,
		_w166_,
		_w1560_
	);
	LUT4 #(
		.INIT('h0777)
	) name1527 (
		_w78_,
		_w65_,
		_w46_,
		_w419_,
		_w1561_
	);
	LUT4 #(
		.INIT('h153f)
	) name1528 (
		_w67_,
		_w93_,
		_w201_,
		_w166_,
		_w1562_
	);
	LUT4 #(
		.INIT('h8000)
	) name1529 (
		_w514_,
		_w1560_,
		_w1561_,
		_w1562_,
		_w1563_
	);
	LUT3 #(
		.INIT('h57)
	) name1530 (
		_w93_,
		_w184_,
		_w236_,
		_w1564_
	);
	LUT2 #(
		.INIT('h4)
	) name1531 (
		_w335_,
		_w1564_,
		_w1565_
	);
	LUT4 #(
		.INIT('h135f)
	) name1532 (
		_w106_,
		_w67_,
		_w90_,
		_w43_,
		_w1566_
	);
	LUT3 #(
		.INIT('h80)
	) name1533 (
		_w143_,
		_w163_,
		_w1566_,
		_w1567_
	);
	LUT3 #(
		.INIT('h80)
	) name1534 (
		_w1565_,
		_w1563_,
		_w1567_,
		_w1568_
	);
	LUT3 #(
		.INIT('h80)
	) name1535 (
		_w1559_,
		_w1553_,
		_w1568_,
		_w1569_
	);
	LUT4 #(
		.INIT('h0777)
	) name1536 (
		_w106_,
		_w110_,
		_w46_,
		_w158_,
		_w1570_
	);
	LUT2 #(
		.INIT('h8)
	) name1537 (
		_w650_,
		_w1570_,
		_w1571_
	);
	LUT3 #(
		.INIT('h57)
	) name1538 (
		_w39_,
		_w65_,
		_w46_,
		_w1572_
	);
	LUT4 #(
		.INIT('h1000)
	) name1539 (
		_w45_,
		_w338_,
		_w1427_,
		_w1572_,
		_w1573_
	);
	LUT2 #(
		.INIT('h8)
	) name1540 (
		_w1571_,
		_w1573_,
		_w1574_
	);
	LUT3 #(
		.INIT('h37)
	) name1541 (
		_w106_,
		_w46_,
		_w201_,
		_w1575_
	);
	LUT4 #(
		.INIT('h0777)
	) name1542 (
		_w122_,
		_w52_,
		_w44_,
		_w201_,
		_w1576_
	);
	LUT4 #(
		.INIT('h8000)
	) name1543 (
		_w1235_,
		_w1483_,
		_w1575_,
		_w1576_,
		_w1577_
	);
	LUT4 #(
		.INIT('h8000)
	) name1544 (
		_w112_,
		_w408_,
		_w990_,
		_w1124_,
		_w1578_
	);
	LUT3 #(
		.INIT('h40)
	) name1545 (
		_w363_,
		_w790_,
		_w1360_,
		_w1579_
	);
	LUT4 #(
		.INIT('h153f)
	) name1546 (
		_w41_,
		_w50_,
		_w184_,
		_w166_,
		_w1580_
	);
	LUT4 #(
		.INIT('h153f)
	) name1547 (
		_w38_,
		_w52_,
		_w72_,
		_w176_,
		_w1581_
	);
	LUT3 #(
		.INIT('h40)
	) name1548 (
		_w346_,
		_w1580_,
		_w1581_,
		_w1582_
	);
	LUT4 #(
		.INIT('h8000)
	) name1549 (
		_w1579_,
		_w1582_,
		_w1577_,
		_w1578_,
		_w1583_
	);
	LUT3 #(
		.INIT('h80)
	) name1550 (
		_w1462_,
		_w1574_,
		_w1583_,
		_w1584_
	);
	LUT4 #(
		.INIT('h135f)
	) name1551 (
		_w122_,
		_w55_,
		_w110_,
		_w78_,
		_w1585_
	);
	LUT4 #(
		.INIT('h0777)
	) name1552 (
		_w72_,
		_w65_,
		_w44_,
		_w236_,
		_w1586_
	);
	LUT4 #(
		.INIT('h0777)
	) name1553 (
		_w90_,
		_w39_,
		_w50_,
		_w378_,
		_w1587_
	);
	LUT4 #(
		.INIT('h8000)
	) name1554 (
		_w1506_,
		_w1585_,
		_w1586_,
		_w1587_,
		_w1588_
	);
	LUT4 #(
		.INIT('h0777)
	) name1555 (
		_w122_,
		_w47_,
		_w44_,
		_w430_,
		_w1589_
	);
	LUT2 #(
		.INIT('h4)
	) name1556 (
		_w362_,
		_w1589_,
		_w1590_
	);
	LUT2 #(
		.INIT('h4)
	) name1557 (
		_w409_,
		_w857_,
		_w1591_
	);
	LUT4 #(
		.INIT('h135f)
	) name1558 (
		_w38_,
		_w55_,
		_w78_,
		_w39_,
		_w1592_
	);
	LUT4 #(
		.INIT('h4000)
	) name1559 (
		_w409_,
		_w890_,
		_w857_,
		_w1592_,
		_w1593_
	);
	LUT3 #(
		.INIT('h80)
	) name1560 (
		_w1590_,
		_w1588_,
		_w1593_,
		_w1594_
	);
	LUT4 #(
		.INIT('h0777)
	) name1561 (
		_w106_,
		_w65_,
		_w46_,
		_w166_,
		_w1595_
	);
	LUT3 #(
		.INIT('h57)
	) name1562 (
		_w110_,
		_w378_,
		_w430_,
		_w1596_
	);
	LUT2 #(
		.INIT('h8)
	) name1563 (
		_w1595_,
		_w1596_,
		_w1597_
	);
	LUT4 #(
		.INIT('h153f)
	) name1564 (
		_w52_,
		_w78_,
		_w44_,
		_w158_,
		_w1598_
	);
	LUT4 #(
		.INIT('h8000)
	) name1565 (
		_w963_,
		_w1247_,
		_w1275_,
		_w1598_,
		_w1599_
	);
	LUT2 #(
		.INIT('h8)
	) name1566 (
		_w1597_,
		_w1599_,
		_w1600_
	);
	LUT2 #(
		.INIT('h4)
	) name1567 (
		_w128_,
		_w54_,
		_w1601_
	);
	LUT4 #(
		.INIT('h135f)
	) name1568 (
		_w85_,
		_w56_,
		_w39_,
		_w259_,
		_w1602_
	);
	LUT4 #(
		.INIT('h0777)
	) name1569 (
		_w78_,
		_w47_,
		_w65_,
		_w430_,
		_w1603_
	);
	LUT3 #(
		.INIT('h80)
	) name1570 (
		_w662_,
		_w1603_,
		_w1602_,
		_w1604_
	);
	LUT4 #(
		.INIT('h8000)
	) name1571 (
		_w1073_,
		_w1076_,
		_w1601_,
		_w1604_,
		_w1605_
	);
	LUT3 #(
		.INIT('h80)
	) name1572 (
		_w1600_,
		_w1594_,
		_w1605_,
		_w1606_
	);
	LUT3 #(
		.INIT('h80)
	) name1573 (
		_w1584_,
		_w1569_,
		_w1606_,
		_w1607_
	);
	LUT3 #(
		.INIT('h80)
	) name1574 (
		_w491_,
		_w660_,
		_w643_,
		_w1608_
	);
	LUT2 #(
		.INIT('h4)
	) name1575 (
		_w369_,
		_w1165_,
		_w1609_
	);
	LUT4 #(
		.INIT('h153f)
	) name1576 (
		_w67_,
		_w41_,
		_w72_,
		_w201_,
		_w1610_
	);
	LUT4 #(
		.INIT('h1000)
	) name1577 (
		_w186_,
		_w477_,
		_w971_,
		_w1610_,
		_w1611_
	);
	LUT3 #(
		.INIT('h80)
	) name1578 (
		_w1609_,
		_w1608_,
		_w1611_,
		_w1612_
	);
	LUT4 #(
		.INIT('h8000)
	) name1579 (
		_w803_,
		_w842_,
		_w937_,
		_w1438_,
		_w1613_
	);
	LUT4 #(
		.INIT('h135f)
	) name1580 (
		_w55_,
		_w47_,
		_w158_,
		_w419_,
		_w1614_
	);
	LUT3 #(
		.INIT('h1f)
	) name1581 (
		_w52_,
		_w59_,
		_w419_,
		_w1615_
	);
	LUT4 #(
		.INIT('h8000)
	) name1582 (
		_w143_,
		_w760_,
		_w1614_,
		_w1615_,
		_w1616_
	);
	LUT4 #(
		.INIT('h153f)
	) name1583 (
		_w78_,
		_w50_,
		_w43_,
		_w46_,
		_w1617_
	);
	LUT4 #(
		.INIT('h4000)
	) name1584 (
		_w285_,
		_w1483_,
		_w1484_,
		_w1617_,
		_w1618_
	);
	LUT3 #(
		.INIT('h80)
	) name1585 (
		_w1613_,
		_w1616_,
		_w1618_,
		_w1619_
	);
	LUT2 #(
		.INIT('h8)
	) name1586 (
		_w1612_,
		_w1619_,
		_w1620_
	);
	LUT4 #(
		.INIT('h153f)
	) name1587 (
		_w38_,
		_w65_,
		_w184_,
		_w158_,
		_w1621_
	);
	LUT3 #(
		.INIT('h1f)
	) name1588 (
		_w59_,
		_w50_,
		_w259_,
		_w1622_
	);
	LUT2 #(
		.INIT('h8)
	) name1589 (
		_w1621_,
		_w1622_,
		_w1623_
	);
	LUT4 #(
		.INIT('h153f)
	) name1590 (
		_w38_,
		_w110_,
		_w236_,
		_w419_,
		_w1624_
	);
	LUT4 #(
		.INIT('h153f)
	) name1591 (
		_w38_,
		_w67_,
		_w236_,
		_w176_,
		_w1625_
	);
	LUT3 #(
		.INIT('h80)
	) name1592 (
		_w964_,
		_w1625_,
		_w1624_,
		_w1626_
	);
	LUT2 #(
		.INIT('h8)
	) name1593 (
		_w1623_,
		_w1626_,
		_w1627_
	);
	LUT4 #(
		.INIT('h0777)
	) name1594 (
		_w55_,
		_w39_,
		_w93_,
		_w378_,
		_w1628_
	);
	LUT4 #(
		.INIT('h135f)
	) name1595 (
		_w122_,
		_w59_,
		_w67_,
		_w158_,
		_w1629_
	);
	LUT4 #(
		.INIT('h8000)
	) name1596 (
		_w1026_,
		_w1164_,
		_w1628_,
		_w1629_,
		_w1630_
	);
	LUT4 #(
		.INIT('h153f)
	) name1597 (
		_w85_,
		_w78_,
		_w56_,
		_w430_,
		_w1631_
	);
	LUT4 #(
		.INIT('h135f)
	) name1598 (
		_w43_,
		_w65_,
		_w46_,
		_w158_,
		_w1632_
	);
	LUT4 #(
		.INIT('h4000)
	) name1599 (
		_w57_,
		_w630_,
		_w1631_,
		_w1632_,
		_w1633_
	);
	LUT4 #(
		.INIT('h153f)
	) name1600 (
		_w65_,
		_w46_,
		_w166_,
		_w259_,
		_w1634_
	);
	LUT4 #(
		.INIT('h153f)
	) name1601 (
		_w52_,
		_w47_,
		_w39_,
		_w259_,
		_w1635_
	);
	LUT4 #(
		.INIT('h135f)
	) name1602 (
		_w38_,
		_w90_,
		_w201_,
		_w236_,
		_w1636_
	);
	LUT3 #(
		.INIT('h80)
	) name1603 (
		_w1635_,
		_w1634_,
		_w1636_,
		_w1637_
	);
	LUT3 #(
		.INIT('h37)
	) name1604 (
		_w38_,
		_w106_,
		_w110_,
		_w1638_
	);
	LUT4 #(
		.INIT('h135f)
	) name1605 (
		_w56_,
		_w47_,
		_w259_,
		_w378_,
		_w1639_
	);
	LUT3 #(
		.INIT('h40)
	) name1606 (
		_w385_,
		_w1638_,
		_w1639_,
		_w1640_
	);
	LUT4 #(
		.INIT('h8000)
	) name1607 (
		_w1637_,
		_w1640_,
		_w1630_,
		_w1633_,
		_w1641_
	);
	LUT2 #(
		.INIT('h8)
	) name1608 (
		_w1627_,
		_w1641_,
		_w1642_
	);
	LUT4 #(
		.INIT('h135f)
	) name1609 (
		_w38_,
		_w59_,
		_w78_,
		_w430_,
		_w1643_
	);
	LUT4 #(
		.INIT('h0777)
	) name1610 (
		_w47_,
		_w72_,
		_w93_,
		_w166_,
		_w1644_
	);
	LUT4 #(
		.INIT('h135f)
	) name1611 (
		_w85_,
		_w46_,
		_w158_,
		_w378_,
		_w1645_
	);
	LUT3 #(
		.INIT('h80)
	) name1612 (
		_w1643_,
		_w1644_,
		_w1645_,
		_w1646_
	);
	LUT4 #(
		.INIT('h153f)
	) name1613 (
		_w110_,
		_w47_,
		_w259_,
		_w419_,
		_w1647_
	);
	LUT4 #(
		.INIT('h0777)
	) name1614 (
		_w122_,
		_w90_,
		_w65_,
		_w419_,
		_w1648_
	);
	LUT4 #(
		.INIT('h0777)
	) name1615 (
		_w110_,
		_w43_,
		_w44_,
		_w166_,
		_w1649_
	);
	LUT3 #(
		.INIT('h80)
	) name1616 (
		_w1648_,
		_w1649_,
		_w1647_,
		_w1650_
	);
	LUT3 #(
		.INIT('h1f)
	) name1617 (
		_w110_,
		_w41_,
		_w158_,
		_w1651_
	);
	LUT4 #(
		.INIT('h135f)
	) name1618 (
		_w110_,
		_w44_,
		_w259_,
		_w176_,
		_w1652_
	);
	LUT4 #(
		.INIT('h8000)
	) name1619 (
		_w997_,
		_w1530_,
		_w1651_,
		_w1652_,
		_w1653_
	);
	LUT3 #(
		.INIT('h80)
	) name1620 (
		_w1646_,
		_w1650_,
		_w1653_,
		_w1654_
	);
	LUT4 #(
		.INIT('h4000)
	) name1621 (
		_w197_,
		_w737_,
		_w804_,
		_w783_,
		_w1655_
	);
	LUT4 #(
		.INIT('h135f)
	) name1622 (
		_w59_,
		_w50_,
		_w43_,
		_w176_,
		_w1656_
	);
	LUT4 #(
		.INIT('h135f)
	) name1623 (
		_w38_,
		_w44_,
		_w166_,
		_w430_,
		_w1657_
	);
	LUT3 #(
		.INIT('h57)
	) name1624 (
		_w46_,
		_w201_,
		_w259_,
		_w1658_
	);
	LUT4 #(
		.INIT('h8000)
	) name1625 (
		_w829_,
		_w1656_,
		_w1657_,
		_w1658_,
		_w1659_
	);
	LUT4 #(
		.INIT('h8000)
	) name1626 (
		_w1115_,
		_w1120_,
		_w1655_,
		_w1659_,
		_w1660_
	);
	LUT4 #(
		.INIT('h8000)
	) name1627 (
		_w1627_,
		_w1641_,
		_w1654_,
		_w1660_,
		_w1661_
	);
	LUT2 #(
		.INIT('h8)
	) name1628 (
		_w1620_,
		_w1661_,
		_w1662_
	);
	LUT2 #(
		.INIT('h1)
	) name1629 (
		_w1607_,
		_w1662_,
		_w1663_
	);
	LUT4 #(
		.INIT('h153f)
	) name1630 (
		_w65_,
		_w44_,
		_w236_,
		_w158_,
		_w1664_
	);
	LUT3 #(
		.INIT('h80)
	) name1631 (
		_w1492_,
		_w1589_,
		_w1664_,
		_w1665_
	);
	LUT4 #(
		.INIT('h135f)
	) name1632 (
		_w38_,
		_w85_,
		_w43_,
		_w176_,
		_w1666_
	);
	LUT4 #(
		.INIT('h2000)
	) name1633 (
		_w364_,
		_w410_,
		_w1168_,
		_w1666_,
		_w1667_
	);
	LUT4 #(
		.INIT('h0777)
	) name1634 (
		_w52_,
		_w39_,
		_w65_,
		_w176_,
		_w1668_
	);
	LUT3 #(
		.INIT('h37)
	) name1635 (
		_w106_,
		_w52_,
		_w176_,
		_w1669_
	);
	LUT2 #(
		.INIT('h4)
	) name1636 (
		_w118_,
		_w1669_,
		_w1670_
	);
	LUT4 #(
		.INIT('h1000)
	) name1637 (
		_w118_,
		_w482_,
		_w1668_,
		_w1669_,
		_w1671_
	);
	LUT3 #(
		.INIT('h80)
	) name1638 (
		_w1665_,
		_w1667_,
		_w1671_,
		_w1672_
	);
	LUT4 #(
		.INIT('h135f)
	) name1639 (
		_w47_,
		_w50_,
		_w201_,
		_w430_,
		_w1673_
	);
	LUT4 #(
		.INIT('h0777)
	) name1640 (
		_w38_,
		_w39_,
		_w46_,
		_w184_,
		_w1674_
	);
	LUT2 #(
		.INIT('h8)
	) name1641 (
		_w1673_,
		_w1674_,
		_w1675_
	);
	LUT4 #(
		.INIT('h0777)
	) name1642 (
		_w122_,
		_w67_,
		_w93_,
		_w201_,
		_w1676_
	);
	LUT4 #(
		.INIT('h153f)
	) name1643 (
		_w122_,
		_w67_,
		_w39_,
		_w65_,
		_w1677_
	);
	LUT4 #(
		.INIT('h4000)
	) name1644 (
		_w129_,
		_w1181_,
		_w1676_,
		_w1677_,
		_w1678_
	);
	LUT4 #(
		.INIT('h0777)
	) name1645 (
		_w78_,
		_w56_,
		_w41_,
		_w236_,
		_w1679_
	);
	LUT3 #(
		.INIT('h40)
	) name1646 (
		_w258_,
		_w1205_,
		_w1679_,
		_w1680_
	);
	LUT4 #(
		.INIT('h135f)
	) name1647 (
		_w55_,
		_w50_,
		_w158_,
		_w419_,
		_w1681_
	);
	LUT4 #(
		.INIT('h135f)
	) name1648 (
		_w106_,
		_w85_,
		_w44_,
		_w236_,
		_w1682_
	);
	LUT3 #(
		.INIT('h37)
	) name1649 (
		_w106_,
		_w47_,
		_w176_,
		_w1683_
	);
	LUT3 #(
		.INIT('h80)
	) name1650 (
		_w1682_,
		_w1683_,
		_w1681_,
		_w1684_
	);
	LUT4 #(
		.INIT('h8000)
	) name1651 (
		_w1675_,
		_w1680_,
		_w1684_,
		_w1678_,
		_w1685_
	);
	LUT3 #(
		.INIT('h80)
	) name1652 (
		_w716_,
		_w1672_,
		_w1685_,
		_w1686_
	);
	LUT4 #(
		.INIT('h135f)
	) name1653 (
		_w122_,
		_w85_,
		_w59_,
		_w78_,
		_w1687_
	);
	LUT4 #(
		.INIT('h135f)
	) name1654 (
		_w122_,
		_w55_,
		_w93_,
		_w378_,
		_w1688_
	);
	LUT3 #(
		.INIT('h80)
	) name1655 (
		_w1551_,
		_w1688_,
		_w1687_,
		_w1689_
	);
	LUT4 #(
		.INIT('h4000)
	) name1656 (
		_w301_,
		_w759_,
		_w1318_,
		_w1437_,
		_w1690_
	);
	LUT2 #(
		.INIT('h8)
	) name1657 (
		_w1689_,
		_w1690_,
		_w1691_
	);
	LUT4 #(
		.INIT('h8000)
	) name1658 (
		_w716_,
		_w1672_,
		_w1685_,
		_w1691_,
		_w1692_
	);
	LUT4 #(
		.INIT('h153f)
	) name1659 (
		_w55_,
		_w52_,
		_w201_,
		_w236_,
		_w1693_
	);
	LUT3 #(
		.INIT('h1f)
	) name1660 (
		_w47_,
		_w44_,
		_w419_,
		_w1694_
	);
	LUT4 #(
		.INIT('h0777)
	) name1661 (
		_w122_,
		_w90_,
		_w44_,
		_w166_,
		_w1695_
	);
	LUT4 #(
		.INIT('h8000)
	) name1662 (
		_w168_,
		_w1695_,
		_w1693_,
		_w1694_,
		_w1696_
	);
	LUT4 #(
		.INIT('h153f)
	) name1663 (
		_w56_,
		_w47_,
		_w72_,
		_w158_,
		_w1697_
	);
	LUT4 #(
		.INIT('h8000)
	) name1664 (
		_w1541_,
		_w1542_,
		_w1624_,
		_w1697_,
		_w1698_
	);
	LUT2 #(
		.INIT('h8)
	) name1665 (
		_w1696_,
		_w1698_,
		_w1699_
	);
	LUT4 #(
		.INIT('h135f)
	) name1666 (
		_w52_,
		_w93_,
		_w378_,
		_w430_,
		_w1700_
	);
	LUT4 #(
		.INIT('h0777)
	) name1667 (
		_w106_,
		_w110_,
		_w46_,
		_w176_,
		_w1701_
	);
	LUT3 #(
		.INIT('h40)
	) name1668 (
		_w450_,
		_w1700_,
		_w1701_,
		_w1702_
	);
	LUT4 #(
		.INIT('h153f)
	) name1669 (
		_w38_,
		_w52_,
		_w78_,
		_w201_,
		_w1703_
	);
	LUT4 #(
		.INIT('h135f)
	) name1670 (
		_w56_,
		_w41_,
		_w72_,
		_w166_,
		_w1704_
	);
	LUT4 #(
		.INIT('h8000)
	) name1671 (
		_w641_,
		_w978_,
		_w1703_,
		_w1704_,
		_w1705_
	);
	LUT3 #(
		.INIT('h80)
	) name1672 (
		_w532_,
		_w1702_,
		_w1705_,
		_w1706_
	);
	LUT4 #(
		.INIT('h153f)
	) name1673 (
		_w52_,
		_w110_,
		_w39_,
		_w43_,
		_w1707_
	);
	LUT2 #(
		.INIT('h4)
	) name1674 (
		_w369_,
		_w1707_,
		_w1708_
	);
	LUT3 #(
		.INIT('h57)
	) name1675 (
		_w90_,
		_w236_,
		_w378_,
		_w1709_
	);
	LUT3 #(
		.INIT('h40)
	) name1676 (
		_w471_,
		_w1458_,
		_w1709_,
		_w1710_
	);
	LUT2 #(
		.INIT('h8)
	) name1677 (
		_w1708_,
		_w1710_,
		_w1711_
	);
	LUT4 #(
		.INIT('h0777)
	) name1678 (
		_w38_,
		_w72_,
		_w65_,
		_w184_,
		_w1712_
	);
	LUT3 #(
		.INIT('h57)
	) name1679 (
		_w78_,
		_w41_,
		_w46_,
		_w1713_
	);
	LUT4 #(
		.INIT('h4000)
	) name1680 (
		_w314_,
		_w391_,
		_w1713_,
		_w1712_,
		_w1714_
	);
	LUT4 #(
		.INIT('h153f)
	) name1681 (
		_w55_,
		_w41_,
		_w378_,
		_w430_,
		_w1715_
	);
	LUT4 #(
		.INIT('h8000)
	) name1682 (
		_w150_,
		_w408_,
		_w1099_,
		_w1715_,
		_w1716_
	);
	LUT4 #(
		.INIT('h153f)
	) name1683 (
		_w59_,
		_w93_,
		_w236_,
		_w166_,
		_w1717_
	);
	LUT4 #(
		.INIT('h0777)
	) name1684 (
		_w106_,
		_w67_,
		_w56_,
		_w39_,
		_w1718_
	);
	LUT4 #(
		.INIT('h153f)
	) name1685 (
		_w122_,
		_w110_,
		_w78_,
		_w56_,
		_w1719_
	);
	LUT3 #(
		.INIT('h80)
	) name1686 (
		_w1717_,
		_w1718_,
		_w1719_,
		_w1720_
	);
	LUT3 #(
		.INIT('h80)
	) name1687 (
		_w635_,
		_w649_,
		_w1180_,
		_w1721_
	);
	LUT4 #(
		.INIT('h8000)
	) name1688 (
		_w1720_,
		_w1721_,
		_w1714_,
		_w1716_,
		_w1722_
	);
	LUT4 #(
		.INIT('h8000)
	) name1689 (
		_w1699_,
		_w1706_,
		_w1711_,
		_w1722_,
		_w1723_
	);
	LUT2 #(
		.INIT('h8)
	) name1690 (
		_w1692_,
		_w1723_,
		_w1724_
	);
	LUT4 #(
		.INIT('h135f)
	) name1691 (
		_w55_,
		_w44_,
		_w184_,
		_w166_,
		_w1725_
	);
	LUT4 #(
		.INIT('h0777)
	) name1692 (
		_w85_,
		_w78_,
		_w41_,
		_w158_,
		_w1726_
	);
	LUT4 #(
		.INIT('h8000)
	) name1693 (
		_w843_,
		_w1683_,
		_w1725_,
		_w1726_,
		_w1727_
	);
	LUT4 #(
		.INIT('h153f)
	) name1694 (
		_w47_,
		_w41_,
		_w39_,
		_w166_,
		_w1728_
	);
	LUT4 #(
		.INIT('h153f)
	) name1695 (
		_w38_,
		_w110_,
		_w72_,
		_w43_,
		_w1729_
	);
	LUT4 #(
		.INIT('h4000)
	) name1696 (
		_w338_,
		_w637_,
		_w1729_,
		_w1728_,
		_w1730_
	);
	LUT2 #(
		.INIT('h8)
	) name1697 (
		_w1727_,
		_w1730_,
		_w1731_
	);
	LUT3 #(
		.INIT('h57)
	) name1698 (
		_w65_,
		_w236_,
		_w166_,
		_w1732_
	);
	LUT2 #(
		.INIT('h8)
	) name1699 (
		_w501_,
		_w1732_,
		_w1733_
	);
	LUT4 #(
		.INIT('h8000)
	) name1700 (
		_w521_,
		_w555_,
		_w697_,
		_w803_,
		_w1734_
	);
	LUT4 #(
		.INIT('h135f)
	) name1701 (
		_w85_,
		_w93_,
		_w201_,
		_w419_,
		_w1735_
	);
	LUT4 #(
		.INIT('h135f)
	) name1702 (
		_w38_,
		_w90_,
		_w176_,
		_w378_,
		_w1736_
	);
	LUT4 #(
		.INIT('h8000)
	) name1703 (
		_w580_,
		_w1276_,
		_w1736_,
		_w1735_,
		_w1737_
	);
	LUT4 #(
		.INIT('h135f)
	) name1704 (
		_w85_,
		_w59_,
		_w419_,
		_w378_,
		_w1738_
	);
	LUT3 #(
		.INIT('h80)
	) name1705 (
		_w863_,
		_w1154_,
		_w1738_,
		_w1739_
	);
	LUT4 #(
		.INIT('h8000)
	) name1706 (
		_w1737_,
		_w1733_,
		_w1739_,
		_w1734_,
		_w1740_
	);
	LUT4 #(
		.INIT('h153f)
	) name1707 (
		_w52_,
		_w50_,
		_w158_,
		_w259_,
		_w1741_
	);
	LUT3 #(
		.INIT('h80)
	) name1708 (
		_w1731_,
		_w1740_,
		_w1741_,
		_w1742_
	);
	LUT4 #(
		.INIT('h4000)
	) name1709 (
		_w334_,
		_w538_,
		_w563_,
		_w886_,
		_w1743_
	);
	LUT4 #(
		.INIT('h135f)
	) name1710 (
		_w93_,
		_w65_,
		_w166_,
		_w259_,
		_w1744_
	);
	LUT4 #(
		.INIT('h0200)
	) name1711 (
		_w361_,
		_w406_,
		_w444_,
		_w1744_,
		_w1745_
	);
	LUT4 #(
		.INIT('h0777)
	) name1712 (
		_w106_,
		_w55_,
		_w46_,
		_w201_,
		_w1746_
	);
	LUT3 #(
		.INIT('h40)
	) name1713 (
		_w197_,
		_w1019_,
		_w1746_,
		_w1747_
	);
	LUT4 #(
		.INIT('h0777)
	) name1714 (
		_w78_,
		_w47_,
		_w50_,
		_w430_,
		_w1748_
	);
	LUT3 #(
		.INIT('h80)
	) name1715 (
		_w918_,
		_w1047_,
		_w1748_,
		_w1749_
	);
	LUT4 #(
		.INIT('h8000)
	) name1716 (
		_w1747_,
		_w1749_,
		_w1743_,
		_w1745_,
		_w1750_
	);
	LUT2 #(
		.INIT('h8)
	) name1717 (
		_w1261_,
		_w1750_,
		_w1751_
	);
	LUT4 #(
		.INIT('h0777)
	) name1718 (
		_w67_,
		_w78_,
		_w46_,
		_w259_,
		_w1752_
	);
	LUT4 #(
		.INIT('h153f)
	) name1719 (
		_w85_,
		_w110_,
		_w184_,
		_w166_,
		_w1753_
	);
	LUT4 #(
		.INIT('h153f)
	) name1720 (
		_w56_,
		_w43_,
		_w93_,
		_w419_,
		_w1754_
	);
	LUT3 #(
		.INIT('h80)
	) name1721 (
		_w1753_,
		_w1754_,
		_w1752_,
		_w1755_
	);
	LUT4 #(
		.INIT('h4000)
	) name1722 (
		_w209_,
		_w274_,
		_w1190_,
		_w1717_,
		_w1756_
	);
	LUT3 #(
		.INIT('h80)
	) name1723 (
		_w599_,
		_w1755_,
		_w1756_,
		_w1757_
	);
	LUT4 #(
		.INIT('h135f)
	) name1724 (
		_w47_,
		_w41_,
		_w72_,
		_w201_,
		_w1758_
	);
	LUT4 #(
		.INIT('h153f)
	) name1725 (
		_w38_,
		_w55_,
		_w158_,
		_w378_,
		_w1759_
	);
	LUT4 #(
		.INIT('h8000)
	) name1726 (
		_w662_,
		_w790_,
		_w1758_,
		_w1759_,
		_w1760_
	);
	LUT4 #(
		.INIT('h135f)
	) name1727 (
		_w106_,
		_w52_,
		_w67_,
		_w158_,
		_w1761_
	);
	LUT4 #(
		.INIT('h135f)
	) name1728 (
		_w38_,
		_w67_,
		_w39_,
		_w184_,
		_w1762_
	);
	LUT4 #(
		.INIT('h2000)
	) name1729 (
		_w68_,
		_w295_,
		_w1761_,
		_w1762_,
		_w1763_
	);
	LUT2 #(
		.INIT('h8)
	) name1730 (
		_w1760_,
		_w1763_,
		_w1764_
	);
	LUT4 #(
		.INIT('h0777)
	) name1731 (
		_w106_,
		_w85_,
		_w72_,
		_w65_,
		_w1765_
	);
	LUT4 #(
		.INIT('h135f)
	) name1732 (
		_w90_,
		_w50_,
		_w184_,
		_w166_,
		_w1766_
	);
	LUT4 #(
		.INIT('h153f)
	) name1733 (
		_w55_,
		_w59_,
		_w419_,
		_w430_,
		_w1767_
	);
	LUT3 #(
		.INIT('h80)
	) name1734 (
		_w1765_,
		_w1766_,
		_w1767_,
		_w1768_
	);
	LUT3 #(
		.INIT('h80)
	) name1735 (
		_w1037_,
		_w1182_,
		_w1278_,
		_w1769_
	);
	LUT3 #(
		.INIT('h80)
	) name1736 (
		_w907_,
		_w1768_,
		_w1769_,
		_w1770_
	);
	LUT3 #(
		.INIT('h80)
	) name1737 (
		_w1757_,
		_w1764_,
		_w1770_,
		_w1771_
	);
	LUT3 #(
		.INIT('h80)
	) name1738 (
		_w1751_,
		_w1742_,
		_w1771_,
		_w1772_
	);
	LUT2 #(
		.INIT('h1)
	) name1739 (
		_w1724_,
		_w1772_,
		_w1773_
	);
	LUT4 #(
		.INIT('h153f)
	) name1740 (
		_w38_,
		_w46_,
		_w236_,
		_w419_,
		_w1774_
	);
	LUT3 #(
		.INIT('h40)
	) name1741 (
		_w220_,
		_w479_,
		_w1774_,
		_w1775_
	);
	LUT4 #(
		.INIT('h153f)
	) name1742 (
		_w67_,
		_w56_,
		_w201_,
		_w166_,
		_w1776_
	);
	LUT4 #(
		.INIT('h0777)
	) name1743 (
		_w122_,
		_w93_,
		_w46_,
		_w378_,
		_w1777_
	);
	LUT4 #(
		.INIT('h0777)
	) name1744 (
		_w122_,
		_w47_,
		_w72_,
		_w50_,
		_w1778_
	);
	LUT4 #(
		.INIT('h4000)
	) name1745 (
		_w320_,
		_w1776_,
		_w1777_,
		_w1778_,
		_w1779_
	);
	LUT3 #(
		.INIT('h80)
	) name1746 (
		_w804_,
		_w864_,
		_w1587_,
		_w1780_
	);
	LUT3 #(
		.INIT('h80)
	) name1747 (
		_w1779_,
		_w1775_,
		_w1780_,
		_w1781_
	);
	LUT2 #(
		.INIT('h4)
	) name1748 (
		_w146_,
		_w1416_,
		_w1782_
	);
	LUT4 #(
		.INIT('h135f)
	) name1749 (
		_w122_,
		_w78_,
		_w41_,
		_w93_,
		_w1783_
	);
	LUT4 #(
		.INIT('h135f)
	) name1750 (
		_w59_,
		_w47_,
		_w43_,
		_w236_,
		_w1784_
	);
	LUT4 #(
		.INIT('h153f)
	) name1751 (
		_w55_,
		_w47_,
		_w166_,
		_w378_,
		_w1785_
	);
	LUT3 #(
		.INIT('h80)
	) name1752 (
		_w1784_,
		_w1785_,
		_w1783_,
		_w1786_
	);
	LUT2 #(
		.INIT('h8)
	) name1753 (
		_w1782_,
		_w1786_,
		_w1787_
	);
	LUT4 #(
		.INIT('h135f)
	) name1754 (
		_w85_,
		_w47_,
		_w201_,
		_w158_,
		_w1788_
	);
	LUT4 #(
		.INIT('h1000)
	) name1755 (
		_w129_,
		_w440_,
		_w1676_,
		_w1788_,
		_w1789_
	);
	LUT4 #(
		.INIT('h153f)
	) name1756 (
		_w90_,
		_w72_,
		_w44_,
		_w419_,
		_w1790_
	);
	LUT4 #(
		.INIT('h0777)
	) name1757 (
		_w122_,
		_w52_,
		_w50_,
		_w430_,
		_w1791_
	);
	LUT4 #(
		.INIT('h153f)
	) name1758 (
		_w55_,
		_w50_,
		_w43_,
		_w158_,
		_w1792_
	);
	LUT4 #(
		.INIT('h4000)
	) name1759 (
		_w83_,
		_w1790_,
		_w1791_,
		_w1792_,
		_w1793_
	);
	LUT4 #(
		.INIT('h8000)
	) name1760 (
		_w1394_,
		_w1396_,
		_w1789_,
		_w1793_,
		_w1794_
	);
	LUT3 #(
		.INIT('h80)
	) name1761 (
		_w1787_,
		_w1781_,
		_w1794_,
		_w1795_
	);
	LUT4 #(
		.INIT('h8000)
	) name1762 (
		_w1261_,
		_w1271_,
		_w1441_,
		_w1453_,
		_w1796_
	);
	LUT2 #(
		.INIT('h8)
	) name1763 (
		_w1795_,
		_w1796_,
		_w1797_
	);
	LUT4 #(
		.INIT('h153f)
	) name1764 (
		_w52_,
		_w65_,
		_w201_,
		_w176_,
		_w1798_
	);
	LUT3 #(
		.INIT('h80)
	) name1765 (
		_w749_,
		_w762_,
		_w1798_,
		_w1799_
	);
	LUT4 #(
		.INIT('h135f)
	) name1766 (
		_w41_,
		_w44_,
		_w184_,
		_w419_,
		_w1800_
	);
	LUT3 #(
		.INIT('h40)
	) name1767 (
		_w141_,
		_w924_,
		_w1800_,
		_w1801_
	);
	LUT4 #(
		.INIT('h153f)
	) name1768 (
		_w59_,
		_w50_,
		_w176_,
		_w419_,
		_w1802_
	);
	LUT2 #(
		.INIT('h8)
	) name1769 (
		_w181_,
		_w1802_,
		_w1803_
	);
	LUT4 #(
		.INIT('h8000)
	) name1770 (
		_w887_,
		_w1222_,
		_w1483_,
		_w1586_,
		_w1804_
	);
	LUT3 #(
		.INIT('h80)
	) name1771 (
		_w1801_,
		_w1803_,
		_w1804_,
		_w1805_
	);
	LUT4 #(
		.INIT('h153f)
	) name1772 (
		_w85_,
		_w56_,
		_w201_,
		_w158_,
		_w1806_
	);
	LUT2 #(
		.INIT('h4)
	) name1773 (
		_w455_,
		_w1806_,
		_w1807_
	);
	LUT4 #(
		.INIT('h135f)
	) name1774 (
		_w110_,
		_w47_,
		_w43_,
		_w201_,
		_w1808_
	);
	LUT4 #(
		.INIT('h4000)
	) name1775 (
		_w282_,
		_w717_,
		_w718_,
		_w1808_,
		_w1809_
	);
	LUT4 #(
		.INIT('h153f)
	) name1776 (
		_w110_,
		_w78_,
		_w44_,
		_w176_,
		_w1810_
	);
	LUT4 #(
		.INIT('h135f)
	) name1777 (
		_w122_,
		_w55_,
		_w56_,
		_w201_,
		_w1811_
	);
	LUT3 #(
		.INIT('h80)
	) name1778 (
		_w1248_,
		_w1811_,
		_w1810_,
		_w1812_
	);
	LUT4 #(
		.INIT('h153f)
	) name1779 (
		_w122_,
		_w106_,
		_w59_,
		_w47_,
		_w1813_
	);
	LUT4 #(
		.INIT('h135f)
	) name1780 (
		_w106_,
		_w47_,
		_w41_,
		_w39_,
		_w1814_
	);
	LUT4 #(
		.INIT('h8000)
	) name1781 (
		_w125_,
		_w1281_,
		_w1813_,
		_w1814_,
		_w1815_
	);
	LUT4 #(
		.INIT('h8000)
	) name1782 (
		_w1807_,
		_w1812_,
		_w1815_,
		_w1809_,
		_w1816_
	);
	LUT2 #(
		.INIT('h8)
	) name1783 (
		_w1805_,
		_w1816_,
		_w1817_
	);
	LUT4 #(
		.INIT('h0777)
	) name1784 (
		_w90_,
		_w72_,
		_w39_,
		_w46_,
		_w1818_
	);
	LUT3 #(
		.INIT('h80)
	) name1785 (
		_w1165_,
		_w1190_,
		_w1818_,
		_w1819_
	);
	LUT2 #(
		.INIT('h8)
	) name1786 (
		_w1013_,
		_w1374_,
		_w1820_
	);
	LUT3 #(
		.INIT('h57)
	) name1787 (
		_w67_,
		_w184_,
		_w158_,
		_w1821_
	);
	LUT4 #(
		.INIT('h1000)
	) name1788 (
		_w451_,
		_w477_,
		_w726_,
		_w1821_,
		_w1822_
	);
	LUT3 #(
		.INIT('h80)
	) name1789 (
		_w1820_,
		_w1819_,
		_w1822_,
		_w1823_
	);
	LUT4 #(
		.INIT('h153f)
	) name1790 (
		_w110_,
		_w67_,
		_w259_,
		_w378_,
		_w1824_
	);
	LUT2 #(
		.INIT('h4)
	) name1791 (
		_w385_,
		_w1824_,
		_w1825_
	);
	LUT4 #(
		.INIT('h135f)
	) name1792 (
		_w67_,
		_w93_,
		_w166_,
		_w430_,
		_w1826_
	);
	LUT4 #(
		.INIT('h135f)
	) name1793 (
		_w56_,
		_w39_,
		_w43_,
		_w65_,
		_w1827_
	);
	LUT4 #(
		.INIT('h153f)
	) name1794 (
		_w47_,
		_w93_,
		_w158_,
		_w176_,
		_w1828_
	);
	LUT3 #(
		.INIT('h80)
	) name1795 (
		_w1826_,
		_w1827_,
		_w1828_,
		_w1829_
	);
	LUT2 #(
		.INIT('h8)
	) name1796 (
		_w1825_,
		_w1829_,
		_w1830_
	);
	LUT4 #(
		.INIT('h8000)
	) name1797 (
		_w538_,
		_w668_,
		_w737_,
		_w991_,
		_w1831_
	);
	LUT3 #(
		.INIT('h1f)
	) name1798 (
		_w55_,
		_w85_,
		_w259_,
		_w1832_
	);
	LUT4 #(
		.INIT('h0777)
	) name1799 (
		_w106_,
		_w90_,
		_w65_,
		_w430_,
		_w1833_
	);
	LUT4 #(
		.INIT('h153f)
	) name1800 (
		_w59_,
		_w72_,
		_w46_,
		_w158_,
		_w1834_
	);
	LUT4 #(
		.INIT('h8000)
	) name1801 (
		_w216_,
		_w1834_,
		_w1832_,
		_w1833_,
		_w1835_
	);
	LUT3 #(
		.INIT('h20)
	) name1802 (
		_w198_,
		_w462_,
		_w1493_,
		_w1836_
	);
	LUT4 #(
		.INIT('h135f)
	) name1803 (
		_w38_,
		_w41_,
		_w43_,
		_w378_,
		_w1837_
	);
	LUT3 #(
		.INIT('h80)
	) name1804 (
		_w1061_,
		_w1216_,
		_w1837_,
		_w1838_
	);
	LUT4 #(
		.INIT('h8000)
	) name1805 (
		_w1836_,
		_w1838_,
		_w1831_,
		_w1835_,
		_w1839_
	);
	LUT3 #(
		.INIT('h80)
	) name1806 (
		_w1830_,
		_w1823_,
		_w1839_,
		_w1840_
	);
	LUT3 #(
		.INIT('h80)
	) name1807 (
		_w1817_,
		_w1799_,
		_w1840_,
		_w1841_
	);
	LUT2 #(
		.INIT('h1)
	) name1808 (
		_w1797_,
		_w1841_,
		_w1842_
	);
	LUT4 #(
		.INIT('h153f)
	) name1809 (
		_w122_,
		_w52_,
		_w72_,
		_w46_,
		_w1843_
	);
	LUT4 #(
		.INIT('h153f)
	) name1810 (
		_w41_,
		_w93_,
		_w158_,
		_w419_,
		_w1844_
	);
	LUT4 #(
		.INIT('h0777)
	) name1811 (
		_w106_,
		_w85_,
		_w39_,
		_w50_,
		_w1845_
	);
	LUT4 #(
		.INIT('h8000)
	) name1812 (
		_w1174_,
		_w1843_,
		_w1844_,
		_w1845_,
		_w1846_
	);
	LUT4 #(
		.INIT('h135f)
	) name1813 (
		_w85_,
		_w56_,
		_w176_,
		_w430_,
		_w1847_
	);
	LUT2 #(
		.INIT('h4)
	) name1814 (
		_w432_,
		_w1847_,
		_w1848_
	);
	LUT4 #(
		.INIT('h0777)
	) name1815 (
		_w55_,
		_w78_,
		_w44_,
		_w166_,
		_w1849_
	);
	LUT4 #(
		.INIT('h4000)
	) name1816 (
		_w83_,
		_w962_,
		_w1790_,
		_w1849_,
		_w1850_
	);
	LUT3 #(
		.INIT('h80)
	) name1817 (
		_w1848_,
		_w1846_,
		_w1850_,
		_w1851_
	);
	LUT4 #(
		.INIT('h153f)
	) name1818 (
		_w38_,
		_w59_,
		_w201_,
		_w236_,
		_w1852_
	);
	LUT4 #(
		.INIT('h153f)
	) name1819 (
		_w90_,
		_w41_,
		_w39_,
		_w378_,
		_w1853_
	);
	LUT2 #(
		.INIT('h8)
	) name1820 (
		_w1852_,
		_w1853_,
		_w1854_
	);
	LUT4 #(
		.INIT('h135f)
	) name1821 (
		_w38_,
		_w106_,
		_w78_,
		_w46_,
		_w1855_
	);
	LUT4 #(
		.INIT('h0200)
	) name1822 (
		_w81_,
		_w193_,
		_w441_,
		_w1855_,
		_w1856_
	);
	LUT2 #(
		.INIT('h8)
	) name1823 (
		_w1854_,
		_w1856_,
		_w1857_
	);
	LUT4 #(
		.INIT('h135f)
	) name1824 (
		_w85_,
		_w90_,
		_w184_,
		_w166_,
		_w1858_
	);
	LUT4 #(
		.INIT('h8000)
	) name1825 (
		_w1273_,
		_w1374_,
		_w1550_,
		_w1858_,
		_w1859_
	);
	LUT3 #(
		.INIT('h40)
	) name1826 (
		_w141_,
		_w384_,
		_w942_,
		_w1860_
	);
	LUT4 #(
		.INIT('h4000)
	) name1827 (
		_w128_,
		_w112_,
		_w139_,
		_w309_,
		_w1861_
	);
	LUT4 #(
		.INIT('h8000)
	) name1828 (
		_w733_,
		_w1860_,
		_w1861_,
		_w1859_,
		_w1862_
	);
	LUT3 #(
		.INIT('h80)
	) name1829 (
		_w1851_,
		_w1857_,
		_w1862_,
		_w1863_
	);
	LUT4 #(
		.INIT('h8000)
	) name1830 (
		_w793_,
		_w768_,
		_w909_,
		_w1437_,
		_w1864_
	);
	LUT4 #(
		.INIT('h0777)
	) name1831 (
		_w122_,
		_w44_,
		_w46_,
		_w430_,
		_w1865_
	);
	LUT4 #(
		.INIT('h0777)
	) name1832 (
		_w85_,
		_w43_,
		_w44_,
		_w158_,
		_w1866_
	);
	LUT4 #(
		.INIT('h0777)
	) name1833 (
		_w52_,
		_w39_,
		_w93_,
		_w166_,
		_w1867_
	);
	LUT4 #(
		.INIT('h8000)
	) name1834 (
		_w534_,
		_w1865_,
		_w1866_,
		_w1867_,
		_w1868_
	);
	LUT2 #(
		.INIT('h8)
	) name1835 (
		_w1864_,
		_w1868_,
		_w1869_
	);
	LUT3 #(
		.INIT('h10)
	) name1836 (
		_w359_,
		_w437_,
		_w1021_,
		_w1870_
	);
	LUT4 #(
		.INIT('h0777)
	) name1837 (
		_w106_,
		_w41_,
		_w65_,
		_w259_,
		_w1871_
	);
	LUT3 #(
		.INIT('h80)
	) name1838 (
		_w1427_,
		_w1664_,
		_w1871_,
		_w1872_
	);
	LUT3 #(
		.INIT('h80)
	) name1839 (
		_w1680_,
		_w1870_,
		_w1872_,
		_w1873_
	);
	LUT2 #(
		.INIT('h8)
	) name1840 (
		_w1869_,
		_w1873_,
		_w1874_
	);
	LUT4 #(
		.INIT('h8000)
	) name1841 (
		_w1612_,
		_w1619_,
		_w1869_,
		_w1873_,
		_w1875_
	);
	LUT2 #(
		.INIT('h8)
	) name1842 (
		_w1863_,
		_w1875_,
		_w1876_
	);
	LUT4 #(
		.INIT('h135f)
	) name1843 (
		_w122_,
		_w39_,
		_w65_,
		_w46_,
		_w1877_
	);
	LUT4 #(
		.INIT('h135f)
	) name1844 (
		_w85_,
		_w93_,
		_w166_,
		_w259_,
		_w1878_
	);
	LUT4 #(
		.INIT('h0777)
	) name1845 (
		_w122_,
		_w85_,
		_w46_,
		_w201_,
		_w1879_
	);
	LUT4 #(
		.INIT('h8000)
	) name1846 (
		_w1410_,
		_w1877_,
		_w1878_,
		_w1879_,
		_w1880_
	);
	LUT2 #(
		.INIT('h4)
	) name1847 (
		_w462_,
		_w1360_,
		_w1881_
	);
	LUT3 #(
		.INIT('h37)
	) name1848 (
		_w78_,
		_w41_,
		_w176_,
		_w1882_
	);
	LUT4 #(
		.INIT('h4000)
	) name1849 (
		_w426_,
		_w817_,
		_w876_,
		_w1882_,
		_w1883_
	);
	LUT3 #(
		.INIT('h80)
	) name1850 (
		_w1881_,
		_w1880_,
		_w1883_,
		_w1884_
	);
	LUT4 #(
		.INIT('h0777)
	) name1851 (
		_w56_,
		_w72_,
		_w46_,
		_w158_,
		_w1885_
	);
	LUT4 #(
		.INIT('h135f)
	) name1852 (
		_w85_,
		_w110_,
		_w236_,
		_w419_,
		_w1886_
	);
	LUT4 #(
		.INIT('h8000)
	) name1853 (
		_w309_,
		_w403_,
		_w1885_,
		_w1886_,
		_w1887_
	);
	LUT4 #(
		.INIT('h135f)
	) name1854 (
		_w106_,
		_w55_,
		_w93_,
		_w201_,
		_w1888_
	);
	LUT4 #(
		.INIT('h1000)
	) name1855 (
		_w40_,
		_w189_,
		_w191_,
		_w1888_,
		_w1889_
	);
	LUT2 #(
		.INIT('h8)
	) name1856 (
		_w1887_,
		_w1889_,
		_w1890_
	);
	LUT4 #(
		.INIT('h135f)
	) name1857 (
		_w122_,
		_w43_,
		_w93_,
		_w46_,
		_w1891_
	);
	LUT4 #(
		.INIT('h135f)
	) name1858 (
		_w110_,
		_w56_,
		_w184_,
		_w430_,
		_w1892_
	);
	LUT3 #(
		.INIT('h80)
	) name1859 (
		_w1126_,
		_w1891_,
		_w1892_,
		_w1893_
	);
	LUT4 #(
		.INIT('h135f)
	) name1860 (
		_w110_,
		_w90_,
		_w72_,
		_w201_,
		_w1894_
	);
	LUT3 #(
		.INIT('h37)
	) name1861 (
		_w106_,
		_w67_,
		_w176_,
		_w1895_
	);
	LUT3 #(
		.INIT('h80)
	) name1862 (
		_w1676_,
		_w1895_,
		_w1894_,
		_w1896_
	);
	LUT3 #(
		.INIT('h80)
	) name1863 (
		_w1424_,
		_w1893_,
		_w1896_,
		_w1897_
	);
	LUT3 #(
		.INIT('h80)
	) name1864 (
		_w1884_,
		_w1890_,
		_w1897_,
		_w1898_
	);
	LUT4 #(
		.INIT('h2000)
	) name1865 (
		_w198_,
		_w398_,
		_w1401_,
		_w1494_,
		_w1899_
	);
	LUT4 #(
		.INIT('h8000)
	) name1866 (
		_w651_,
		_w750_,
		_w1138_,
		_w1333_,
		_w1900_
	);
	LUT4 #(
		.INIT('h153f)
	) name1867 (
		_w85_,
		_w78_,
		_w56_,
		_w201_,
		_w1901_
	);
	LUT4 #(
		.INIT('h0200)
	) name1868 (
		_w254_,
		_w397_,
		_w440_,
		_w1901_,
		_w1902_
	);
	LUT3 #(
		.INIT('h80)
	) name1869 (
		_w1899_,
		_w1900_,
		_w1902_,
		_w1903_
	);
	LUT4 #(
		.INIT('h135f)
	) name1870 (
		_w59_,
		_w50_,
		_w259_,
		_w378_,
		_w1904_
	);
	LUT4 #(
		.INIT('h153f)
	) name1871 (
		_w38_,
		_w110_,
		_w236_,
		_w378_,
		_w1905_
	);
	LUT3 #(
		.INIT('h80)
	) name1872 (
		_w1113_,
		_w1905_,
		_w1904_,
		_w1906_
	);
	LUT4 #(
		.INIT('h135f)
	) name1873 (
		_w110_,
		_w67_,
		_w78_,
		_w166_,
		_w1907_
	);
	LUT4 #(
		.INIT('h135f)
	) name1874 (
		_w38_,
		_w122_,
		_w106_,
		_w52_,
		_w1908_
	);
	LUT4 #(
		.INIT('h4000)
	) name1875 (
		_w413_,
		_w843_,
		_w1908_,
		_w1907_,
		_w1909_
	);
	LUT4 #(
		.INIT('h135f)
	) name1876 (
		_w38_,
		_w41_,
		_w201_,
		_w236_,
		_w1910_
	);
	LUT4 #(
		.INIT('h0777)
	) name1877 (
		_w110_,
		_w43_,
		_w46_,
		_w184_,
		_w1911_
	);
	LUT2 #(
		.INIT('h8)
	) name1878 (
		_w1910_,
		_w1911_,
		_w1912_
	);
	LUT4 #(
		.INIT('h1000)
	) name1879 (
		_w226_,
		_w294_,
		_w538_,
		_w1211_,
		_w1913_
	);
	LUT4 #(
		.INIT('h8000)
	) name1880 (
		_w1912_,
		_w1906_,
		_w1909_,
		_w1913_,
		_w1914_
	);
	LUT4 #(
		.INIT('h135f)
	) name1881 (
		_w50_,
		_w93_,
		_w184_,
		_w430_,
		_w1915_
	);
	LUT2 #(
		.INIT('h8)
	) name1882 (
		_w1359_,
		_w1915_,
		_w1916_
	);
	LUT4 #(
		.INIT('h4000)
	) name1883 (
		_w206_,
		_w824_,
		_w1656_,
		_w1657_,
		_w1917_
	);
	LUT2 #(
		.INIT('h8)
	) name1884 (
		_w1916_,
		_w1917_,
		_w1918_
	);
	LUT4 #(
		.INIT('h135f)
	) name1885 (
		_w59_,
		_w50_,
		_w236_,
		_w259_,
		_w1919_
	);
	LUT3 #(
		.INIT('h1f)
	) name1886 (
		_w67_,
		_w44_,
		_w419_,
		_w1920_
	);
	LUT4 #(
		.INIT('h135f)
	) name1887 (
		_w44_,
		_w46_,
		_w176_,
		_w419_,
		_w1921_
	);
	LUT4 #(
		.INIT('h153f)
	) name1888 (
		_w52_,
		_w46_,
		_w236_,
		_w166_,
		_w1922_
	);
	LUT4 #(
		.INIT('h8000)
	) name1889 (
		_w1921_,
		_w1922_,
		_w1919_,
		_w1920_,
		_w1923_
	);
	LUT4 #(
		.INIT('h153f)
	) name1890 (
		_w55_,
		_w50_,
		_w166_,
		_w158_,
		_w1924_
	);
	LUT3 #(
		.INIT('h80)
	) name1891 (
		_w1334_,
		_w1783_,
		_w1924_,
		_w1925_
	);
	LUT4 #(
		.INIT('h8000)
	) name1892 (
		_w768_,
		_w789_,
		_w950_,
		_w1257_,
		_w1926_
	);
	LUT3 #(
		.INIT('h80)
	) name1893 (
		_w1923_,
		_w1925_,
		_w1926_,
		_w1927_
	);
	LUT4 #(
		.INIT('h8000)
	) name1894 (
		_w1903_,
		_w1914_,
		_w1918_,
		_w1927_,
		_w1928_
	);
	LUT2 #(
		.INIT('h8)
	) name1895 (
		_w1898_,
		_w1928_,
		_w1929_
	);
	LUT4 #(
		.INIT('h0777)
	) name1896 (
		_w1863_,
		_w1875_,
		_w1898_,
		_w1928_,
		_w1930_
	);
	LUT4 #(
		.INIT('h135f)
	) name1897 (
		_w55_,
		_w93_,
		_w201_,
		_w430_,
		_w1931_
	);
	LUT2 #(
		.INIT('h8)
	) name1898 (
		_w1910_,
		_w1931_,
		_w1932_
	);
	LUT4 #(
		.INIT('h4000)
	) name1899 (
		_w230_,
		_w944_,
		_w1359_,
		_w1506_,
		_w1933_
	);
	LUT2 #(
		.INIT('h8)
	) name1900 (
		_w1932_,
		_w1933_,
		_w1934_
	);
	LUT4 #(
		.INIT('h135f)
	) name1901 (
		_w122_,
		_w90_,
		_w50_,
		_w236_,
		_w1935_
	);
	LUT4 #(
		.INIT('h135f)
	) name1902 (
		_w85_,
		_w67_,
		_w419_,
		_w430_,
		_w1936_
	);
	LUT3 #(
		.INIT('h80)
	) name1903 (
		_w1179_,
		_w1936_,
		_w1935_,
		_w1937_
	);
	LUT3 #(
		.INIT('h80)
	) name1904 (
		_w1436_,
		_w1779_,
		_w1937_,
		_w1938_
	);
	LUT2 #(
		.INIT('h8)
	) name1905 (
		_w1934_,
		_w1938_,
		_w1939_
	);
	LUT3 #(
		.INIT('h40)
	) name1906 (
		_w209_,
		_w260_,
		_w403_,
		_w1940_
	);
	LUT4 #(
		.INIT('h4000)
	) name1907 (
		_w167_,
		_w760_,
		_w1791_,
		_w1792_,
		_w1941_
	);
	LUT3 #(
		.INIT('h80)
	) name1908 (
		_w302_,
		_w584_,
		_w1184_,
		_w1942_
	);
	LUT3 #(
		.INIT('h80)
	) name1909 (
		_w1941_,
		_w1942_,
		_w1940_,
		_w1943_
	);
	LUT3 #(
		.INIT('h80)
	) name1910 (
		_w997_,
		_w1416_,
		_w1664_,
		_w1944_
	);
	LUT4 #(
		.INIT('h153f)
	) name1911 (
		_w90_,
		_w39_,
		_w46_,
		_w166_,
		_w1945_
	);
	LUT4 #(
		.INIT('h135f)
	) name1912 (
		_w52_,
		_w110_,
		_w78_,
		_w378_,
		_w1946_
	);
	LUT4 #(
		.INIT('h4000)
	) name1913 (
		_w339_,
		_w906_,
		_w1945_,
		_w1946_,
		_w1947_
	);
	LUT4 #(
		.INIT('h8000)
	) name1914 (
		_w1065_,
		_w1105_,
		_w1944_,
		_w1947_,
		_w1948_
	);
	LUT4 #(
		.INIT('h8000)
	) name1915 (
		_w1934_,
		_w1938_,
		_w1943_,
		_w1948_,
		_w1949_
	);
	LUT2 #(
		.INIT('h8)
	) name1916 (
		_w1501_,
		_w1949_,
		_w1950_
	);
	LUT4 #(
		.INIT('h135f)
	) name1917 (
		_w122_,
		_w85_,
		_w93_,
		_w419_,
		_w1951_
	);
	LUT2 #(
		.INIT('h8)
	) name1918 (
		_w767_,
		_w1951_,
		_w1952_
	);
	LUT4 #(
		.INIT('h135f)
	) name1919 (
		_w67_,
		_w93_,
		_w184_,
		_w378_,
		_w1953_
	);
	LUT4 #(
		.INIT('h8000)
	) name1920 (
		_w1089_,
		_w1127_,
		_w1879_,
		_w1953_,
		_w1954_
	);
	LUT3 #(
		.INIT('h80)
	) name1921 (
		_w1331_,
		_w1952_,
		_w1954_,
		_w1955_
	);
	LUT4 #(
		.INIT('h135f)
	) name1922 (
		_w110_,
		_w56_,
		_w201_,
		_w419_,
		_w1956_
	);
	LUT3 #(
		.INIT('h80)
	) name1923 (
		_w867_,
		_w1112_,
		_w1956_,
		_w1957_
	);
	LUT4 #(
		.INIT('h0400)
	) name1924 (
		_w239_,
		_w342_,
		_w455_,
		_w1806_,
		_w1958_
	);
	LUT2 #(
		.INIT('h8)
	) name1925 (
		_w1957_,
		_w1958_,
		_w1959_
	);
	LUT4 #(
		.INIT('h8000)
	) name1926 (
		_w150_,
		_w1147_,
		_w1148_,
		_w1715_,
		_w1960_
	);
	LUT4 #(
		.INIT('h135f)
	) name1927 (
		_w56_,
		_w41_,
		_w184_,
		_w259_,
		_w1961_
	);
	LUT4 #(
		.INIT('h153f)
	) name1928 (
		_w110_,
		_w56_,
		_w236_,
		_w166_,
		_w1962_
	);
	LUT4 #(
		.INIT('h135f)
	) name1929 (
		_w85_,
		_w46_,
		_w259_,
		_w176_,
		_w1963_
	);
	LUT2 #(
		.INIT('h8)
	) name1930 (
		_w1962_,
		_w1963_,
		_w1964_
	);
	LUT4 #(
		.INIT('h8000)
	) name1931 (
		_w902_,
		_w1961_,
		_w1962_,
		_w1963_,
		_w1965_
	);
	LUT4 #(
		.INIT('h0777)
	) name1932 (
		_w122_,
		_w90_,
		_w47_,
		_w184_,
		_w1966_
	);
	LUT3 #(
		.INIT('h1f)
	) name1933 (
		_w85_,
		_w59_,
		_w184_,
		_w1967_
	);
	LUT4 #(
		.INIT('h8000)
	) name1934 (
		_w663_,
		_w1844_,
		_w1967_,
		_w1966_,
		_w1968_
	);
	LUT4 #(
		.INIT('h153f)
	) name1935 (
		_w110_,
		_w46_,
		_w184_,
		_w378_,
		_w1969_
	);
	LUT4 #(
		.INIT('h135f)
	) name1936 (
		_w59_,
		_w50_,
		_w419_,
		_w430_,
		_w1970_
	);
	LUT4 #(
		.INIT('h4000)
	) name1937 (
		_w468_,
		_w882_,
		_w1969_,
		_w1970_,
		_w1971_
	);
	LUT4 #(
		.INIT('h8000)
	) name1938 (
		_w1968_,
		_w1971_,
		_w1960_,
		_w1965_,
		_w1972_
	);
	LUT3 #(
		.INIT('h80)
	) name1939 (
		_w1959_,
		_w1955_,
		_w1972_,
		_w1973_
	);
	LUT4 #(
		.INIT('h153f)
	) name1940 (
		_w110_,
		_w65_,
		_w201_,
		_w236_,
		_w1974_
	);
	LUT4 #(
		.INIT('h135f)
	) name1941 (
		_w55_,
		_w47_,
		_w176_,
		_w430_,
		_w1975_
	);
	LUT4 #(
		.INIT('h153f)
	) name1942 (
		_w67_,
		_w78_,
		_w65_,
		_w201_,
		_w1976_
	);
	LUT3 #(
		.INIT('h80)
	) name1943 (
		_w1975_,
		_w1976_,
		_w1974_,
		_w1977_
	);
	LUT4 #(
		.INIT('h0777)
	) name1944 (
		_w110_,
		_w78_,
		_w44_,
		_w166_,
		_w1978_
	);
	LUT4 #(
		.INIT('h4000)
	) name1945 (
		_w390_,
		_w863_,
		_w1603_,
		_w1978_,
		_w1979_
	);
	LUT3 #(
		.INIT('h80)
	) name1946 (
		_w1932_,
		_w1977_,
		_w1979_,
		_w1980_
	);
	LUT3 #(
		.INIT('h80)
	) name1947 (
		_w861_,
		_w948_,
		_w1014_,
		_w1981_
	);
	LUT4 #(
		.INIT('h153f)
	) name1948 (
		_w59_,
		_w78_,
		_w56_,
		_w259_,
		_w1982_
	);
	LUT4 #(
		.INIT('h153f)
	) name1949 (
		_w38_,
		_w90_,
		_w158_,
		_w378_,
		_w1983_
	);
	LUT4 #(
		.INIT('h01ff)
	) name1950 (
		_w90_,
		_w56_,
		_w47_,
		_w378_,
		_w1984_
	);
	LUT3 #(
		.INIT('h80)
	) name1951 (
		_w1982_,
		_w1983_,
		_w1984_,
		_w1985_
	);
	LUT4 #(
		.INIT('h135f)
	) name1952 (
		_w106_,
		_w41_,
		_w44_,
		_w201_,
		_w1986_
	);
	LUT4 #(
		.INIT('h4000)
	) name1953 (
		_w190_,
		_w479_,
		_w1726_,
		_w1986_,
		_w1987_
	);
	LUT4 #(
		.INIT('h8000)
	) name1954 (
		_w1422_,
		_w1987_,
		_w1981_,
		_w1985_,
		_w1988_
	);
	LUT4 #(
		.INIT('h153f)
	) name1955 (
		_w110_,
		_w65_,
		_w166_,
		_w158_,
		_w1989_
	);
	LUT2 #(
		.INIT('h4)
	) name1956 (
		_w363_,
		_w1989_,
		_w1990_
	);
	LUT3 #(
		.INIT('h1f)
	) name1957 (
		_w85_,
		_w65_,
		_w378_,
		_w1991_
	);
	LUT4 #(
		.INIT('h0777)
	) name1958 (
		_w122_,
		_w55_,
		_w78_,
		_w50_,
		_w1992_
	);
	LUT4 #(
		.INIT('h153f)
	) name1959 (
		_w38_,
		_w59_,
		_w201_,
		_w259_,
		_w1993_
	);
	LUT4 #(
		.INIT('h8000)
	) name1960 (
		_w562_,
		_w1991_,
		_w1992_,
		_w1993_,
		_w1994_
	);
	LUT2 #(
		.INIT('h8)
	) name1961 (
		_w1990_,
		_w1994_,
		_w1995_
	);
	LUT4 #(
		.INIT('h8000)
	) name1962 (
		_w82_,
		_w92_,
		_w1990_,
		_w1994_,
		_w1996_
	);
	LUT4 #(
		.INIT('h8000)
	) name1963 (
		_w76_,
		_w1980_,
		_w1988_,
		_w1996_,
		_w1997_
	);
	LUT2 #(
		.INIT('h8)
	) name1964 (
		_w1973_,
		_w1997_,
		_w1998_
	);
	LUT4 #(
		.INIT('h0777)
	) name1965 (
		_w1501_,
		_w1949_,
		_w1973_,
		_w1997_,
		_w1999_
	);
	LUT4 #(
		.INIT('h153f)
	) name1966 (
		_w85_,
		_w90_,
		_w236_,
		_w176_,
		_w2000_
	);
	LUT4 #(
		.INIT('h8000)
	) name1967 (
		_w641_,
		_w974_,
		_w1643_,
		_w2000_,
		_w2001_
	);
	LUT2 #(
		.INIT('h4)
	) name1968 (
		_w167_,
		_w343_,
		_w2002_
	);
	LUT4 #(
		.INIT('h153f)
	) name1969 (
		_w110_,
		_w46_,
		_w166_,
		_w176_,
		_w2003_
	);
	LUT4 #(
		.INIT('h153f)
	) name1970 (
		_w41_,
		_w44_,
		_w259_,
		_w419_,
		_w2004_
	);
	LUT4 #(
		.INIT('h0777)
	) name1971 (
		_w38_,
		_w39_,
		_w50_,
		_w201_,
		_w2005_
	);
	LUT4 #(
		.INIT('h8000)
	) name1972 (
		_w311_,
		_w2005_,
		_w2003_,
		_w2004_,
		_w2006_
	);
	LUT3 #(
		.INIT('h80)
	) name1973 (
		_w2002_,
		_w2001_,
		_w2006_,
		_w2007_
	);
	LUT4 #(
		.INIT('h135f)
	) name1974 (
		_w85_,
		_w65_,
		_w236_,
		_w158_,
		_w2008_
	);
	LUT2 #(
		.INIT('h4)
	) name1975 (
		_w355_,
		_w2008_,
		_w2009_
	);
	LUT4 #(
		.INIT('h153f)
	) name1976 (
		_w52_,
		_w59_,
		_w201_,
		_w176_,
		_w2010_
	);
	LUT4 #(
		.INIT('h135f)
	) name1977 (
		_w122_,
		_w85_,
		_w56_,
		_w378_,
		_w2011_
	);
	LUT4 #(
		.INIT('h0777)
	) name1978 (
		_w106_,
		_w85_,
		_w90_,
		_w72_,
		_w2012_
	);
	LUT4 #(
		.INIT('h8000)
	) name1979 (
		_w687_,
		_w2012_,
		_w2010_,
		_w2011_,
		_w2013_
	);
	LUT2 #(
		.INIT('h8)
	) name1980 (
		_w2009_,
		_w2013_,
		_w2014_
	);
	LUT4 #(
		.INIT('h0777)
	) name1981 (
		_w110_,
		_w72_,
		_w65_,
		_w419_,
		_w2015_
	);
	LUT4 #(
		.INIT('h153f)
	) name1982 (
		_w38_,
		_w106_,
		_w56_,
		_w72_,
		_w2016_
	);
	LUT4 #(
		.INIT('h8000)
	) name1983 (
		_w1401_,
		_w1683_,
		_w2015_,
		_w2016_,
		_w2017_
	);
	LUT4 #(
		.INIT('h8000)
	) name1984 (
		_w580_,
		_w611_,
		_w1174_,
		_w1265_,
		_w2018_
	);
	LUT4 #(
		.INIT('h0777)
	) name1985 (
		_w67_,
		_w72_,
		_w44_,
		_w236_,
		_w2019_
	);
	LUT4 #(
		.INIT('h153f)
	) name1986 (
		_w55_,
		_w47_,
		_w158_,
		_w176_,
		_w2020_
	);
	LUT4 #(
		.INIT('h4000)
	) name1987 (
		_w275_,
		_w706_,
		_w2019_,
		_w2020_,
		_w2021_
	);
	LUT3 #(
		.INIT('h80)
	) name1988 (
		_w2017_,
		_w2018_,
		_w2021_,
		_w2022_
	);
	LUT3 #(
		.INIT('h80)
	) name1989 (
		_w2014_,
		_w2007_,
		_w2022_,
		_w2023_
	);
	LUT4 #(
		.INIT('h135f)
	) name1990 (
		_w85_,
		_w93_,
		_w184_,
		_w419_,
		_w2024_
	);
	LUT4 #(
		.INIT('h0800)
	) name1991 (
		_w115_,
		_w211_,
		_w476_,
		_w2024_,
		_w2025_
	);
	LUT4 #(
		.INIT('h1000)
	) name1992 (
		_w473_,
		_w469_,
		_w1356_,
		_w1587_,
		_w2026_
	);
	LUT4 #(
		.INIT('h135f)
	) name1993 (
		_w55_,
		_w110_,
		_w43_,
		_w158_,
		_w2027_
	);
	LUT3 #(
		.INIT('h40)
	) name1994 (
		_w124_,
		_w621_,
		_w2027_,
		_w2028_
	);
	LUT3 #(
		.INIT('h80)
	) name1995 (
		_w2026_,
		_w2028_,
		_w2025_,
		_w2029_
	);
	LUT4 #(
		.INIT('h153f)
	) name1996 (
		_w55_,
		_w59_,
		_w236_,
		_w158_,
		_w2030_
	);
	LUT4 #(
		.INIT('h135f)
	) name1997 (
		_w110_,
		_w41_,
		_w43_,
		_w158_,
		_w2031_
	);
	LUT4 #(
		.INIT('h4000)
	) name1998 (
		_w263_,
		_w750_,
		_w2031_,
		_w2030_,
		_w2032_
	);
	LUT4 #(
		.INIT('h1000)
	) name1999 (
		_w339_,
		_w383_,
		_w1141_,
		_w1945_,
		_w2033_
	);
	LUT3 #(
		.INIT('h80)
	) name2000 (
		_w817_,
		_w863_,
		_w1269_,
		_w2034_
	);
	LUT4 #(
		.INIT('h8000)
	) name2001 (
		_w1579_,
		_w2034_,
		_w2032_,
		_w2033_,
		_w2035_
	);
	LUT2 #(
		.INIT('h8)
	) name2002 (
		_w2029_,
		_w2035_,
		_w2036_
	);
	LUT4 #(
		.INIT('h135f)
	) name2003 (
		_w38_,
		_w93_,
		_w259_,
		_w378_,
		_w2037_
	);
	LUT2 #(
		.INIT('h4)
	) name2004 (
		_w478_,
		_w2037_,
		_w2038_
	);
	LUT4 #(
		.INIT('h153f)
	) name2005 (
		_w38_,
		_w122_,
		_w90_,
		_w419_,
		_w2039_
	);
	LUT4 #(
		.INIT('h135f)
	) name2006 (
		_w78_,
		_w47_,
		_w41_,
		_w184_,
		_w2040_
	);
	LUT4 #(
		.INIT('h153f)
	) name2007 (
		_w59_,
		_w67_,
		_w201_,
		_w158_,
		_w2041_
	);
	LUT3 #(
		.INIT('h80)
	) name2008 (
		_w2039_,
		_w2040_,
		_w2041_,
		_w2042_
	);
	LUT2 #(
		.INIT('h8)
	) name2009 (
		_w2038_,
		_w2042_,
		_w2043_
	);
	LUT4 #(
		.INIT('h0777)
	) name2010 (
		_w38_,
		_w106_,
		_w78_,
		_w56_,
		_w2044_
	);
	LUT2 #(
		.INIT('h4)
	) name2011 (
		_w241_,
		_w2044_,
		_w2045_
	);
	LUT4 #(
		.INIT('h0777)
	) name2012 (
		_w56_,
		_w43_,
		_w46_,
		_w259_,
		_w2046_
	);
	LUT4 #(
		.INIT('h0777)
	) name2013 (
		_w39_,
		_w50_,
		_w93_,
		_w201_,
		_w2047_
	);
	LUT4 #(
		.INIT('h153f)
	) name2014 (
		_w52_,
		_w56_,
		_w236_,
		_w378_,
		_w2048_
	);
	LUT4 #(
		.INIT('h4000)
	) name2015 (
		_w346_,
		_w2046_,
		_w2047_,
		_w2048_,
		_w2049_
	);
	LUT4 #(
		.INIT('h135f)
	) name2016 (
		_w106_,
		_w90_,
		_w93_,
		_w158_,
		_w2050_
	);
	LUT4 #(
		.INIT('h153f)
	) name2017 (
		_w38_,
		_w67_,
		_w43_,
		_w166_,
		_w2051_
	);
	LUT4 #(
		.INIT('h4000)
	) name2018 (
		_w455_,
		_w807_,
		_w2051_,
		_w2050_,
		_w2052_
	);
	LUT4 #(
		.INIT('h8000)
	) name2019 (
		_w562_,
		_w975_,
		_w1082_,
		_w1190_,
		_w2053_
	);
	LUT4 #(
		.INIT('h8000)
	) name2020 (
		_w2045_,
		_w2052_,
		_w2053_,
		_w2049_,
		_w2054_
	);
	LUT4 #(
		.INIT('h8000)
	) name2021 (
		_w2029_,
		_w2035_,
		_w2043_,
		_w2054_,
		_w2055_
	);
	LUT2 #(
		.INIT('h8)
	) name2022 (
		_w2023_,
		_w2055_,
		_w2056_
	);
	LUT4 #(
		.INIT('h153f)
	) name2023 (
		_w122_,
		_w59_,
		_w78_,
		_w65_,
		_w2057_
	);
	LUT4 #(
		.INIT('h153f)
	) name2024 (
		_w85_,
		_w50_,
		_w158_,
		_w176_,
		_w2058_
	);
	LUT2 #(
		.INIT('h8)
	) name2025 (
		_w2057_,
		_w2058_,
		_w2059_
	);
	LUT4 #(
		.INIT('h153f)
	) name2026 (
		_w59_,
		_w72_,
		_w65_,
		_w201_,
		_w2060_
	);
	LUT3 #(
		.INIT('h80)
	) name2027 (
		_w1435_,
		_w1598_,
		_w2060_,
		_w2061_
	);
	LUT2 #(
		.INIT('h8)
	) name2028 (
		_w2059_,
		_w2061_,
		_w2062_
	);
	LUT4 #(
		.INIT('h135f)
	) name2029 (
		_w67_,
		_w44_,
		_w176_,
		_w378_,
		_w2063_
	);
	LUT4 #(
		.INIT('h1000)
	) name2030 (
		_w185_,
		_w458_,
		_w690_,
		_w2063_,
		_w2064_
	);
	LUT2 #(
		.INIT('h4)
	) name2031 (
		_w261_,
		_w760_,
		_w2065_
	);
	LUT4 #(
		.INIT('h1000)
	) name2032 (
		_w261_,
		_w473_,
		_w760_,
		_w1356_,
		_w2066_
	);
	LUT4 #(
		.INIT('h135f)
	) name2033 (
		_w55_,
		_w41_,
		_w43_,
		_w419_,
		_w2067_
	);
	LUT4 #(
		.INIT('h0777)
	) name2034 (
		_w55_,
		_w78_,
		_w43_,
		_w93_,
		_w2068_
	);
	LUT4 #(
		.INIT('h135f)
	) name2035 (
		_w38_,
		_w110_,
		_w201_,
		_w176_,
		_w2069_
	);
	LUT3 #(
		.INIT('h80)
	) name2036 (
		_w2067_,
		_w2068_,
		_w2069_,
		_w2070_
	);
	LUT4 #(
		.INIT('h135f)
	) name2037 (
		_w106_,
		_w52_,
		_w110_,
		_w236_,
		_w2071_
	);
	LUT4 #(
		.INIT('h153f)
	) name2038 (
		_w122_,
		_w56_,
		_w72_,
		_w50_,
		_w2072_
	);
	LUT3 #(
		.INIT('h1f)
	) name2039 (
		_w85_,
		_w46_,
		_w201_,
		_w2073_
	);
	LUT4 #(
		.INIT('h8000)
	) name2040 (
		_w1416_,
		_w2072_,
		_w2073_,
		_w2071_,
		_w2074_
	);
	LUT4 #(
		.INIT('h8000)
	) name2041 (
		_w2070_,
		_w2074_,
		_w2064_,
		_w2066_,
		_w2075_
	);
	LUT3 #(
		.INIT('h80)
	) name2042 (
		_w1591_,
		_w2062_,
		_w2075_,
		_w2076_
	);
	LUT4 #(
		.INIT('h135f)
	) name2043 (
		_w85_,
		_w110_,
		_w184_,
		_w201_,
		_w2077_
	);
	LUT4 #(
		.INIT('h153f)
	) name2044 (
		_w110_,
		_w90_,
		_w419_,
		_w430_,
		_w2078_
	);
	LUT2 #(
		.INIT('h8)
	) name2045 (
		_w2077_,
		_w2078_,
		_w2079_
	);
	LUT4 #(
		.INIT('h153f)
	) name2046 (
		_w47_,
		_w39_,
		_w50_,
		_w43_,
		_w2080_
	);
	LUT4 #(
		.INIT('h8000)
	) name2047 (
		_w150_,
		_w513_,
		_w1303_,
		_w2080_,
		_w2081_
	);
	LUT4 #(
		.INIT('h135f)
	) name2048 (
		_w122_,
		_w52_,
		_w110_,
		_w43_,
		_w2082_
	);
	LUT4 #(
		.INIT('h135f)
	) name2049 (
		_w55_,
		_w41_,
		_w201_,
		_w158_,
		_w2083_
	);
	LUT4 #(
		.INIT('h8000)
	) name2050 (
		_w1514_,
		_w1783_,
		_w2082_,
		_w2083_,
		_w2084_
	);
	LUT4 #(
		.INIT('h8000)
	) name2051 (
		_w934_,
		_w2079_,
		_w2084_,
		_w2081_,
		_w2085_
	);
	LUT4 #(
		.INIT('h153f)
	) name2052 (
		_w52_,
		_w59_,
		_w43_,
		_w430_,
		_w2086_
	);
	LUT2 #(
		.INIT('h4)
	) name2053 (
		_w358_,
		_w2086_,
		_w2087_
	);
	LUT4 #(
		.INIT('h135f)
	) name2054 (
		_w67_,
		_w90_,
		_w43_,
		_w259_,
		_w2088_
	);
	LUT3 #(
		.INIT('h40)
	) name2055 (
		_w358_,
		_w2086_,
		_w2088_,
		_w2089_
	);
	LUT4 #(
		.INIT('h135f)
	) name2056 (
		_w85_,
		_w41_,
		_w72_,
		_w184_,
		_w2090_
	);
	LUT3 #(
		.INIT('h80)
	) name2057 (
		_w1037_,
		_w1683_,
		_w2090_,
		_w2091_
	);
	LUT3 #(
		.INIT('h37)
	) name2058 (
		_w90_,
		_w43_,
		_w46_,
		_w2092_
	);
	LUT4 #(
		.INIT('h135f)
	) name2059 (
		_w41_,
		_w39_,
		_w43_,
		_w44_,
		_w2093_
	);
	LUT4 #(
		.INIT('h8000)
	) name2060 (
		_w265_,
		_w713_,
		_w2092_,
		_w2093_,
		_w2094_
	);
	LUT3 #(
		.INIT('h80)
	) name2061 (
		_w2089_,
		_w2091_,
		_w2094_,
		_w2095_
	);
	LUT4 #(
		.INIT('h153f)
	) name2062 (
		_w55_,
		_w59_,
		_w166_,
		_w176_,
		_w2096_
	);
	LUT3 #(
		.INIT('h20)
	) name2063 (
		_w149_,
		_w392_,
		_w2096_,
		_w2097_
	);
	LUT4 #(
		.INIT('h8000)
	) name2064 (
		_w915_,
		_w1906_,
		_w1909_,
		_w2097_,
		_w2098_
	);
	LUT3 #(
		.INIT('h80)
	) name2065 (
		_w2085_,
		_w2095_,
		_w2098_,
		_w2099_
	);
	LUT3 #(
		.INIT('h80)
	) name2066 (
		_w1874_,
		_w2076_,
		_w2099_,
		_w2100_
	);
	LUT2 #(
		.INIT('h1)
	) name2067 (
		_w2056_,
		_w2100_,
		_w2101_
	);
	LUT4 #(
		.INIT('h153f)
	) name2068 (
		_w106_,
		_w47_,
		_w39_,
		_w65_,
		_w2102_
	);
	LUT4 #(
		.INIT('h8000)
	) name2069 (
		_w1198_,
		_w1826_,
		_w1837_,
		_w2102_,
		_w2103_
	);
	LUT4 #(
		.INIT('h153f)
	) name2070 (
		_w85_,
		_w65_,
		_w201_,
		_w430_,
		_w2104_
	);
	LUT4 #(
		.INIT('h8000)
	) name2071 (
		_w495_,
		_w960_,
		_w948_,
		_w2104_,
		_w2105_
	);
	LUT4 #(
		.INIT('h135f)
	) name2072 (
		_w90_,
		_w56_,
		_w166_,
		_w158_,
		_w2106_
	);
	LUT4 #(
		.INIT('h153f)
	) name2073 (
		_w38_,
		_w85_,
		_w158_,
		_w176_,
		_w2107_
	);
	LUT2 #(
		.INIT('h8)
	) name2074 (
		_w2106_,
		_w2107_,
		_w2108_
	);
	LUT4 #(
		.INIT('h8000)
	) name2075 (
		_w1079_,
		_w1190_,
		_w2106_,
		_w2107_,
		_w2109_
	);
	LUT3 #(
		.INIT('h80)
	) name2076 (
		_w2103_,
		_w2105_,
		_w2109_,
		_w2110_
	);
	LUT4 #(
		.INIT('h0777)
	) name2077 (
		_w52_,
		_w78_,
		_w50_,
		_w201_,
		_w2111_
	);
	LUT4 #(
		.INIT('h153f)
	) name2078 (
		_w52_,
		_w67_,
		_w43_,
		_w184_,
		_w2112_
	);
	LUT4 #(
		.INIT('h2000)
	) name2079 (
		_w58_,
		_w301_,
		_w2112_,
		_w2111_,
		_w2113_
	);
	LUT3 #(
		.INIT('h20)
	) name2080 (
		_w394_,
		_w436_,
		_w971_,
		_w2114_
	);
	LUT3 #(
		.INIT('h80)
	) name2081 (
		_w606_,
		_w2114_,
		_w2113_,
		_w2115_
	);
	LUT4 #(
		.INIT('h135f)
	) name2082 (
		_w90_,
		_w46_,
		_w236_,
		_w176_,
		_w2116_
	);
	LUT3 #(
		.INIT('h1f)
	) name2083 (
		_w93_,
		_w44_,
		_w259_,
		_w2117_
	);
	LUT4 #(
		.INIT('h153f)
	) name2084 (
		_w55_,
		_w39_,
		_w93_,
		_w184_,
		_w2118_
	);
	LUT4 #(
		.INIT('h8000)
	) name2085 (
		_w1956_,
		_w2116_,
		_w2117_,
		_w2118_,
		_w2119_
	);
	LUT4 #(
		.INIT('h0777)
	) name2086 (
		_w122_,
		_w56_,
		_w41_,
		_w259_,
		_w2120_
	);
	LUT4 #(
		.INIT('h153f)
	) name2087 (
		_w41_,
		_w72_,
		_w46_,
		_w201_,
		_w2121_
	);
	LUT4 #(
		.INIT('h2000)
	) name2088 (
		_w81_,
		_w366_,
		_w2121_,
		_w2120_,
		_w2122_
	);
	LUT4 #(
		.INIT('h8000)
	) name2089 (
		_w943_,
		_w947_,
		_w2119_,
		_w2122_,
		_w2123_
	);
	LUT3 #(
		.INIT('h80)
	) name2090 (
		_w2110_,
		_w2115_,
		_w2123_,
		_w2124_
	);
	LUT3 #(
		.INIT('h57)
	) name2091 (
		_w90_,
		_w43_,
		_w184_,
		_w2125_
	);
	LUT4 #(
		.INIT('h153f)
	) name2092 (
		_w85_,
		_w67_,
		_w78_,
		_w43_,
		_w2126_
	);
	LUT3 #(
		.INIT('h80)
	) name2093 (
		_w1967_,
		_w2126_,
		_w2125_,
		_w2127_
	);
	LUT4 #(
		.INIT('h8000)
	) name2094 (
		_w311_,
		_w361_,
		_w893_,
		_w856_,
		_w2128_
	);
	LUT4 #(
		.INIT('h0777)
	) name2095 (
		_w122_,
		_w47_,
		_w72_,
		_w44_,
		_w2129_
	);
	LUT4 #(
		.INIT('h0777)
	) name2096 (
		_w106_,
		_w67_,
		_w39_,
		_w46_,
		_w2130_
	);
	LUT4 #(
		.INIT('h8000)
	) name2097 (
		_w501_,
		_w502_,
		_w2129_,
		_w2130_,
		_w2131_
	);
	LUT4 #(
		.INIT('h8000)
	) name2098 (
		_w1197_,
		_w2127_,
		_w2128_,
		_w2131_,
		_w2132_
	);
	LUT3 #(
		.INIT('h80)
	) name2099 (
		_w2062_,
		_w2075_,
		_w2132_,
		_w2133_
	);
	LUT2 #(
		.INIT('h8)
	) name2100 (
		_w2124_,
		_w2133_,
		_w2134_
	);
	LUT4 #(
		.INIT('h153f)
	) name2101 (
		_w85_,
		_w52_,
		_w236_,
		_w259_,
		_w2135_
	);
	LUT4 #(
		.INIT('h153f)
	) name2102 (
		_w55_,
		_w93_,
		_w166_,
		_w176_,
		_w2136_
	);
	LUT4 #(
		.INIT('h153f)
	) name2103 (
		_w47_,
		_w50_,
		_w201_,
		_w236_,
		_w2137_
	);
	LUT3 #(
		.INIT('h80)
	) name2104 (
		_w2136_,
		_w2137_,
		_w2135_,
		_w2138_
	);
	LUT4 #(
		.INIT('h153f)
	) name2105 (
		_w90_,
		_w41_,
		_w39_,
		_w176_,
		_w2139_
	);
	LUT4 #(
		.INIT('h135f)
	) name2106 (
		_w55_,
		_w56_,
		_w158_,
		_w378_,
		_w2140_
	);
	LUT4 #(
		.INIT('h2000)
	) name2107 (
		_w260_,
		_w410_,
		_w2140_,
		_w2139_,
		_w2141_
	);
	LUT3 #(
		.INIT('h80)
	) name2108 (
		_w2065_,
		_w2138_,
		_w2141_,
		_w2142_
	);
	LUT4 #(
		.INIT('h153f)
	) name2109 (
		_w50_,
		_w46_,
		_w184_,
		_w176_,
		_w2143_
	);
	LUT2 #(
		.INIT('h8)
	) name2110 (
		_w172_,
		_w2143_,
		_w2144_
	);
	LUT3 #(
		.INIT('h37)
	) name2111 (
		_w56_,
		_w43_,
		_w65_,
		_w2145_
	);
	LUT3 #(
		.INIT('h37)
	) name2112 (
		_w122_,
		_w55_,
		_w72_,
		_w2146_
	);
	LUT4 #(
		.INIT('h4000)
	) name2113 (
		_w282_,
		_w381_,
		_w2146_,
		_w2145_,
		_w2147_
	);
	LUT2 #(
		.INIT('h8)
	) name2114 (
		_w2144_,
		_w2147_,
		_w2148_
	);
	LUT4 #(
		.INIT('h153f)
	) name2115 (
		_w67_,
		_w93_,
		_w236_,
		_w259_,
		_w2149_
	);
	LUT3 #(
		.INIT('h80)
	) name2116 (
		_w1560_,
		_w1783_,
		_w2149_,
		_w2150_
	);
	LUT3 #(
		.INIT('h57)
	) name2117 (
		_w56_,
		_w184_,
		_w430_,
		_w2151_
	);
	LUT2 #(
		.INIT('h8)
	) name2118 (
		_w583_,
		_w2151_,
		_w2152_
	);
	LUT4 #(
		.INIT('h8000)
	) name2119 (
		_w902_,
		_w1080_,
		_w1248_,
		_w1506_,
		_w2153_
	);
	LUT3 #(
		.INIT('h80)
	) name2120 (
		_w2152_,
		_w2150_,
		_w2153_,
		_w2154_
	);
	LUT3 #(
		.INIT('h80)
	) name2121 (
		_w2148_,
		_w2142_,
		_w2154_,
		_w2155_
	);
	LUT4 #(
		.INIT('h8000)
	) name2122 (
		_w1146_,
		_w1160_,
		_w1376_,
		_w1380_,
		_w2156_
	);
	LUT2 #(
		.INIT('h8)
	) name2123 (
		_w2155_,
		_w2156_,
		_w2157_
	);
	LUT4 #(
		.INIT('h0777)
	) name2124 (
		_w2124_,
		_w2133_,
		_w2155_,
		_w2156_,
		_w2158_
	);
	LUT3 #(
		.INIT('h40)
	) name2125 (
		_w84_,
		_w660_,
		_w894_,
		_w2159_
	);
	LUT4 #(
		.INIT('h153f)
	) name2126 (
		_w90_,
		_w39_,
		_w44_,
		_w201_,
		_w2160_
	);
	LUT4 #(
		.INIT('h8000)
	) name2127 (
		_w580_,
		_w1281_,
		_w2000_,
		_w2160_,
		_w2161_
	);
	LUT4 #(
		.INIT('h0777)
	) name2128 (
		_w106_,
		_w59_,
		_w43_,
		_w65_,
		_w2162_
	);
	LUT4 #(
		.INIT('h153f)
	) name2129 (
		_w67_,
		_w90_,
		_w166_,
		_w419_,
		_w2163_
	);
	LUT4 #(
		.INIT('h4000)
	) name2130 (
		_w353_,
		_w1810_,
		_w2162_,
		_w2163_,
		_w2164_
	);
	LUT3 #(
		.INIT('h80)
	) name2131 (
		_w2159_,
		_w2161_,
		_w2164_,
		_w2165_
	);
	LUT3 #(
		.INIT('h37)
	) name2132 (
		_w67_,
		_w39_,
		_w50_,
		_w2166_
	);
	LUT4 #(
		.INIT('h153f)
	) name2133 (
		_w56_,
		_w46_,
		_w201_,
		_w166_,
		_w2167_
	);
	LUT2 #(
		.INIT('h8)
	) name2134 (
		_w2166_,
		_w2167_,
		_w2168_
	);
	LUT4 #(
		.INIT('h153f)
	) name2135 (
		_w56_,
		_w47_,
		_w236_,
		_w176_,
		_w2169_
	);
	LUT4 #(
		.INIT('h153f)
	) name2136 (
		_w110_,
		_w65_,
		_w236_,
		_w259_,
		_w2170_
	);
	LUT3 #(
		.INIT('h80)
	) name2137 (
		_w876_,
		_w2170_,
		_w2169_,
		_w2171_
	);
	LUT2 #(
		.INIT('h8)
	) name2138 (
		_w2168_,
		_w2171_,
		_w2172_
	);
	LUT4 #(
		.INIT('h0777)
	) name2139 (
		_w122_,
		_w110_,
		_w39_,
		_w46_,
		_w2173_
	);
	LUT2 #(
		.INIT('h4)
	) name2140 (
		_w237_,
		_w2173_,
		_w2174_
	);
	LUT4 #(
		.INIT('h1000)
	) name2141 (
		_w206_,
		_w444_,
		_w713_,
		_w1744_,
		_w2175_
	);
	LUT4 #(
		.INIT('h135f)
	) name2142 (
		_w78_,
		_w41_,
		_w46_,
		_w184_,
		_w2176_
	);
	LUT4 #(
		.INIT('h135f)
	) name2143 (
		_w55_,
		_w110_,
		_w201_,
		_w166_,
		_w2177_
	);
	LUT4 #(
		.INIT('h8000)
	) name2144 (
		_w292_,
		_w1628_,
		_w2176_,
		_w2177_,
		_w2178_
	);
	LUT4 #(
		.INIT('h0777)
	) name2145 (
		_w55_,
		_w78_,
		_w46_,
		_w430_,
		_w2179_
	);
	LUT3 #(
		.INIT('h37)
	) name2146 (
		_w38_,
		_w78_,
		_w90_,
		_w2180_
	);
	LUT4 #(
		.INIT('h2000)
	) name2147 (
		_w130_,
		_w432_,
		_w2180_,
		_w2179_,
		_w2181_
	);
	LUT4 #(
		.INIT('h8000)
	) name2148 (
		_w2174_,
		_w2178_,
		_w2181_,
		_w2175_,
		_w2182_
	);
	LUT3 #(
		.INIT('h80)
	) name2149 (
		_w2165_,
		_w2172_,
		_w2182_,
		_w2183_
	);
	LUT4 #(
		.INIT('h8000)
	) name2150 (
		_w512_,
		_w1137_,
		_w1703_,
		_w1668_,
		_w2184_
	);
	LUT4 #(
		.INIT('h153f)
	) name2151 (
		_w38_,
		_w43_,
		_w44_,
		_w158_,
		_w2185_
	);
	LUT4 #(
		.INIT('h1000)
	) name2152 (
		_w369_,
		_w450_,
		_w1165_,
		_w2185_,
		_w2186_
	);
	LUT2 #(
		.INIT('h4)
	) name2153 (
		_w243_,
		_w502_,
		_w2187_
	);
	LUT4 #(
		.INIT('h0777)
	) name2154 (
		_w90_,
		_w72_,
		_w44_,
		_w158_,
		_w2188_
	);
	LUT3 #(
		.INIT('h40)
	) name2155 (
		_w243_,
		_w502_,
		_w2188_,
		_w2189_
	);
	LUT3 #(
		.INIT('h57)
	) name2156 (
		_w106_,
		_w67_,
		_w46_,
		_w2190_
	);
	LUT3 #(
		.INIT('h80)
	) name2157 (
		_w1725_,
		_w2117_,
		_w2190_,
		_w2191_
	);
	LUT4 #(
		.INIT('h8000)
	) name2158 (
		_w2189_,
		_w2191_,
		_w2184_,
		_w2186_,
		_w2192_
	);
	LUT2 #(
		.INIT('h8)
	) name2159 (
		_w1536_,
		_w2192_,
		_w2193_
	);
	LUT4 #(
		.INIT('h135f)
	) name2160 (
		_w67_,
		_w90_,
		_w176_,
		_w419_,
		_w2194_
	);
	LUT3 #(
		.INIT('h40)
	) name2161 (
		_w295_,
		_w951_,
		_w2194_,
		_w2195_
	);
	LUT4 #(
		.INIT('h0777)
	) name2162 (
		_w78_,
		_w50_,
		_w65_,
		_w430_,
		_w2196_
	);
	LUT2 #(
		.INIT('h4)
	) name2163 (
		_w468_,
		_w2196_,
		_w2197_
	);
	LUT4 #(
		.INIT('h135f)
	) name2164 (
		_w52_,
		_w90_,
		_w236_,
		_w158_,
		_w2198_
	);
	LUT3 #(
		.INIT('h40)
	) name2165 (
		_w60_,
		_w2015_,
		_w2198_,
		_w2199_
	);
	LUT3 #(
		.INIT('h80)
	) name2166 (
		_w2197_,
		_w2195_,
		_w2199_,
		_w2200_
	);
	LUT2 #(
		.INIT('h4)
	) name2167 (
		_w477_,
		_w1139_,
		_w2201_
	);
	LUT3 #(
		.INIT('h80)
	) name2168 (
		_w1157_,
		_w1589_,
		_w1843_,
		_w2202_
	);
	LUT2 #(
		.INIT('h8)
	) name2169 (
		_w2201_,
		_w2202_,
		_w2203_
	);
	LUT4 #(
		.INIT('h8000)
	) name2170 (
		_w81_,
		_w384_,
		_w496_,
		_w1602_,
		_w2204_
	);
	LUT4 #(
		.INIT('h153f)
	) name2171 (
		_w52_,
		_w56_,
		_w236_,
		_w176_,
		_w2205_
	);
	LUT4 #(
		.INIT('h153f)
	) name2172 (
		_w85_,
		_w59_,
		_w72_,
		_w236_,
		_w2206_
	);
	LUT4 #(
		.INIT('h4000)
	) name2173 (
		_w451_,
		_w1561_,
		_w2205_,
		_w2206_,
		_w2207_
	);
	LUT3 #(
		.INIT('h40)
	) name2174 (
		_w215_,
		_w662_,
		_w834_,
		_w2208_
	);
	LUT3 #(
		.INIT('h1f)
	) name2175 (
		_w59_,
		_w41_,
		_w39_,
		_w2209_
	);
	LUT3 #(
		.INIT('h37)
	) name2176 (
		_w106_,
		_w93_,
		_w430_,
		_w2210_
	);
	LUT3 #(
		.INIT('h80)
	) name2177 (
		_w2016_,
		_w2210_,
		_w2209_,
		_w2211_
	);
	LUT4 #(
		.INIT('h8000)
	) name2178 (
		_w2208_,
		_w2211_,
		_w2204_,
		_w2207_,
		_w2212_
	);
	LUT3 #(
		.INIT('h80)
	) name2179 (
		_w2200_,
		_w2203_,
		_w2212_,
		_w2213_
	);
	LUT3 #(
		.INIT('h80)
	) name2180 (
		_w2193_,
		_w2183_,
		_w2213_,
		_w2214_
	);
	LUT3 #(
		.INIT('h20)
	) name2181 (
		_w87_,
		_w135_,
		_w992_,
		_w2215_
	);
	LUT2 #(
		.INIT('h8)
	) name2182 (
		_w1030_,
		_w2215_,
		_w2216_
	);
	LUT4 #(
		.INIT('h135f)
	) name2183 (
		_w52_,
		_w41_,
		_w72_,
		_w176_,
		_w2217_
	);
	LUT3 #(
		.INIT('h80)
	) name2184 (
		_w538_,
		_w752_,
		_w2217_,
		_w2218_
	);
	LUT4 #(
		.INIT('h135f)
	) name2185 (
		_w122_,
		_w52_,
		_w93_,
		_w259_,
		_w2219_
	);
	LUT4 #(
		.INIT('h8000)
	) name2186 (
		_w820_,
		_w1472_,
		_w1844_,
		_w2219_,
		_w2220_
	);
	LUT4 #(
		.INIT('h153f)
	) name2187 (
		_w67_,
		_w41_,
		_w39_,
		_w236_,
		_w2221_
	);
	LUT4 #(
		.INIT('h135f)
	) name2188 (
		_w38_,
		_w52_,
		_w184_,
		_w158_,
		_w2222_
	);
	LUT4 #(
		.INIT('h153f)
	) name2189 (
		_w90_,
		_w56_,
		_w39_,
		_w184_,
		_w2223_
	);
	LUT4 #(
		.INIT('h4000)
	) name2190 (
		_w469_,
		_w2222_,
		_w2223_,
		_w2221_,
		_w2224_
	);
	LUT4 #(
		.INIT('h153f)
	) name2191 (
		_w59_,
		_w78_,
		_w50_,
		_w158_,
		_w2225_
	);
	LUT3 #(
		.INIT('h80)
	) name2192 (
		_w908_,
		_w1082_,
		_w2225_,
		_w2226_
	);
	LUT4 #(
		.INIT('h8000)
	) name2193 (
		_w2224_,
		_w2226_,
		_w2218_,
		_w2220_,
		_w2227_
	);
	LUT2 #(
		.INIT('h8)
	) name2194 (
		_w2216_,
		_w2227_,
		_w2228_
	);
	LUT4 #(
		.INIT('h135f)
	) name2195 (
		_w38_,
		_w90_,
		_w378_,
		_w430_,
		_w2229_
	);
	LUT3 #(
		.INIT('h40)
	) name2196 (
		_w235_,
		_w1450_,
		_w2229_,
		_w2230_
	);
	LUT4 #(
		.INIT('h153f)
	) name2197 (
		_w110_,
		_w47_,
		_w201_,
		_w259_,
		_w2231_
	);
	LUT4 #(
		.INIT('h8000)
	) name2198 (
		_w1403_,
		_w1473_,
		_w2137_,
		_w2231_,
		_w2232_
	);
	LUT3 #(
		.INIT('h80)
	) name2199 (
		_w2089_,
		_w2230_,
		_w2232_,
		_w2233_
	);
	LUT3 #(
		.INIT('h1f)
	) name2200 (
		_w55_,
		_w67_,
		_w166_,
		_w2234_
	);
	LUT4 #(
		.INIT('h153f)
	) name2201 (
		_w52_,
		_w56_,
		_w43_,
		_w166_,
		_w2235_
	);
	LUT4 #(
		.INIT('h8000)
	) name2202 (
		_w553_,
		_w1359_,
		_w2234_,
		_w2235_,
		_w2236_
	);
	LUT4 #(
		.INIT('h0777)
	) name2203 (
		_w106_,
		_w85_,
		_w90_,
		_w378_,
		_w2237_
	);
	LUT4 #(
		.INIT('h153f)
	) name2204 (
		_w47_,
		_w46_,
		_w201_,
		_w158_,
		_w2238_
	);
	LUT4 #(
		.INIT('h153f)
	) name2205 (
		_w67_,
		_w65_,
		_w259_,
		_w378_,
		_w2239_
	);
	LUT4 #(
		.INIT('h8000)
	) name2206 (
		_w1158_,
		_w2237_,
		_w2238_,
		_w2239_,
		_w2240_
	);
	LUT3 #(
		.INIT('h57)
	) name2207 (
		_w52_,
		_w78_,
		_w419_,
		_w2241_
	);
	LUT4 #(
		.INIT('h8000)
	) name2208 (
		_w296_,
		_w281_,
		_w1012_,
		_w2241_,
		_w2242_
	);
	LUT2 #(
		.INIT('h4)
	) name2209 (
		_w224_,
		_w555_,
		_w2243_
	);
	LUT4 #(
		.INIT('h4000)
	) name2210 (
		_w224_,
		_w555_,
		_w834_,
		_w1047_,
		_w2244_
	);
	LUT4 #(
		.INIT('h8000)
	) name2211 (
		_w2236_,
		_w2240_,
		_w2242_,
		_w2244_,
		_w2245_
	);
	LUT4 #(
		.INIT('h153f)
	) name2212 (
		_w110_,
		_w39_,
		_w46_,
		_w430_,
		_w2246_
	);
	LUT4 #(
		.INIT('h8000)
	) name2213 (
		_w1628_,
		_w1852_,
		_w1895_,
		_w2246_,
		_w2247_
	);
	LUT4 #(
		.INIT('h0757)
	) name2214 (
		_w72_,
		_w50_,
		_w93_,
		_w430_,
		_w2248_
	);
	LUT3 #(
		.INIT('h80)
	) name2215 (
		_w1269_,
		_w1483_,
		_w2248_,
		_w2249_
	);
	LUT2 #(
		.INIT('h8)
	) name2216 (
		_w2247_,
		_w2249_,
		_w2250_
	);
	LUT4 #(
		.INIT('h8000)
	) name2217 (
		_w68_,
		_w252_,
		_w491_,
		_w668_,
		_w2251_
	);
	LUT4 #(
		.INIT('h153f)
	) name2218 (
		_w85_,
		_w78_,
		_w41_,
		_w39_,
		_w2252_
	);
	LUT4 #(
		.INIT('h0777)
	) name2219 (
		_w78_,
		_w47_,
		_w50_,
		_w184_,
		_w2253_
	);
	LUT4 #(
		.INIT('h153f)
	) name2220 (
		_w44_,
		_w46_,
		_w259_,
		_w378_,
		_w2254_
	);
	LUT4 #(
		.INIT('h8000)
	) name2221 (
		_w1910_,
		_w2252_,
		_w2253_,
		_w2254_,
		_w2255_
	);
	LUT4 #(
		.INIT('h135f)
	) name2222 (
		_w122_,
		_w72_,
		_w65_,
		_w46_,
		_w2256_
	);
	LUT4 #(
		.INIT('h135f)
	) name2223 (
		_w38_,
		_w47_,
		_w72_,
		_w176_,
		_w2257_
	);
	LUT3 #(
		.INIT('h57)
	) name2224 (
		_w67_,
		_w72_,
		_w430_,
		_w2258_
	);
	LUT3 #(
		.INIT('h80)
	) name2225 (
		_w2257_,
		_w2258_,
		_w2256_,
		_w2259_
	);
	LUT4 #(
		.INIT('h8000)
	) name2226 (
		_w1173_,
		_w1687_,
		_w1725_,
		_w1982_,
		_w2260_
	);
	LUT4 #(
		.INIT('h8000)
	) name2227 (
		_w2259_,
		_w2260_,
		_w2251_,
		_w2255_,
		_w2261_
	);
	LUT4 #(
		.INIT('h8000)
	) name2228 (
		_w2250_,
		_w2233_,
		_w2245_,
		_w2261_,
		_w2262_
	);
	LUT2 #(
		.INIT('h8)
	) name2229 (
		_w2228_,
		_w2262_,
		_w2263_
	);
	LUT4 #(
		.INIT('h8000)
	) name2230 (
		_w191_,
		_w513_,
		_w649_,
		_w905_,
		_w2264_
	);
	LUT3 #(
		.INIT('h57)
	) name2231 (
		_w59_,
		_w72_,
		_w184_,
		_w2265_
	);
	LUT4 #(
		.INIT('h4000)
	) name2232 (
		_w237_,
		_w1504_,
		_w1505_,
		_w2265_,
		_w2266_
	);
	LUT4 #(
		.INIT('h135f)
	) name2233 (
		_w106_,
		_w55_,
		_w41_,
		_w158_,
		_w2267_
	);
	LUT4 #(
		.INIT('h0800)
	) name2234 (
		_w292_,
		_w384_,
		_w437_,
		_w2267_,
		_w2268_
	);
	LUT3 #(
		.INIT('h80)
	) name2235 (
		_w2264_,
		_w2266_,
		_w2268_,
		_w2269_
	);
	LUT4 #(
		.INIT('h115f)
	) name2236 (
		_w38_,
		_w110_,
		_w43_,
		_w176_,
		_w2270_
	);
	LUT4 #(
		.INIT('h2000)
	) name2237 (
		_w95_,
		_w347_,
		_w1308_,
		_w2270_,
		_w2271_
	);
	LUT3 #(
		.INIT('h80)
	) name2238 (
		_w2038_,
		_w2042_,
		_w2271_,
		_w2272_
	);
	LUT2 #(
		.INIT('h8)
	) name2239 (
		_w2269_,
		_w2272_,
		_w2273_
	);
	LUT4 #(
		.INIT('h135f)
	) name2240 (
		_w122_,
		_w39_,
		_w44_,
		_w46_,
		_w2274_
	);
	LUT4 #(
		.INIT('h135f)
	) name2241 (
		_w52_,
		_w50_,
		_w43_,
		_w158_,
		_w2275_
	);
	LUT4 #(
		.INIT('h8000)
	) name2242 (
		_w867_,
		_w1374_,
		_w2274_,
		_w2275_,
		_w2276_
	);
	LUT4 #(
		.INIT('h0777)
	) name2243 (
		_w38_,
		_w122_,
		_w106_,
		_w47_,
		_w2277_
	);
	LUT3 #(
		.INIT('h40)
	) name2244 (
		_w275_,
		_w1754_,
		_w2277_,
		_w2278_
	);
	LUT4 #(
		.INIT('h8000)
	) name2245 (
		_w188_,
		_w2026_,
		_w2278_,
		_w2276_,
		_w2279_
	);
	LUT4 #(
		.INIT('h135f)
	) name2246 (
		_w67_,
		_w41_,
		_w72_,
		_w166_,
		_w2280_
	);
	LUT4 #(
		.INIT('h0777)
	) name2247 (
		_w106_,
		_w85_,
		_w78_,
		_w56_,
		_w2281_
	);
	LUT4 #(
		.INIT('h153f)
	) name2248 (
		_w56_,
		_w39_,
		_w93_,
		_w166_,
		_w2282_
	);
	LUT4 #(
		.INIT('h8000)
	) name2249 (
		_w2116_,
		_w2280_,
		_w2281_,
		_w2282_,
		_w2283_
	);
	LUT4 #(
		.INIT('h153f)
	) name2250 (
		_w67_,
		_w65_,
		_w184_,
		_w236_,
		_w2284_
	);
	LUT4 #(
		.INIT('h0777)
	) name2251 (
		_w106_,
		_w90_,
		_w93_,
		_w176_,
		_w2285_
	);
	LUT4 #(
		.INIT('h8000)
	) name2252 (
		_w1643_,
		_w2083_,
		_w2284_,
		_w2285_,
		_w2286_
	);
	LUT2 #(
		.INIT('h8)
	) name2253 (
		_w2283_,
		_w2286_,
		_w2287_
	);
	LUT4 #(
		.INIT('h153f)
	) name2254 (
		_w78_,
		_w39_,
		_w65_,
		_w46_,
		_w2288_
	);
	LUT2 #(
		.INIT('h8)
	) name2255 (
		_w895_,
		_w2288_,
		_w2289_
	);
	LUT4 #(
		.INIT('h0777)
	) name2256 (
		_w47_,
		_w39_,
		_w93_,
		_w166_,
		_w2290_
	);
	LUT4 #(
		.INIT('h4000)
	) name2257 (
		_w398_,
		_w492_,
		_w611_,
		_w2290_,
		_w2291_
	);
	LUT4 #(
		.INIT('h8000)
	) name2258 (
		_w2289_,
		_w2283_,
		_w2286_,
		_w2291_,
		_w2292_
	);
	LUT4 #(
		.INIT('h8000)
	) name2259 (
		_w1536_,
		_w2192_,
		_w2279_,
		_w2292_,
		_w2293_
	);
	LUT2 #(
		.INIT('h8)
	) name2260 (
		_w2273_,
		_w2293_,
		_w2294_
	);
	LUT4 #(
		.INIT('heec8)
	) name2261 (
		_w2157_,
		_w2214_,
		_w2263_,
		_w2294_,
		_w2295_
	);
	LUT4 #(
		.INIT('h8000)
	) name2262 (
		_w2124_,
		_w2133_,
		_w2155_,
		_w2156_,
		_w2296_
	);
	LUT4 #(
		.INIT('h7888)
	) name2263 (
		_w2124_,
		_w2133_,
		_w2155_,
		_w2156_,
		_w2297_
	);
	LUT2 #(
		.INIT('h6)
	) name2264 (
		_w2100_,
		_w2134_,
		_w2298_
	);
	LUT4 #(
		.INIT('hecc8)
	) name2265 (
		_w2100_,
		_w2134_,
		_w2157_,
		_w2295_,
		_w2299_
	);
	LUT2 #(
		.INIT('h8)
	) name2266 (
		_w2056_,
		_w2100_,
		_w2300_
	);
	LUT2 #(
		.INIT('h6)
	) name2267 (
		_w2056_,
		_w2100_,
		_w2301_
	);
	LUT4 #(
		.INIT('h7888)
	) name2268 (
		_w1973_,
		_w1997_,
		_w2023_,
		_w2055_,
		_w2302_
	);
	LUT4 #(
		.INIT('hecc8)
	) name2269 (
		_w1998_,
		_w2056_,
		_w2100_,
		_w2299_,
		_w2303_
	);
	LUT4 #(
		.INIT('h8000)
	) name2270 (
		_w1501_,
		_w1949_,
		_w1973_,
		_w1997_,
		_w2304_
	);
	LUT4 #(
		.INIT('h7888)
	) name2271 (
		_w1501_,
		_w1949_,
		_w1973_,
		_w1997_,
		_w2305_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2272 (
		_w1501_,
		_w1898_,
		_w1928_,
		_w1949_,
		_w2306_
	);
	LUT4 #(
		.INIT('hecc8)
	) name2273 (
		_w1929_,
		_w1950_,
		_w1998_,
		_w2303_,
		_w2307_
	);
	LUT4 #(
		.INIT('h8000)
	) name2274 (
		_w1863_,
		_w1875_,
		_w1898_,
		_w1928_,
		_w2308_
	);
	LUT4 #(
		.INIT('h7888)
	) name2275 (
		_w1863_,
		_w1875_,
		_w1898_,
		_w1928_,
		_w2309_
	);
	LUT2 #(
		.INIT('h6)
	) name2276 (
		_w1841_,
		_w1876_,
		_w2310_
	);
	LUT4 #(
		.INIT('hecc8)
	) name2277 (
		_w1841_,
		_w1876_,
		_w1929_,
		_w2307_,
		_w2311_
	);
	LUT2 #(
		.INIT('h8)
	) name2278 (
		_w1797_,
		_w1841_,
		_w2312_
	);
	LUT2 #(
		.INIT('h6)
	) name2279 (
		_w1797_,
		_w1841_,
		_w2313_
	);
	LUT2 #(
		.INIT('h6)
	) name2280 (
		_w1772_,
		_w1797_,
		_w2314_
	);
	LUT4 #(
		.INIT('hecc8)
	) name2281 (
		_w1772_,
		_w1797_,
		_w1841_,
		_w2311_,
		_w2315_
	);
	LUT2 #(
		.INIT('h8)
	) name2282 (
		_w1724_,
		_w1772_,
		_w2316_
	);
	LUT2 #(
		.INIT('h6)
	) name2283 (
		_w1724_,
		_w1772_,
		_w2317_
	);
	LUT4 #(
		.INIT('h7888)
	) name2284 (
		_w1620_,
		_w1661_,
		_w1692_,
		_w1723_,
		_w2318_
	);
	LUT4 #(
		.INIT('hecc8)
	) name2285 (
		_w1662_,
		_w1724_,
		_w1772_,
		_w2315_,
		_w2319_
	);
	LUT2 #(
		.INIT('h8)
	) name2286 (
		_w1607_,
		_w1662_,
		_w2320_
	);
	LUT2 #(
		.INIT('h6)
	) name2287 (
		_w1607_,
		_w1662_,
		_w2321_
	);
	LUT2 #(
		.INIT('h6)
	) name2288 (
		_w1546_,
		_w1607_,
		_w2322_
	);
	LUT4 #(
		.INIT('hecc8)
	) name2289 (
		_w1546_,
		_w1607_,
		_w1662_,
		_w2319_,
		_w2323_
	);
	LUT2 #(
		.INIT('h8)
	) name2290 (
		_w1479_,
		_w1546_,
		_w2324_
	);
	LUT2 #(
		.INIT('h6)
	) name2291 (
		_w1479_,
		_w1546_,
		_w2325_
	);
	LUT2 #(
		.INIT('h6)
	) name2292 (
		_w1399_,
		_w1479_,
		_w2326_
	);
	LUT4 #(
		.INIT('hecc8)
	) name2293 (
		_w1399_,
		_w1479_,
		_w1546_,
		_w2323_,
		_w2327_
	);
	LUT4 #(
		.INIT('h8000)
	) name2294 (
		_w1325_,
		_w1367_,
		_w1381_,
		_w1398_,
		_w2328_
	);
	LUT4 #(
		.INIT('h7888)
	) name2295 (
		_w1325_,
		_w1367_,
		_w1381_,
		_w1398_,
		_w2329_
	);
	LUT4 #(
		.INIT('h7888)
	) name2296 (
		_w1253_,
		_w1294_,
		_w1325_,
		_w1367_,
		_w2330_
	);
	LUT4 #(
		.INIT('hecc8)
	) name2297 (
		_w1295_,
		_w1368_,
		_w1399_,
		_w2327_,
		_w2331_
	);
	LUT4 #(
		.INIT('h8000)
	) name2298 (
		_w1202_,
		_w1233_,
		_w1253_,
		_w1294_,
		_w2332_
	);
	LUT4 #(
		.INIT('h7888)
	) name2299 (
		_w1202_,
		_w1233_,
		_w1253_,
		_w1294_,
		_w2333_
	);
	LUT4 #(
		.INIT('h7888)
	) name2300 (
		_w1136_,
		_w1187_,
		_w1202_,
		_w1233_,
		_w2334_
	);
	LUT4 #(
		.INIT('hecc8)
	) name2301 (
		_w1188_,
		_w1234_,
		_w1295_,
		_w2331_,
		_w2335_
	);
	LUT4 #(
		.INIT('h8000)
	) name2302 (
		_w1071_,
		_w1102_,
		_w1136_,
		_w1187_,
		_w2336_
	);
	LUT4 #(
		.INIT('h7888)
	) name2303 (
		_w1071_,
		_w1102_,
		_w1136_,
		_w1187_,
		_w2337_
	);
	LUT4 #(
		.INIT('h7888)
	) name2304 (
		_w1009_,
		_w1050_,
		_w1071_,
		_w1102_,
		_w2338_
	);
	LUT4 #(
		.INIT('hecc8)
	) name2305 (
		_w1051_,
		_w1103_,
		_w1188_,
		_w2335_,
		_w2339_
	);
	LUT4 #(
		.INIT('h8000)
	) name2306 (
		_w763_,
		_w983_,
		_w1009_,
		_w1050_,
		_w2340_
	);
	LUT4 #(
		.INIT('h7888)
	) name2307 (
		_w763_,
		_w983_,
		_w1009_,
		_w1050_,
		_w2341_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name2308 (
		_w763_,
		_w871_,
		_w927_,
		_w983_,
		_w2342_
	);
	LUT4 #(
		.INIT('hecc8)
	) name2309 (
		_w928_,
		_w984_,
		_w1051_,
		_w2339_,
		_w2343_
	);
	LUT4 #(
		.INIT('h8000)
	) name2310 (
		_w801_,
		_w851_,
		_w871_,
		_w927_,
		_w2344_
	);
	LUT4 #(
		.INIT('h7888)
	) name2311 (
		_w801_,
		_w851_,
		_w871_,
		_w927_,
		_w2345_
	);
	LUT4 #(
		.INIT('h7888)
	) name2312 (
		_w725_,
		_w764_,
		_w801_,
		_w851_,
		_w2346_
	);
	LUT4 #(
		.INIT('hecc8)
	) name2313 (
		_w765_,
		_w852_,
		_w928_,
		_w2343_,
		_w2347_
	);
	LUT4 #(
		.INIT('h8000)
	) name2314 (
		_w666_,
		_w694_,
		_w725_,
		_w764_,
		_w2348_
	);
	LUT4 #(
		.INIT('h7888)
	) name2315 (
		_w666_,
		_w694_,
		_w725_,
		_w764_,
		_w2349_
	);
	LUT2 #(
		.INIT('h6)
	) name2316 (
		_w625_,
		_w695_,
		_w2350_
	);
	LUT4 #(
		.INIT('hecc8)
	) name2317 (
		_w625_,
		_w695_,
		_w765_,
		_w2347_,
		_w2351_
	);
	LUT2 #(
		.INIT('h8)
	) name2318 (
		_w559_,
		_w625_,
		_w2352_
	);
	LUT2 #(
		.INIT('h6)
	) name2319 (
		_w559_,
		_w625_,
		_w2353_
	);
	LUT2 #(
		.INIT('h6)
	) name2320 (
		_w510_,
		_w559_,
		_w2354_
	);
	LUT4 #(
		.INIT('hecc8)
	) name2321 (
		_w510_,
		_w559_,
		_w625_,
		_w2351_,
		_w2355_
	);
	LUT2 #(
		.INIT('h8)
	) name2322 (
		_w423_,
		_w510_,
		_w2356_
	);
	LUT2 #(
		.INIT('h6)
	) name2323 (
		_w423_,
		_w510_,
		_w2357_
	);
	LUT4 #(
		.INIT('h2000)
	) name2324 (
		_w121_,
		_w352_,
		_w418_,
		_w422_,
		_w2358_
	);
	LUT2 #(
		.INIT('h2)
	) name2325 (
		_w374_,
		_w423_,
		_w2359_
	);
	LUT3 #(
		.INIT('h0d)
	) name2326 (
		_w374_,
		_w423_,
		_w2358_,
		_w2360_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2327 (
		_w423_,
		_w510_,
		_w2355_,
		_w2360_,
		_w2361_
	);
	LUT4 #(
		.INIT('h4454)
	) name2328 (
		_w374_,
		_w376_,
		_w377_,
		_w2361_,
		_w2362_
	);
	LUT2 #(
		.INIT('h6)
	) name2329 (
		_w333_,
		_w2362_,
		_w2363_
	);
	LUT3 #(
		.INIT('h37)
	) name2330 (
		_w78_,
		_w47_,
		_w184_,
		_w2364_
	);
	LUT4 #(
		.INIT('h135f)
	) name2331 (
		_w67_,
		_w65_,
		_w184_,
		_w236_,
		_w2365_
	);
	LUT3 #(
		.INIT('h80)
	) name2332 (
		_w2246_,
		_w2365_,
		_w2364_,
		_w2366_
	);
	LUT4 #(
		.INIT('h8000)
	) name2333 (
		_w856_,
		_w1401_,
		_w1519_,
		_w2137_,
		_w2367_
	);
	LUT3 #(
		.INIT('h80)
	) name2334 (
		_w1702_,
		_w2366_,
		_w2367_,
		_w2368_
	);
	LUT4 #(
		.INIT('h135f)
	) name2335 (
		_w59_,
		_w44_,
		_w184_,
		_w259_,
		_w2369_
	);
	LUT4 #(
		.INIT('h153f)
	) name2336 (
		_w110_,
		_w65_,
		_w184_,
		_w176_,
		_w2370_
	);
	LUT4 #(
		.INIT('h8000)
	) name2337 (
		_w216_,
		_w1541_,
		_w2369_,
		_w2370_,
		_w2371_
	);
	LUT3 #(
		.INIT('h1f)
	) name2338 (
		_w122_,
		_w106_,
		_w47_,
		_w2372_
	);
	LUT4 #(
		.INIT('h135f)
	) name2339 (
		_w110_,
		_w72_,
		_w39_,
		_w46_,
		_w2373_
	);
	LUT4 #(
		.INIT('h0777)
	) name2340 (
		_w72_,
		_w93_,
		_w44_,
		_w184_,
		_w2374_
	);
	LUT4 #(
		.INIT('h4000)
	) name2341 (
		_w452_,
		_w2372_,
		_w2373_,
		_w2374_,
		_w2375_
	);
	LUT2 #(
		.INIT('h8)
	) name2342 (
		_w2371_,
		_w2375_,
		_w2376_
	);
	LUT4 #(
		.INIT('h0777)
	) name2343 (
		_w56_,
		_w39_,
		_w44_,
		_w378_,
		_w2377_
	);
	LUT4 #(
		.INIT('h8000)
	) name2344 (
		_w305_,
		_w1318_,
		_w1319_,
		_w2377_,
		_w2378_
	);
	LUT3 #(
		.INIT('h57)
	) name2345 (
		_w52_,
		_w158_,
		_w176_,
		_w2379_
	);
	LUT4 #(
		.INIT('h4000)
	) name2346 (
		_w243_,
		_w283_,
		_w502_,
		_w2379_,
		_w2380_
	);
	LUT4 #(
		.INIT('h8000)
	) name2347 (
		_w1123_,
		_w1128_,
		_w2378_,
		_w2380_,
		_w2381_
	);
	LUT3 #(
		.INIT('h80)
	) name2348 (
		_w2376_,
		_w2368_,
		_w2381_,
		_w2382_
	);
	LUT3 #(
		.INIT('h80)
	) name2349 (
		_w828_,
		_w1075_,
		_w1904_,
		_w2383_
	);
	LUT4 #(
		.INIT('h135f)
	) name2350 (
		_w106_,
		_w55_,
		_w65_,
		_w184_,
		_w2384_
	);
	LUT3 #(
		.INIT('h57)
	) name2351 (
		_w55_,
		_w176_,
		_w378_,
		_w2385_
	);
	LUT4 #(
		.INIT('h8000)
	) name2352 (
		_w553_,
		_w574_,
		_w2384_,
		_w2385_,
		_w2386_
	);
	LUT3 #(
		.INIT('h80)
	) name2353 (
		_w131_,
		_w2383_,
		_w2386_,
		_w2387_
	);
	LUT2 #(
		.INIT('h4)
	) name2354 (
		_w73_,
		_w743_,
		_w2388_
	);
	LUT4 #(
		.INIT('h8000)
	) name2355 (
		_w131_,
		_w2383_,
		_w2386_,
		_w2388_,
		_w2389_
	);
	LUT3 #(
		.INIT('h80)
	) name2356 (
		_w1376_,
		_w1380_,
		_w2389_,
		_w2390_
	);
	LUT2 #(
		.INIT('h8)
	) name2357 (
		_w2382_,
		_w2390_,
		_w2391_
	);
	LUT4 #(
		.INIT('h153f)
	) name2358 (
		_w67_,
		_w43_,
		_w65_,
		_w259_,
		_w2392_
	);
	LUT3 #(
		.INIT('h40)
	) name2359 (
		_w268_,
		_w1198_,
		_w2392_,
		_w2393_
	);
	LUT4 #(
		.INIT('h8000)
	) name2360 (
		_w526_,
		_w537_,
		_w543_,
		_w2393_,
		_w2394_
	);
	LUT2 #(
		.INIT('h4)
	) name2361 (
		_w80_,
		_w348_,
		_w2395_
	);
	LUT4 #(
		.INIT('h153f)
	) name2362 (
		_w38_,
		_w39_,
		_w46_,
		_w259_,
		_w2396_
	);
	LUT4 #(
		.INIT('h0777)
	) name2363 (
		_w122_,
		_w90_,
		_w72_,
		_w46_,
		_w2397_
	);
	LUT4 #(
		.INIT('h8000)
	) name2364 (
		_w1481_,
		_w1704_,
		_w2397_,
		_w2396_,
		_w2398_
	);
	LUT4 #(
		.INIT('h8000)
	) name2365 (
		_w127_,
		_w133_,
		_w2395_,
		_w2398_,
		_w2399_
	);
	LUT3 #(
		.INIT('h80)
	) name2366 (
		_w200_,
		_w449_,
		_w2399_,
		_w2400_
	);
	LUT3 #(
		.INIT('h80)
	) name2367 (
		_w179_,
		_w2394_,
		_w2400_,
		_w2401_
	);
	LUT4 #(
		.INIT('h044c)
	) name2368 (
		\a[29] ,
		_w330_,
		_w2391_,
		_w2401_,
		_w2402_
	);
	LUT4 #(
		.INIT('h3220)
	) name2369 (
		\a[29] ,
		_w330_,
		_w2391_,
		_w2401_,
		_w2403_
	);
	LUT4 #(
		.INIT('h1700)
	) name2370 (
		_w423_,
		_w510_,
		_w2355_,
		_w2359_,
		_w2404_
	);
	LUT4 #(
		.INIT('hcc40)
	) name2371 (
		_w374_,
		_w377_,
		_w2361_,
		_w2404_,
		_w2405_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2372 (
		_w121_,
		_w376_,
		_w418_,
		_w422_,
		_w2406_
	);
	LUT3 #(
		.INIT('h18)
	) name2373 (
		\a[29] ,
		\a[30] ,
		\a[31] ,
		_w2407_
	);
	LUT3 #(
		.INIT('h70)
	) name2374 (
		_w352_,
		_w373_,
		_w2407_,
		_w2408_
	);
	LUT2 #(
		.INIT('h1)
	) name2375 (
		_w2406_,
		_w2408_,
		_w2409_
	);
	LUT4 #(
		.INIT('h4544)
	) name2376 (
		_w2402_,
		_w2403_,
		_w2405_,
		_w2409_,
		_w2410_
	);
	LUT2 #(
		.INIT('h2)
	) name2377 (
		_w2363_,
		_w2410_,
		_w2411_
	);
	LUT2 #(
		.INIT('h9)
	) name2378 (
		_w2363_,
		_w2410_,
		_w2412_
	);
	LUT4 #(
		.INIT('h135f)
	) name2379 (
		_w59_,
		_w50_,
		_w43_,
		_w430_,
		_w2413_
	);
	LUT4 #(
		.INIT('h4000)
	) name2380 (
		_w440_,
		_w1037_,
		_w1198_,
		_w2413_,
		_w2414_
	);
	LUT4 #(
		.INIT('h135f)
	) name2381 (
		_w39_,
		_w50_,
		_w44_,
		_w166_,
		_w2415_
	);
	LUT4 #(
		.INIT('h1000)
	) name2382 (
		_w358_,
		_w458_,
		_w1845_,
		_w2415_,
		_w2416_
	);
	LUT2 #(
		.INIT('h8)
	) name2383 (
		_w2414_,
		_w2416_,
		_w2417_
	);
	LUT4 #(
		.INIT('h153f)
	) name2384 (
		_w56_,
		_w46_,
		_w236_,
		_w419_,
		_w2418_
	);
	LUT4 #(
		.INIT('h8000)
	) name2385 (
		_w978_,
		_w1156_,
		_w2369_,
		_w2418_,
		_w2419_
	);
	LUT3 #(
		.INIT('h80)
	) name2386 (
		_w1893_,
		_w2025_,
		_w2419_,
		_w2420_
	);
	LUT3 #(
		.INIT('h80)
	) name2387 (
		_w1980_,
		_w2417_,
		_w2420_,
		_w2421_
	);
	LUT4 #(
		.INIT('h135f)
	) name2388 (
		_w52_,
		_w67_,
		_w72_,
		_w158_,
		_w2422_
	);
	LUT2 #(
		.INIT('h4)
	) name2389 (
		_w369_,
		_w2422_,
		_w2423_
	);
	LUT4 #(
		.INIT('h0777)
	) name2390 (
		_w85_,
		_w78_,
		_w90_,
		_w39_,
		_w2424_
	);
	LUT4 #(
		.INIT('h135f)
	) name2391 (
		_w85_,
		_w93_,
		_w259_,
		_w378_,
		_w2425_
	);
	LUT4 #(
		.INIT('h8000)
	) name2392 (
		_w1354_,
		_w1355_,
		_w2424_,
		_w2425_,
		_w2426_
	);
	LUT4 #(
		.INIT('h135f)
	) name2393 (
		_w38_,
		_w93_,
		_w184_,
		_w236_,
		_w2427_
	);
	LUT3 #(
		.INIT('h80)
	) name2394 (
		_w2027_,
		_w2146_,
		_w2427_,
		_w2428_
	);
	LUT4 #(
		.INIT('h8000)
	) name2395 (
		_w464_,
		_w857_,
		_w1278_,
		_w1474_,
		_w2429_
	);
	LUT4 #(
		.INIT('h8000)
	) name2396 (
		_w2423_,
		_w2428_,
		_w2429_,
		_w2426_,
		_w2430_
	);
	LUT3 #(
		.INIT('h37)
	) name2397 (
		_w59_,
		_w78_,
		_w41_,
		_w2431_
	);
	LUT4 #(
		.INIT('h0737)
	) name2398 (
		_w122_,
		_w59_,
		_w78_,
		_w41_,
		_w2432_
	);
	LUT4 #(
		.INIT('h0777)
	) name2399 (
		_w106_,
		_w55_,
		_w90_,
		_w43_,
		_w2433_
	);
	LUT4 #(
		.INIT('h0200)
	) name2400 (
		_w132_,
		_w261_,
		_w432_,
		_w2433_,
		_w2434_
	);
	LUT4 #(
		.INIT('h8000)
	) name2401 (
		_w790_,
		_w829_,
		_w1047_,
		_w1652_,
		_w2435_
	);
	LUT4 #(
		.INIT('h153f)
	) name2402 (
		_w52_,
		_w47_,
		_w158_,
		_w259_,
		_w2436_
	);
	LUT4 #(
		.INIT('h0777)
	) name2403 (
		_w38_,
		_w122_,
		_w78_,
		_w46_,
		_w2437_
	);
	LUT4 #(
		.INIT('h4000)
	) name2404 (
		_w386_,
		_w381_,
		_w2437_,
		_w2436_,
		_w2438_
	);
	LUT4 #(
		.INIT('h8000)
	) name2405 (
		_w2432_,
		_w2435_,
		_w2438_,
		_w2434_,
		_w2439_
	);
	LUT4 #(
		.INIT('h135f)
	) name2406 (
		_w52_,
		_w110_,
		_w43_,
		_w419_,
		_w2440_
	);
	LUT4 #(
		.INIT('h8000)
	) name2407 (
		_w1079_,
		_w1154_,
		_w1321_,
		_w2440_,
		_w2441_
	);
	LUT3 #(
		.INIT('h57)
	) name2408 (
		_w65_,
		_w158_,
		_w419_,
		_w2442_
	);
	LUT4 #(
		.INIT('h153f)
	) name2409 (
		_w110_,
		_w67_,
		_w184_,
		_w201_,
		_w2443_
	);
	LUT4 #(
		.INIT('h4000)
	) name2410 (
		_w392_,
		_w840_,
		_w2443_,
		_w2442_,
		_w2444_
	);
	LUT4 #(
		.INIT('h8000)
	) name2411 (
		_w915_,
		_w920_,
		_w2441_,
		_w2444_,
		_w2445_
	);
	LUT3 #(
		.INIT('h80)
	) name2412 (
		_w2430_,
		_w2439_,
		_w2445_,
		_w2446_
	);
	LUT2 #(
		.INIT('h8)
	) name2413 (
		_w2421_,
		_w2446_,
		_w2447_
	);
	LUT4 #(
		.INIT('h0888)
	) name2414 (
		_w2382_,
		_w2390_,
		_w2421_,
		_w2446_,
		_w2448_
	);
	LUT4 #(
		.INIT('h8777)
	) name2415 (
		_w2382_,
		_w2390_,
		_w2421_,
		_w2446_,
		_w2449_
	);
	LUT4 #(
		.INIT('h0777)
	) name2416 (
		_w122_,
		_w55_,
		_w41_,
		_w72_,
		_w2450_
	);
	LUT4 #(
		.INIT('h153f)
	) name2417 (
		_w52_,
		_w72_,
		_w44_,
		_w236_,
		_w2451_
	);
	LUT4 #(
		.INIT('h4000)
	) name2418 (
		_w218_,
		_w1681_,
		_w2451_,
		_w2450_,
		_w2452_
	);
	LUT4 #(
		.INIT('h135f)
	) name2419 (
		_w50_,
		_w65_,
		_w166_,
		_w419_,
		_w2453_
	);
	LUT4 #(
		.INIT('h0777)
	) name2420 (
		_w72_,
		_w50_,
		_w44_,
		_w259_,
		_w2454_
	);
	LUT4 #(
		.INIT('h1000)
	) name2421 (
		_w393_,
		_w462_,
		_w2453_,
		_w2454_,
		_w2455_
	);
	LUT2 #(
		.INIT('h8)
	) name2422 (
		_w2452_,
		_w2455_,
		_w2456_
	);
	LUT4 #(
		.INIT('h01ff)
	) name2423 (
		_w110_,
		_w56_,
		_w46_,
		_w419_,
		_w2457_
	);
	LUT4 #(
		.INIT('h0777)
	) name2424 (
		_w110_,
		_w78_,
		_w39_,
		_w50_,
		_w2458_
	);
	LUT4 #(
		.INIT('h4000)
	) name2425 (
		_w383_,
		_w978_,
		_w935_,
		_w2458_,
		_w2459_
	);
	LUT4 #(
		.INIT('h135f)
	) name2426 (
		_w110_,
		_w50_,
		_w158_,
		_w430_,
		_w2460_
	);
	LUT4 #(
		.INIT('h135f)
	) name2427 (
		_w67_,
		_w90_,
		_w201_,
		_w419_,
		_w2461_
	);
	LUT4 #(
		.INIT('h4000)
	) name2428 (
		_w261_,
		_w2433_,
		_w2460_,
		_w2461_,
		_w2462_
	);
	LUT4 #(
		.INIT('h8000)
	) name2429 (
		_w1472_,
		_w1753_,
		_w1798_,
		_w2229_,
		_w2463_
	);
	LUT4 #(
		.INIT('h8000)
	) name2430 (
		_w2457_,
		_w2462_,
		_w2463_,
		_w2459_,
		_w2464_
	);
	LUT4 #(
		.INIT('h0777)
	) name2431 (
		_w67_,
		_w43_,
		_w44_,
		_w166_,
		_w2465_
	);
	LUT4 #(
		.INIT('h135f)
	) name2432 (
		_w85_,
		_w93_,
		_w201_,
		_w176_,
		_w2466_
	);
	LUT4 #(
		.INIT('h8000)
	) name2433 (
		_w742_,
		_w1936_,
		_w2465_,
		_w2466_,
		_w2467_
	);
	LUT4 #(
		.INIT('h153f)
	) name2434 (
		_w55_,
		_w67_,
		_w184_,
		_w419_,
		_w2468_
	);
	LUT4 #(
		.INIT('h8000)
	) name2435 (
		_w937_,
		_w1783_,
		_w2116_,
		_w2468_,
		_w2469_
	);
	LUT4 #(
		.INIT('h8000)
	) name2436 (
		_w96_,
		_w171_,
		_w491_,
		_w687_,
		_w2470_
	);
	LUT3 #(
		.INIT('h80)
	) name2437 (
		_w2467_,
		_w2469_,
		_w2470_,
		_w2471_
	);
	LUT4 #(
		.INIT('h153f)
	) name2438 (
		_w38_,
		_w65_,
		_w184_,
		_w259_,
		_w2472_
	);
	LUT3 #(
		.INIT('h80)
	) name2439 (
		_w1635_,
		_w2225_,
		_w2472_,
		_w2473_
	);
	LUT4 #(
		.INIT('h0777)
	) name2440 (
		_w52_,
		_w78_,
		_w56_,
		_w236_,
		_w2474_
	);
	LUT4 #(
		.INIT('h135f)
	) name2441 (
		_w110_,
		_w41_,
		_w201_,
		_w259_,
		_w2475_
	);
	LUT4 #(
		.INIT('h8000)
	) name2442 (
		_w797_,
		_w1004_,
		_w2474_,
		_w2475_,
		_w2476_
	);
	LUT4 #(
		.INIT('h135f)
	) name2443 (
		_w41_,
		_w50_,
		_w176_,
		_w378_,
		_w2477_
	);
	LUT2 #(
		.INIT('h4)
	) name2444 (
		_w51_,
		_w2477_,
		_w2478_
	);
	LUT4 #(
		.INIT('h0777)
	) name2445 (
		_w85_,
		_w39_,
		_w50_,
		_w236_,
		_w2479_
	);
	LUT4 #(
		.INIT('h4000)
	) name2446 (
		_w412_,
		_w403_,
		_w663_,
		_w2479_,
		_w2480_
	);
	LUT4 #(
		.INIT('h8000)
	) name2447 (
		_w2473_,
		_w2476_,
		_w2478_,
		_w2480_,
		_w2481_
	);
	LUT4 #(
		.INIT('h8000)
	) name2448 (
		_w2456_,
		_w2464_,
		_w2471_,
		_w2481_,
		_w2482_
	);
	LUT2 #(
		.INIT('h8)
	) name2449 (
		_w1584_,
		_w2482_,
		_w2483_
	);
	LUT3 #(
		.INIT('h1f)
	) name2450 (
		_w38_,
		_w41_,
		_w201_,
		_w2484_
	);
	LUT4 #(
		.INIT('h135f)
	) name2451 (
		_w110_,
		_w67_,
		_w236_,
		_w176_,
		_w2485_
	);
	LUT2 #(
		.INIT('h8)
	) name2452 (
		_w2484_,
		_w2485_,
		_w2486_
	);
	LUT3 #(
		.INIT('h80)
	) name2453 (
		_w916_,
		_w1483_,
		_w1651_,
		_w2487_
	);
	LUT2 #(
		.INIT('h8)
	) name2454 (
		_w2486_,
		_w2487_,
		_w2488_
	);
	LUT3 #(
		.INIT('h37)
	) name2455 (
		_w72_,
		_w50_,
		_w184_,
		_w2489_
	);
	LUT2 #(
		.INIT('h4)
	) name2456 (
		_w392_,
		_w2489_,
		_w2490_
	);
	LUT4 #(
		.INIT('h153f)
	) name2457 (
		_w38_,
		_w56_,
		_w158_,
		_w259_,
		_w2491_
	);
	LUT4 #(
		.INIT('h1000)
	) name2458 (
		_w452_,
		_w439_,
		_w442_,
		_w2491_,
		_w2492_
	);
	LUT4 #(
		.INIT('h153f)
	) name2459 (
		_w55_,
		_w85_,
		_w72_,
		_w158_,
		_w2493_
	);
	LUT4 #(
		.INIT('h153f)
	) name2460 (
		_w41_,
		_w50_,
		_w259_,
		_w430_,
		_w2494_
	);
	LUT4 #(
		.INIT('h153f)
	) name2461 (
		_w67_,
		_w39_,
		_w93_,
		_w158_,
		_w2495_
	);
	LUT4 #(
		.INIT('h8000)
	) name2462 (
		_w1519_,
		_w2493_,
		_w2494_,
		_w2495_,
		_w2496_
	);
	LUT4 #(
		.INIT('h8000)
	) name2463 (
		_w738_,
		_w863_,
		_w957_,
		_w1092_,
		_w2497_
	);
	LUT4 #(
		.INIT('h8000)
	) name2464 (
		_w2490_,
		_w2496_,
		_w2497_,
		_w2492_,
		_w2498_
	);
	LUT2 #(
		.INIT('h8)
	) name2465 (
		_w2488_,
		_w2498_,
		_w2499_
	);
	LUT4 #(
		.INIT('h135f)
	) name2466 (
		_w85_,
		_w90_,
		_w184_,
		_w176_,
		_w2500_
	);
	LUT3 #(
		.INIT('h20)
	) name2467 (
		_w343_,
		_w369_,
		_w2500_,
		_w2501_
	);
	LUT4 #(
		.INIT('h135f)
	) name2468 (
		_w106_,
		_w67_,
		_w47_,
		_w201_,
		_w2502_
	);
	LUT3 #(
		.INIT('h37)
	) name2469 (
		_w122_,
		_w55_,
		_w78_,
		_w2503_
	);
	LUT2 #(
		.INIT('h8)
	) name2470 (
		_w2502_,
		_w2503_,
		_w2504_
	);
	LUT4 #(
		.INIT('h153f)
	) name2471 (
		_w38_,
		_w106_,
		_w110_,
		_w72_,
		_w2505_
	);
	LUT3 #(
		.INIT('h57)
	) name2472 (
		_w110_,
		_w78_,
		_w166_,
		_w2506_
	);
	LUT4 #(
		.INIT('h8000)
	) name2473 (
		_w697_,
		_w820_,
		_w2505_,
		_w2506_,
		_w2507_
	);
	LUT3 #(
		.INIT('h80)
	) name2474 (
		_w2504_,
		_w2501_,
		_w2507_,
		_w2508_
	);
	LUT4 #(
		.INIT('h8000)
	) name2475 (
		_w876_,
		_w966_,
		_w1131_,
		_w1427_,
		_w2509_
	);
	LUT4 #(
		.INIT('h153f)
	) name2476 (
		_w38_,
		_w72_,
		_w46_,
		_w158_,
		_w2510_
	);
	LUT2 #(
		.INIT('h8)
	) name2477 (
		_w1371_,
		_w2510_,
		_w2511_
	);
	LUT4 #(
		.INIT('h153f)
	) name2478 (
		_w50_,
		_w46_,
		_w166_,
		_w378_,
		_w2512_
	);
	LUT4 #(
		.INIT('h8000)
	) name2479 (
		_w760_,
		_w1371_,
		_w2510_,
		_w2512_,
		_w2513_
	);
	LUT4 #(
		.INIT('h135f)
	) name2480 (
		_w106_,
		_w85_,
		_w52_,
		_w43_,
		_w2514_
	);
	LUT3 #(
		.INIT('h40)
	) name2481 (
		_w94_,
		_w408_,
		_w2514_,
		_w2515_
	);
	LUT3 #(
		.INIT('h1f)
	) name2482 (
		_w47_,
		_w46_,
		_w176_,
		_w2516_
	);
	LUT4 #(
		.INIT('h0777)
	) name2483 (
		_w122_,
		_w85_,
		_w90_,
		_w43_,
		_w2517_
	);
	LUT3 #(
		.INIT('h80)
	) name2484 (
		_w1586_,
		_w2517_,
		_w2516_,
		_w2518_
	);
	LUT4 #(
		.INIT('h8000)
	) name2485 (
		_w2515_,
		_w2518_,
		_w2509_,
		_w2513_,
		_w2519_
	);
	LUT4 #(
		.INIT('h8000)
	) name2486 (
		_w2233_,
		_w2245_,
		_w2508_,
		_w2519_,
		_w2520_
	);
	LUT2 #(
		.INIT('h8)
	) name2487 (
		_w2499_,
		_w2520_,
		_w2521_
	);
	LUT4 #(
		.INIT('h0777)
	) name2488 (
		_w1584_,
		_w2482_,
		_w2499_,
		_w2520_,
		_w2522_
	);
	LUT4 #(
		.INIT('h8000)
	) name2489 (
		_w1584_,
		_w2482_,
		_w2499_,
		_w2520_,
		_w2523_
	);
	LUT4 #(
		.INIT('h044c)
	) name2490 (
		\a[26] ,
		_w2447_,
		_w2483_,
		_w2521_,
		_w2524_
	);
	LUT4 #(
		.INIT('h3220)
	) name2491 (
		\a[26] ,
		_w2447_,
		_w2483_,
		_w2521_,
		_w2525_
	);
	LUT4 #(
		.INIT('h54ab)
	) name2492 (
		_w626_,
		_w2351_,
		_w2352_,
		_w2354_,
		_w2526_
	);
	LUT3 #(
		.INIT('h06)
	) name2493 (
		\a[29] ,
		\a[30] ,
		\a[31] ,
		_w2527_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2494 (
		_w486_,
		_w487_,
		_w509_,
		_w2527_,
		_w2528_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name2495 (
		_w376_,
		_w587_,
		_w608_,
		_w624_,
		_w2529_
	);
	LUT3 #(
		.INIT('h70)
	) name2496 (
		_w544_,
		_w558_,
		_w2407_,
		_w2530_
	);
	LUT3 #(
		.INIT('h01)
	) name2497 (
		_w2528_,
		_w2529_,
		_w2530_,
		_w2531_
	);
	LUT4 #(
		.INIT('h2033)
	) name2498 (
		_w377_,
		_w2525_,
		_w2526_,
		_w2531_,
		_w2532_
	);
	LUT4 #(
		.INIT('h1115)
	) name2499 (
		_w2448_,
		_w2449_,
		_w2524_,
		_w2532_,
		_w2533_
	);
	LUT3 #(
		.INIT('h96)
	) name2500 (
		\a[29] ,
		_w2391_,
		_w2401_,
		_w2534_
	);
	LUT4 #(
		.INIT('hab54)
	) name2501 (
		_w511_,
		_w2355_,
		_w2356_,
		_w2360_,
		_w2535_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name2502 (
		_w376_,
		_w486_,
		_w487_,
		_w509_,
		_w2536_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2503 (
		_w121_,
		_w418_,
		_w422_,
		_w2407_,
		_w2537_
	);
	LUT3 #(
		.INIT('h70)
	) name2504 (
		_w352_,
		_w373_,
		_w2527_,
		_w2538_
	);
	LUT3 #(
		.INIT('h01)
	) name2505 (
		_w2536_,
		_w2537_,
		_w2538_,
		_w2539_
	);
	LUT3 #(
		.INIT('h70)
	) name2506 (
		_w377_,
		_w2535_,
		_w2539_,
		_w2540_
	);
	LUT3 #(
		.INIT('he8)
	) name2507 (
		_w2533_,
		_w2534_,
		_w2540_,
		_w2541_
	);
	LUT4 #(
		.INIT('hc993)
	) name2508 (
		\a[29] ,
		_w330_,
		_w2391_,
		_w2401_,
		_w2542_
	);
	LUT3 #(
		.INIT('h4b)
	) name2509 (
		_w2405_,
		_w2409_,
		_w2542_,
		_w2543_
	);
	LUT2 #(
		.INIT('h4)
	) name2510 (
		_w2541_,
		_w2543_,
		_w2544_
	);
	LUT2 #(
		.INIT('h2)
	) name2511 (
		_w2541_,
		_w2543_,
		_w2545_
	);
	LUT2 #(
		.INIT('h9)
	) name2512 (
		_w2541_,
		_w2543_,
		_w2546_
	);
	LUT3 #(
		.INIT('h69)
	) name2513 (
		_w2533_,
		_w2534_,
		_w2540_,
		_w2547_
	);
	LUT2 #(
		.INIT('h9)
	) name2514 (
		\a[26] ,
		\a[27] ,
		_w2548_
	);
	LUT4 #(
		.INIT('h0180)
	) name2515 (
		\a[26] ,
		\a[27] ,
		\a[28] ,
		\a[29] ,
		_w2549_
	);
	LUT4 #(
		.INIT('h0660)
	) name2516 (
		\a[26] ,
		\a[27] ,
		\a[28] ,
		\a[29] ,
		_w2550_
	);
	LUT4 #(
		.INIT('h5150)
	) name2517 (
		_w374_,
		_w2361_,
		_w2549_,
		_w2550_,
		_w2551_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2518 (
		_w486_,
		_w487_,
		_w509_,
		_w2407_,
		_w2552_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2519 (
		_w121_,
		_w418_,
		_w422_,
		_w2527_,
		_w2553_
	);
	LUT3 #(
		.INIT('h2a)
	) name2520 (
		_w376_,
		_w544_,
		_w558_,
		_w2554_
	);
	LUT3 #(
		.INIT('h01)
	) name2521 (
		_w2552_,
		_w2553_,
		_w2554_,
		_w2555_
	);
	LUT4 #(
		.INIT('h7d00)
	) name2522 (
		_w377_,
		_w2355_,
		_w2357_,
		_w2555_,
		_w2556_
	);
	LUT3 #(
		.INIT('h56)
	) name2523 (
		_w2449_,
		_w2524_,
		_w2532_,
		_w2557_
	);
	LUT4 #(
		.INIT('h6f06)
	) name2524 (
		\a[29] ,
		_w2551_,
		_w2556_,
		_w2557_,
		_w2558_
	);
	LUT2 #(
		.INIT('h8)
	) name2525 (
		_w2547_,
		_w2558_,
		_w2559_
	);
	LUT4 #(
		.INIT('h153f)
	) name2526 (
		_w47_,
		_w65_,
		_w176_,
		_w430_,
		_w2560_
	);
	LUT4 #(
		.INIT('h135f)
	) name2527 (
		_w106_,
		_w52_,
		_w56_,
		_w184_,
		_w2561_
	);
	LUT4 #(
		.INIT('h8000)
	) name2528 (
		_w96_,
		_w1656_,
		_w2560_,
		_w2561_,
		_w2562_
	);
	LUT4 #(
		.INIT('h135f)
	) name2529 (
		_w78_,
		_w90_,
		_w50_,
		_w184_,
		_w2563_
	);
	LUT4 #(
		.INIT('h0200)
	) name2530 (
		_w130_,
		_w74_,
		_w386_,
		_w2563_,
		_w2564_
	);
	LUT2 #(
		.INIT('h8)
	) name2531 (
		_w2562_,
		_w2564_,
		_w2565_
	);
	LUT3 #(
		.INIT('h80)
	) name2532 (
		_w1077_,
		_w1086_,
		_w2565_,
		_w2566_
	);
	LUT3 #(
		.INIT('h80)
	) name2533 (
		_w662_,
		_w1416_,
		_w1587_,
		_w2567_
	);
	LUT4 #(
		.INIT('h0777)
	) name2534 (
		_w78_,
		_w90_,
		_w44_,
		_w158_,
		_w2568_
	);
	LUT4 #(
		.INIT('h8000)
	) name2535 (
		_w132_,
		_w260_,
		_w490_,
		_w2568_,
		_w2569_
	);
	LUT4 #(
		.INIT('h135f)
	) name2536 (
		_w106_,
		_w55_,
		_w110_,
		_w236_,
		_w2570_
	);
	LUT4 #(
		.INIT('h4000)
	) name2537 (
		_w407_,
		_w1026_,
		_w1027_,
		_w2570_,
		_w2571_
	);
	LUT3 #(
		.INIT('h80)
	) name2538 (
		_w2567_,
		_w2569_,
		_w2571_,
		_w2572_
	);
	LUT4 #(
		.INIT('h153f)
	) name2539 (
		_w47_,
		_w72_,
		_w93_,
		_w166_,
		_w2573_
	);
	LUT4 #(
		.INIT('h0777)
	) name2540 (
		_w90_,
		_w43_,
		_w46_,
		_w236_,
		_w2574_
	);
	LUT3 #(
		.INIT('h80)
	) name2541 (
		_w474_,
		_w2573_,
		_w2574_,
		_w2575_
	);
	LUT4 #(
		.INIT('h135f)
	) name2542 (
		_w52_,
		_w110_,
		_w78_,
		_w39_,
		_w2576_
	);
	LUT3 #(
		.INIT('h80)
	) name2543 (
		_w1974_,
		_w2140_,
		_w2576_,
		_w2577_
	);
	LUT3 #(
		.INIT('h80)
	) name2544 (
		_w1582_,
		_w2575_,
		_w2577_,
		_w2578_
	);
	LUT4 #(
		.INIT('h153f)
	) name2545 (
		_w59_,
		_w39_,
		_w65_,
		_w176_,
		_w2579_
	);
	LUT2 #(
		.INIT('h4)
	) name2546 (
		_w443_,
		_w2579_,
		_w2580_
	);
	LUT3 #(
		.INIT('h57)
	) name2547 (
		_w56_,
		_w419_,
		_w430_,
		_w2581_
	);
	LUT4 #(
		.INIT('h135f)
	) name2548 (
		_w55_,
		_w59_,
		_w39_,
		_w430_,
		_w2582_
	);
	LUT4 #(
		.INIT('h4000)
	) name2549 (
		_w186_,
		_w1931_,
		_w2581_,
		_w2582_,
		_w2583_
	);
	LUT4 #(
		.INIT('h0777)
	) name2550 (
		_w78_,
		_w56_,
		_w44_,
		_w184_,
		_w2584_
	);
	LUT2 #(
		.INIT('h4)
	) name2551 (
		_w194_,
		_w2584_,
		_w2585_
	);
	LUT4 #(
		.INIT('h2000)
	) name2552 (
		_w54_,
		_w205_,
		_w956_,
		_w1986_,
		_w2586_
	);
	LUT4 #(
		.INIT('h8000)
	) name2553 (
		_w2585_,
		_w2580_,
		_w2583_,
		_w2586_,
		_w2587_
	);
	LUT3 #(
		.INIT('h80)
	) name2554 (
		_w2572_,
		_w2578_,
		_w2587_,
		_w2588_
	);
	LUT4 #(
		.INIT('h8000)
	) name2555 (
		_w367_,
		_w514_,
		_w1683_,
		_w2495_,
		_w2589_
	);
	LUT2 #(
		.INIT('h4)
	) name2556 (
		_w230_,
		_w2235_,
		_w2590_
	);
	LUT4 #(
		.INIT('h153f)
	) name2557 (
		_w38_,
		_w122_,
		_w41_,
		_w39_,
		_w2591_
	);
	LUT4 #(
		.INIT('h135f)
	) name2558 (
		_w122_,
		_w44_,
		_w46_,
		_w378_,
		_w2592_
	);
	LUT4 #(
		.INIT('h8000)
	) name2559 (
		_w496_,
		_w806_,
		_w2591_,
		_w2592_,
		_w2593_
	);
	LUT3 #(
		.INIT('h80)
	) name2560 (
		_w2590_,
		_w2589_,
		_w2593_,
		_w2594_
	);
	LUT4 #(
		.INIT('h8000)
	) name2561 (
		_w2572_,
		_w2578_,
		_w2587_,
		_w2594_,
		_w2595_
	);
	LUT4 #(
		.INIT('h0888)
	) name2562 (
		_w1584_,
		_w2482_,
		_w2566_,
		_w2595_,
		_w2596_
	);
	LUT4 #(
		.INIT('h8777)
	) name2563 (
		_w1584_,
		_w2482_,
		_w2566_,
		_w2595_,
		_w2597_
	);
	LUT4 #(
		.INIT('h54ab)
	) name2564 (
		_w766_,
		_w2347_,
		_w2348_,
		_w2350_,
		_w2598_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2565 (
		_w587_,
		_w608_,
		_w624_,
		_w2527_,
		_w2599_
	);
	LUT3 #(
		.INIT('h2a)
	) name2566 (
		_w376_,
		_w725_,
		_w764_,
		_w2600_
	);
	LUT3 #(
		.INIT('h70)
	) name2567 (
		_w666_,
		_w694_,
		_w2407_,
		_w2601_
	);
	LUT3 #(
		.INIT('h01)
	) name2568 (
		_w2600_,
		_w2601_,
		_w2599_,
		_w2602_
	);
	LUT4 #(
		.INIT('h80cc)
	) name2569 (
		_w377_,
		_w2597_,
		_w2598_,
		_w2602_,
		_w2603_
	);
	LUT3 #(
		.INIT('ha9)
	) name2570 (
		\a[26] ,
		_w2522_,
		_w2523_,
		_w2604_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2571 (
		_w587_,
		_w608_,
		_w624_,
		_w2407_,
		_w2605_
	);
	LUT3 #(
		.INIT('h2a)
	) name2572 (
		_w376_,
		_w666_,
		_w694_,
		_w2606_
	);
	LUT3 #(
		.INIT('h70)
	) name2573 (
		_w544_,
		_w558_,
		_w2527_,
		_w2607_
	);
	LUT3 #(
		.INIT('h01)
	) name2574 (
		_w2606_,
		_w2607_,
		_w2605_,
		_w2608_
	);
	LUT4 #(
		.INIT('h7d00)
	) name2575 (
		_w377_,
		_w2351_,
		_w2353_,
		_w2608_,
		_w2609_
	);
	LUT4 #(
		.INIT('hf110)
	) name2576 (
		_w2596_,
		_w2603_,
		_w2604_,
		_w2609_,
		_w2610_
	);
	LUT4 #(
		.INIT('h3c39)
	) name2577 (
		\a[26] ,
		_w2447_,
		_w2522_,
		_w2523_,
		_w2611_
	);
	LUT4 #(
		.INIT('h708f)
	) name2578 (
		_w377_,
		_w2526_,
		_w2531_,
		_w2611_,
		_w2612_
	);
	LUT2 #(
		.INIT('h4)
	) name2579 (
		_w2610_,
		_w2612_,
		_w2613_
	);
	LUT2 #(
		.INIT('h2)
	) name2580 (
		_w2610_,
		_w2612_,
		_w2614_
	);
	LUT4 #(
		.INIT('hf400)
	) name2581 (
		_w374_,
		_w2361_,
		_w2404_,
		_w2550_,
		_w2615_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2582 (
		_w121_,
		_w418_,
		_w422_,
		_w2549_,
		_w2616_
	);
	LUT3 #(
		.INIT('h18)
	) name2583 (
		\a[26] ,
		\a[27] ,
		\a[28] ,
		_w2617_
	);
	LUT3 #(
		.INIT('h70)
	) name2584 (
		_w352_,
		_w373_,
		_w2617_,
		_w2618_
	);
	LUT2 #(
		.INIT('h1)
	) name2585 (
		_w2616_,
		_w2618_,
		_w2619_
	);
	LUT4 #(
		.INIT('h1211)
	) name2586 (
		\a[29] ,
		_w2614_,
		_w2615_,
		_w2619_,
		_w2620_
	);
	LUT4 #(
		.INIT('h6996)
	) name2587 (
		\a[29] ,
		_w2551_,
		_w2556_,
		_w2557_,
		_w2621_
	);
	LUT3 #(
		.INIT('h0e)
	) name2588 (
		_w2613_,
		_w2620_,
		_w2621_,
		_w2622_
	);
	LUT4 #(
		.INIT('h6c33)
	) name2589 (
		_w377_,
		_w2597_,
		_w2598_,
		_w2602_,
		_w2623_
	);
	LUT4 #(
		.INIT('h135f)
	) name2590 (
		_w47_,
		_w50_,
		_w201_,
		_w378_,
		_w2624_
	);
	LUT4 #(
		.INIT('h153f)
	) name2591 (
		_w55_,
		_w78_,
		_w65_,
		_w184_,
		_w2625_
	);
	LUT3 #(
		.INIT('h80)
	) name2592 (
		_w886_,
		_w2625_,
		_w2624_,
		_w2626_
	);
	LUT4 #(
		.INIT('h135f)
	) name2593 (
		_w106_,
		_w85_,
		_w50_,
		_w158_,
		_w2627_
	);
	LUT4 #(
		.INIT('h0777)
	) name2594 (
		_w122_,
		_w67_,
		_w90_,
		_w158_,
		_w2628_
	);
	LUT4 #(
		.INIT('h4000)
	) name2595 (
		_w478_,
		_w698_,
		_w2628_,
		_w2627_,
		_w2629_
	);
	LUT4 #(
		.INIT('h4000)
	) name2596 (
		_w380_,
		_w824_,
		_w825_,
		_w1521_,
		_w2630_
	);
	LUT3 #(
		.INIT('h80)
	) name2597 (
		_w2626_,
		_w2629_,
		_w2630_,
		_w2631_
	);
	LUT4 #(
		.INIT('h0777)
	) name2598 (
		_w106_,
		_w67_,
		_w41_,
		_w43_,
		_w2632_
	);
	LUT3 #(
		.INIT('h80)
	) name2599 (
		_w974_,
		_w1748_,
		_w2632_,
		_w2633_
	);
	LUT4 #(
		.INIT('h0777)
	) name2600 (
		_w85_,
		_w78_,
		_w90_,
		_w259_,
		_w2634_
	);
	LUT4 #(
		.INIT('h1000)
	) name2601 (
		_w321_,
		_w354_,
		_w790_,
		_w2634_,
		_w2635_
	);
	LUT4 #(
		.INIT('h8000)
	) name2602 (
		_w2201_,
		_w2202_,
		_w2633_,
		_w2635_,
		_w2636_
	);
	LUT4 #(
		.INIT('h153f)
	) name2603 (
		_w47_,
		_w44_,
		_w201_,
		_w166_,
		_w2637_
	);
	LUT4 #(
		.INIT('h135f)
	) name2604 (
		_w122_,
		_w55_,
		_w93_,
		_w166_,
		_w2638_
	);
	LUT2 #(
		.INIT('h8)
	) name2605 (
		_w2637_,
		_w2638_,
		_w2639_
	);
	LUT4 #(
		.INIT('h135f)
	) name2606 (
		_w67_,
		_w90_,
		_w184_,
		_w419_,
		_w2640_
	);
	LUT3 #(
		.INIT('h80)
	) name2607 (
		_w808_,
		_w1455_,
		_w2640_,
		_w2641_
	);
	LUT4 #(
		.INIT('h0777)
	) name2608 (
		_w52_,
		_w78_,
		_w56_,
		_w166_,
		_w2642_
	);
	LUT2 #(
		.INIT('h4)
	) name2609 (
		_w382_,
		_w2642_,
		_w2643_
	);
	LUT4 #(
		.INIT('h0777)
	) name2610 (
		_w110_,
		_w72_,
		_w65_,
		_w378_,
		_w2644_
	);
	LUT3 #(
		.INIT('h80)
	) name2611 (
		_w54_,
		_w2516_,
		_w2644_,
		_w2645_
	);
	LUT2 #(
		.INIT('h8)
	) name2612 (
		_w2643_,
		_w2645_,
		_w2646_
	);
	LUT4 #(
		.INIT('h8000)
	) name2613 (
		_w2639_,
		_w2641_,
		_w2643_,
		_w2645_,
		_w2647_
	);
	LUT3 #(
		.INIT('h80)
	) name2614 (
		_w2631_,
		_w2636_,
		_w2647_,
		_w2648_
	);
	LUT4 #(
		.INIT('h153f)
	) name2615 (
		_w52_,
		_w47_,
		_w39_,
		_w176_,
		_w2649_
	);
	LUT2 #(
		.INIT('h8)
	) name2616 (
		_w1514_,
		_w2649_,
		_w2650_
	);
	LUT4 #(
		.INIT('h0777)
	) name2617 (
		_w122_,
		_w41_,
		_w44_,
		_w158_,
		_w2651_
	);
	LUT4 #(
		.INIT('h153f)
	) name2618 (
		_w110_,
		_w65_,
		_w236_,
		_w419_,
		_w2652_
	);
	LUT4 #(
		.INIT('h4000)
	) name2619 (
		_w261_,
		_w760_,
		_w2651_,
		_w2652_,
		_w2653_
	);
	LUT4 #(
		.INIT('h153f)
	) name2620 (
		_w90_,
		_w47_,
		_w43_,
		_w176_,
		_w2654_
	);
	LUT4 #(
		.INIT('h135f)
	) name2621 (
		_w106_,
		_w78_,
		_w41_,
		_w46_,
		_w2655_
	);
	LUT3 #(
		.INIT('h40)
	) name2622 (
		_w424_,
		_w2654_,
		_w2655_,
		_w2656_
	);
	LUT4 #(
		.INIT('h8000)
	) name2623 (
		_w238_,
		_w1124_,
		_w1519_,
		_w1837_,
		_w2657_
	);
	LUT4 #(
		.INIT('h8000)
	) name2624 (
		_w2650_,
		_w2656_,
		_w2657_,
		_w2653_,
		_w2658_
	);
	LUT4 #(
		.INIT('h135f)
	) name2625 (
		_w56_,
		_w41_,
		_w43_,
		_w184_,
		_w2659_
	);
	LUT2 #(
		.INIT('h4)
	) name2626 (
		_w461_,
		_w2659_,
		_w2660_
	);
	LUT3 #(
		.INIT('h57)
	) name2627 (
		_w59_,
		_w236_,
		_w158_,
		_w2661_
	);
	LUT4 #(
		.INIT('h153f)
	) name2628 (
		_w110_,
		_w67_,
		_w201_,
		_w176_,
		_w2662_
	);
	LUT3 #(
		.INIT('h80)
	) name2629 (
		_w348_,
		_w2662_,
		_w2661_,
		_w2663_
	);
	LUT4 #(
		.INIT('h8000)
	) name2630 (
		_w1449_,
		_w1452_,
		_w2660_,
		_w2663_,
		_w2664_
	);
	LUT2 #(
		.INIT('h8)
	) name2631 (
		_w2658_,
		_w2664_,
		_w2665_
	);
	LUT2 #(
		.INIT('h8)
	) name2632 (
		_w2648_,
		_w2665_,
		_w2666_
	);
	LUT4 #(
		.INIT('h153f)
	) name2633 (
		_w38_,
		_w67_,
		_w259_,
		_w176_,
		_w2667_
	);
	LUT3 #(
		.INIT('h40)
	) name2634 (
		_w354_,
		_w2457_,
		_w2667_,
		_w2668_
	);
	LUT4 #(
		.INIT('h0777)
	) name2635 (
		_w38_,
		_w122_,
		_w106_,
		_w110_,
		_w2669_
	);
	LUT2 #(
		.INIT('h4)
	) name2636 (
		_w167_,
		_w2669_,
		_w2670_
	);
	LUT4 #(
		.INIT('h135f)
	) name2637 (
		_w38_,
		_w39_,
		_w43_,
		_w65_,
		_w2671_
	);
	LUT4 #(
		.INIT('h135f)
	) name2638 (
		_w106_,
		_w55_,
		_w41_,
		_w39_,
		_w2672_
	);
	LUT4 #(
		.INIT('h4000)
	) name2639 (
		_w167_,
		_w2669_,
		_w2671_,
		_w2672_,
		_w2673_
	);
	LUT2 #(
		.INIT('h8)
	) name2640 (
		_w2668_,
		_w2673_,
		_w2674_
	);
	LUT3 #(
		.INIT('h80)
	) name2641 (
		_w1004_,
		_w1182_,
		_w1910_,
		_w2675_
	);
	LUT4 #(
		.INIT('h8000)
	) name2642 (
		_w296_,
		_w527_,
		_w521_,
		_w660_,
		_w2676_
	);
	LUT3 #(
		.INIT('h80)
	) name2643 (
		_w733_,
		_w2675_,
		_w2676_,
		_w2677_
	);
	LUT4 #(
		.INIT('h8000)
	) name2644 (
		_w1198_,
		_w1403_,
		_w1651_,
		_w1844_,
		_w2678_
	);
	LUT4 #(
		.INIT('h153f)
	) name2645 (
		_w67_,
		_w50_,
		_w166_,
		_w430_,
		_w2679_
	);
	LUT4 #(
		.INIT('h8000)
	) name2646 (
		_w68_,
		_w222_,
		_w1337_,
		_w2679_,
		_w2680_
	);
	LUT4 #(
		.INIT('h8000)
	) name2647 (
		_w862_,
		_w2501_,
		_w2680_,
		_w2678_,
		_w2681_
	);
	LUT4 #(
		.INIT('h153f)
	) name2648 (
		_w90_,
		_w65_,
		_w236_,
		_w378_,
		_w2682_
	);
	LUT2 #(
		.INIT('h4)
	) name2649 (
		_w431_,
		_w2682_,
		_w2683_
	);
	LUT4 #(
		.INIT('h0777)
	) name2650 (
		_w38_,
		_w78_,
		_w90_,
		_w43_,
		_w2684_
	);
	LUT4 #(
		.INIT('h8000)
	) name2651 (
		_w936_,
		_w1137_,
		_w1180_,
		_w2684_,
		_w2685_
	);
	LUT4 #(
		.INIT('h8000)
	) name2652 (
		_w1555_,
		_w1558_,
		_w2683_,
		_w2685_,
		_w2686_
	);
	LUT4 #(
		.INIT('h8000)
	) name2653 (
		_w2674_,
		_w2677_,
		_w2681_,
		_w2686_,
		_w2687_
	);
	LUT3 #(
		.INIT('h80)
	) name2654 (
		_w567_,
		_w857_,
		_w1982_,
		_w2688_
	);
	LUT4 #(
		.INIT('h135f)
	) name2655 (
		_w55_,
		_w67_,
		_w78_,
		_w184_,
		_w2689_
	);
	LUT3 #(
		.INIT('h40)
	) name2656 (
		_w323_,
		_w906_,
		_w2689_,
		_w2690_
	);
	LUT4 #(
		.INIT('h135f)
	) name2657 (
		_w65_,
		_w46_,
		_w201_,
		_w176_,
		_w2691_
	);
	LUT4 #(
		.INIT('h2000)
	) name2658 (
		_w130_,
		_w478_,
		_w2169_,
		_w2691_,
		_w2692_
	);
	LUT3 #(
		.INIT('h80)
	) name2659 (
		_w2690_,
		_w2688_,
		_w2692_,
		_w2693_
	);
	LUT4 #(
		.INIT('h135f)
	) name2660 (
		_w55_,
		_w85_,
		_w378_,
		_w430_,
		_w2694_
	);
	LUT2 #(
		.INIT('h8)
	) name2661 (
		_w1415_,
		_w2694_,
		_w2695_
	);
	LUT4 #(
		.INIT('h135f)
	) name2662 (
		_w55_,
		_w72_,
		_w43_,
		_w65_,
		_w2696_
	);
	LUT3 #(
		.INIT('h80)
	) name2663 (
		_w1603_,
		_w2370_,
		_w2696_,
		_w2697_
	);
	LUT2 #(
		.INIT('h8)
	) name2664 (
		_w2695_,
		_w2697_,
		_w2698_
	);
	LUT4 #(
		.INIT('h135f)
	) name2665 (
		_w55_,
		_w90_,
		_w166_,
		_w158_,
		_w2699_
	);
	LUT3 #(
		.INIT('h1f)
	) name2666 (
		_w110_,
		_w56_,
		_w72_,
		_w2700_
	);
	LUT4 #(
		.INIT('h4000)
	) name2667 (
		_w389_,
		_w979_,
		_w2700_,
		_w2699_,
		_w2701_
	);
	LUT4 #(
		.INIT('h153f)
	) name2668 (
		_w122_,
		_w59_,
		_w39_,
		_w50_,
		_w2702_
	);
	LUT4 #(
		.INIT('h135f)
	) name2669 (
		_w106_,
		_w52_,
		_w50_,
		_w430_,
		_w2703_
	);
	LUT4 #(
		.INIT('h4000)
	) name2670 (
		_w451_,
		_w1122_,
		_w2702_,
		_w2703_,
		_w2704_
	);
	LUT4 #(
		.INIT('h153f)
	) name2671 (
		_w59_,
		_w41_,
		_w39_,
		_w430_,
		_w2705_
	);
	LUT4 #(
		.INIT('h135f)
	) name2672 (
		_w90_,
		_w50_,
		_w259_,
		_w419_,
		_w2706_
	);
	LUT3 #(
		.INIT('h80)
	) name2673 (
		_w1132_,
		_w2706_,
		_w2705_,
		_w2707_
	);
	LUT4 #(
		.INIT('h8000)
	) name2674 (
		_w1322_,
		_w2707_,
		_w2701_,
		_w2704_,
		_w2708_
	);
	LUT3 #(
		.INIT('h80)
	) name2675 (
		_w2693_,
		_w2698_,
		_w2708_,
		_w2709_
	);
	LUT2 #(
		.INIT('h8)
	) name2676 (
		_w2687_,
		_w2709_,
		_w2710_
	);
	LUT4 #(
		.INIT('h0777)
	) name2677 (
		_w2648_,
		_w2665_,
		_w2687_,
		_w2709_,
		_w2711_
	);
	LUT4 #(
		.INIT('h8000)
	) name2678 (
		_w2648_,
		_w2665_,
		_w2687_,
		_w2709_,
		_w2712_
	);
	LUT4 #(
		.INIT('h3220)
	) name2679 (
		\a[23] ,
		_w2483_,
		_w2666_,
		_w2710_,
		_w2713_
	);
	LUT4 #(
		.INIT('h044c)
	) name2680 (
		\a[23] ,
		_w2483_,
		_w2666_,
		_w2710_,
		_w2714_
	);
	LUT3 #(
		.INIT('h70)
	) name2681 (
		_w725_,
		_w764_,
		_w2407_,
		_w2715_
	);
	LUT3 #(
		.INIT('h2a)
	) name2682 (
		_w376_,
		_w801_,
		_w851_,
		_w2716_
	);
	LUT3 #(
		.INIT('h70)
	) name2683 (
		_w666_,
		_w694_,
		_w2527_,
		_w2717_
	);
	LUT3 #(
		.INIT('h01)
	) name2684 (
		_w2716_,
		_w2717_,
		_w2715_,
		_w2718_
	);
	LUT4 #(
		.INIT('h7d00)
	) name2685 (
		_w377_,
		_w2347_,
		_w2349_,
		_w2718_,
		_w2719_
	);
	LUT3 #(
		.INIT('h45)
	) name2686 (
		_w2713_,
		_w2714_,
		_w2719_,
		_w2720_
	);
	LUT2 #(
		.INIT('h8)
	) name2687 (
		_w2623_,
		_w2720_,
		_w2721_
	);
	LUT2 #(
		.INIT('h6)
	) name2688 (
		_w2623_,
		_w2720_,
		_w2722_
	);
	LUT3 #(
		.INIT('ha9)
	) name2689 (
		\a[23] ,
		_w2711_,
		_w2712_,
		_w2723_
	);
	LUT4 #(
		.INIT('h54ab)
	) name2690 (
		_w929_,
		_w2343_,
		_w2344_,
		_w2346_,
		_w2724_
	);
	LUT3 #(
		.INIT('h70)
	) name2691 (
		_w725_,
		_w764_,
		_w2527_,
		_w2725_
	);
	LUT3 #(
		.INIT('h70)
	) name2692 (
		_w801_,
		_w851_,
		_w2407_,
		_w2726_
	);
	LUT3 #(
		.INIT('h2a)
	) name2693 (
		_w376_,
		_w871_,
		_w927_,
		_w2727_
	);
	LUT3 #(
		.INIT('h01)
	) name2694 (
		_w2726_,
		_w2727_,
		_w2725_,
		_w2728_
	);
	LUT4 #(
		.INIT('h2033)
	) name2695 (
		_w377_,
		_w2723_,
		_w2724_,
		_w2728_,
		_w2729_
	);
	LUT2 #(
		.INIT('h2)
	) name2696 (
		_w240_,
		_w424_,
		_w2730_
	);
	LUT4 #(
		.INIT('h153f)
	) name2697 (
		_w56_,
		_w47_,
		_w39_,
		_w430_,
		_w2731_
	);
	LUT3 #(
		.INIT('h80)
	) name2698 (
		_w1351_,
		_w1429_,
		_w2731_,
		_w2732_
	);
	LUT2 #(
		.INIT('h8)
	) name2699 (
		_w2730_,
		_w2732_,
		_w2733_
	);
	LUT4 #(
		.INIT('h8000)
	) name2700 (
		_w949_,
		_w1060_,
		_w1158_,
		_w1785_,
		_w2734_
	);
	LUT4 #(
		.INIT('h135f)
	) name2701 (
		_w78_,
		_w50_,
		_w44_,
		_w166_,
		_w2735_
	);
	LUT4 #(
		.INIT('h4000)
	) name2702 (
		_w440_,
		_w834_,
		_w1047_,
		_w2735_,
		_w2736_
	);
	LUT4 #(
		.INIT('h135f)
	) name2703 (
		_w106_,
		_w90_,
		_w46_,
		_w236_,
		_w2737_
	);
	LUT3 #(
		.INIT('h40)
	) name2704 (
		_w379_,
		_w512_,
		_w2737_,
		_w2738_
	);
	LUT4 #(
		.INIT('h8000)
	) name2705 (
		_w1032_,
		_w2738_,
		_w2734_,
		_w2736_,
		_w2739_
	);
	LUT3 #(
		.INIT('h80)
	) name2706 (
		_w1213_,
		_w2733_,
		_w2739_,
		_w2740_
	);
	LUT4 #(
		.INIT('h135f)
	) name2707 (
		_w67_,
		_w90_,
		_w201_,
		_w158_,
		_w2741_
	);
	LUT4 #(
		.INIT('h4000)
	) name2708 (
		_w97_,
		_w1891_,
		_w2364_,
		_w2741_,
		_w2742_
	);
	LUT2 #(
		.INIT('h8)
	) name2709 (
		_w2230_,
		_w2742_,
		_w2743_
	);
	LUT4 #(
		.INIT('h135f)
	) name2710 (
		_w106_,
		_w55_,
		_w93_,
		_w166_,
		_w2744_
	);
	LUT3 #(
		.INIT('h57)
	) name2711 (
		_w110_,
		_w184_,
		_w236_,
		_w2745_
	);
	LUT4 #(
		.INIT('h8000)
	) name2712 (
		_w609_,
		_w957_,
		_w2744_,
		_w2745_,
		_w2746_
	);
	LUT4 #(
		.INIT('h153f)
	) name2713 (
		_w41_,
		_w46_,
		_w236_,
		_w259_,
		_w2747_
	);
	LUT4 #(
		.INIT('h4000)
	) name2714 (
		_w291_,
		_w518_,
		_w584_,
		_w2747_,
		_w2748_
	);
	LUT4 #(
		.INIT('h135f)
	) name2715 (
		_w122_,
		_w65_,
		_w46_,
		_w184_,
		_w2749_
	);
	LUT4 #(
		.INIT('h2000)
	) name2716 (
		_w68_,
		_w392_,
		_w1761_,
		_w2749_,
		_w2750_
	);
	LUT3 #(
		.INIT('h80)
	) name2717 (
		_w2746_,
		_w2748_,
		_w2750_,
		_w2751_
	);
	LUT4 #(
		.INIT('h8000)
	) name2718 (
		_w2029_,
		_w2035_,
		_w2743_,
		_w2751_,
		_w2752_
	);
	LUT2 #(
		.INIT('h8)
	) name2719 (
		_w2740_,
		_w2752_,
		_w2753_
	);
	LUT4 #(
		.INIT('h0888)
	) name2720 (
		_w2648_,
		_w2665_,
		_w2740_,
		_w2752_,
		_w2754_
	);
	LUT4 #(
		.INIT('h8777)
	) name2721 (
		_w2648_,
		_w2665_,
		_w2740_,
		_w2752_,
		_w2755_
	);
	LUT2 #(
		.INIT('h8)
	) name2722 (
		_w944_,
		_w990_,
		_w2756_
	);
	LUT4 #(
		.INIT('h8000)
	) name2723 (
		_w1013_,
		_w1191_,
		_w1472_,
		_w1844_,
		_w2757_
	);
	LUT3 #(
		.INIT('h1f)
	) name2724 (
		_w41_,
		_w44_,
		_w184_,
		_w2758_
	);
	LUT3 #(
		.INIT('h80)
	) name2725 (
		_w817_,
		_w1091_,
		_w2758_,
		_w2759_
	);
	LUT4 #(
		.INIT('h153f)
	) name2726 (
		_w59_,
		_w72_,
		_w65_,
		_w430_,
		_w2760_
	);
	LUT4 #(
		.INIT('h4000)
	) name2727 (
		_w476_,
		_w479_,
		_w519_,
		_w2760_,
		_w2761_
	);
	LUT4 #(
		.INIT('h8000)
	) name2728 (
		_w2756_,
		_w2759_,
		_w2761_,
		_w2757_,
		_w2762_
	);
	LUT3 #(
		.INIT('h80)
	) name2729 (
		_w1313_,
		_w1553_,
		_w2762_,
		_w2763_
	);
	LUT4 #(
		.INIT('h135f)
	) name2730 (
		_w85_,
		_w44_,
		_w259_,
		_w176_,
		_w2764_
	);
	LUT4 #(
		.INIT('h8000)
	) name2731 (
		_w2274_,
		_w2460_,
		_w2493_,
		_w2764_,
		_w2765_
	);
	LUT3 #(
		.INIT('h1f)
	) name2732 (
		_w55_,
		_w52_,
		_w201_,
		_w2766_
	);
	LUT4 #(
		.INIT('h8000)
	) name2733 (
		_w96_,
		_w1045_,
		_w1726_,
		_w2766_,
		_w2767_
	);
	LUT3 #(
		.INIT('h80)
	) name2734 (
		_w2730_,
		_w2765_,
		_w2767_,
		_w2768_
	);
	LUT4 #(
		.INIT('h0777)
	) name2735 (
		_w122_,
		_w55_,
		_w90_,
		_w72_,
		_w2769_
	);
	LUT4 #(
		.INIT('h8000)
	) name2736 (
		_w809_,
		_w1124_,
		_w1935_,
		_w2769_,
		_w2770_
	);
	LUT4 #(
		.INIT('h135f)
	) name2737 (
		_w85_,
		_w65_,
		_w184_,
		_w419_,
		_w2771_
	);
	LUT4 #(
		.INIT('h1000)
	) name2738 (
		_w358_,
		_w379_,
		_w2415_,
		_w2771_,
		_w2772_
	);
	LUT2 #(
		.INIT('h8)
	) name2739 (
		_w2770_,
		_w2772_,
		_w2773_
	);
	LUT4 #(
		.INIT('h8000)
	) name2740 (
		_w1782_,
		_w1786_,
		_w2770_,
		_w2772_,
		_w2774_
	);
	LUT2 #(
		.INIT('h8)
	) name2741 (
		_w2768_,
		_w2774_,
		_w2775_
	);
	LUT4 #(
		.INIT('h0200)
	) name2742 (
		_w132_,
		_w253_,
		_w432_,
		_w1429_,
		_w2776_
	);
	LUT2 #(
		.INIT('h8)
	) name2743 (
		_w2289_,
		_w2776_,
		_w2777_
	);
	LUT3 #(
		.INIT('h80)
	) name2744 (
		_w651_,
		_w1519_,
		_w1761_,
		_w2778_
	);
	LUT4 #(
		.INIT('h153f)
	) name2745 (
		_w52_,
		_w72_,
		_w50_,
		_w236_,
		_w2779_
	);
	LUT4 #(
		.INIT('h2000)
	) name2746 (
		_w198_,
		_w360_,
		_w668_,
		_w2779_,
		_w2780_
	);
	LUT3 #(
		.INIT('h10)
	) name2747 (
		_w246_,
		_w167_,
		_w343_,
		_w2781_
	);
	LUT4 #(
		.INIT('h153f)
	) name2748 (
		_w110_,
		_w44_,
		_w236_,
		_w176_,
		_w2782_
	);
	LUT4 #(
		.INIT('h4000)
	) name2749 (
		_w276_,
		_w394_,
		_w1975_,
		_w2782_,
		_w2783_
	);
	LUT4 #(
		.INIT('h8000)
	) name2750 (
		_w2781_,
		_w2783_,
		_w2778_,
		_w2780_,
		_w2784_
	);
	LUT2 #(
		.INIT('h8)
	) name2751 (
		_w2777_,
		_w2784_,
		_w2785_
	);
	LUT4 #(
		.INIT('h8000)
	) name2752 (
		_w2768_,
		_w2774_,
		_w2777_,
		_w2784_,
		_w2786_
	);
	LUT2 #(
		.INIT('h8)
	) name2753 (
		_w2763_,
		_w2786_,
		_w2787_
	);
	LUT3 #(
		.INIT('h1f)
	) name2754 (
		_w90_,
		_w46_,
		_w166_,
		_w2788_
	);
	LUT3 #(
		.INIT('h40)
	) name2755 (
		_w355_,
		_w1438_,
		_w2788_,
		_w2789_
	);
	LUT4 #(
		.INIT('h153f)
	) name2756 (
		_w38_,
		_w55_,
		_w236_,
		_w378_,
		_w2790_
	);
	LUT4 #(
		.INIT('h4000)
	) name2757 (
		_w431_,
		_w863_,
		_w1401_,
		_w2790_,
		_w2791_
	);
	LUT4 #(
		.INIT('h1000)
	) name2758 (
		_w146_,
		_w308_,
		_w868_,
		_w1012_,
		_w2792_
	);
	LUT3 #(
		.INIT('h80)
	) name2759 (
		_w2789_,
		_w2791_,
		_w2792_,
		_w2793_
	);
	LUT4 #(
		.INIT('h0777)
	) name2760 (
		_w122_,
		_w67_,
		_w43_,
		_w44_,
		_w2794_
	);
	LUT4 #(
		.INIT('h8000)
	) name2761 (
		_w361_,
		_w533_,
		_w582_,
		_w2794_,
		_w2795_
	);
	LUT4 #(
		.INIT('h135f)
	) name2762 (
		_w50_,
		_w46_,
		_w166_,
		_w176_,
		_w2796_
	);
	LUT4 #(
		.INIT('h135f)
	) name2763 (
		_w106_,
		_w85_,
		_w90_,
		_w430_,
		_w2797_
	);
	LUT4 #(
		.INIT('h4000)
	) name2764 (
		_w74_,
		_w1014_,
		_w2796_,
		_w2797_,
		_w2798_
	);
	LUT4 #(
		.INIT('h8000)
	) name2765 (
		_w1601_,
		_w1604_,
		_w2795_,
		_w2798_,
		_w2799_
	);
	LUT2 #(
		.INIT('h8)
	) name2766 (
		_w2793_,
		_w2799_,
		_w2800_
	);
	LUT4 #(
		.INIT('h135f)
	) name2767 (
		_w56_,
		_w50_,
		_w378_,
		_w430_,
		_w2801_
	);
	LUT4 #(
		.INIT('h8000)
	) name2768 (
		_w148_,
		_w512_,
		_w678_,
		_w2801_,
		_w2802_
	);
	LUT4 #(
		.INIT('h153f)
	) name2769 (
		_w38_,
		_w106_,
		_w41_,
		_w39_,
		_w2803_
	);
	LUT4 #(
		.INIT('h8000)
	) name2770 (
		_w302_,
		_w839_,
		_w2706_,
		_w2803_,
		_w2804_
	);
	LUT2 #(
		.INIT('h8)
	) name2771 (
		_w2802_,
		_w2804_,
		_w2805_
	);
	LUT4 #(
		.INIT('h131f)
	) name2772 (
		_w38_,
		_w52_,
		_w184_,
		_w430_,
		_w2806_
	);
	LUT4 #(
		.INIT('h0777)
	) name2773 (
		_w122_,
		_w52_,
		_w93_,
		_w184_,
		_w2807_
	);
	LUT3 #(
		.INIT('h80)
	) name2774 (
		_w2258_,
		_w2807_,
		_w2806_,
		_w2808_
	);
	LUT4 #(
		.INIT('h135f)
	) name2775 (
		_w38_,
		_w85_,
		_w72_,
		_w419_,
		_w2809_
	);
	LUT4 #(
		.INIT('h153f)
	) name2776 (
		_w55_,
		_w110_,
		_w201_,
		_w166_,
		_w2810_
	);
	LUT3 #(
		.INIT('h80)
	) name2777 (
		_w2000_,
		_w2810_,
		_w2809_,
		_w2811_
	);
	LUT4 #(
		.INIT('h8000)
	) name2778 (
		_w944_,
		_w1158_,
		_w1334_,
		_w1362_,
		_w2812_
	);
	LUT3 #(
		.INIT('h80)
	) name2779 (
		_w2808_,
		_w2811_,
		_w2812_,
		_w2813_
	);
	LUT2 #(
		.INIT('h8)
	) name2780 (
		_w2805_,
		_w2813_,
		_w2814_
	);
	LUT4 #(
		.INIT('h8000)
	) name2781 (
		_w737_,
		_w808_,
		_w937_,
		_w1079_,
		_w2815_
	);
	LUT3 #(
		.INIT('h37)
	) name2782 (
		_w90_,
		_w72_,
		_w44_,
		_w2816_
	);
	LUT4 #(
		.INIT('h135f)
	) name2783 (
		_w106_,
		_w110_,
		_w47_,
		_w378_,
		_w2817_
	);
	LUT4 #(
		.INIT('h4000)
	) name2784 (
		_w241_,
		_w2044_,
		_w2816_,
		_w2817_,
		_w2818_
	);
	LUT3 #(
		.INIT('h80)
	) name2785 (
		_w684_,
		_w2815_,
		_w2818_,
		_w2819_
	);
	LUT4 #(
		.INIT('h0777)
	) name2786 (
		_w106_,
		_w55_,
		_w85_,
		_w259_,
		_w2820_
	);
	LUT2 #(
		.INIT('h8)
	) name2787 (
		_w95_,
		_w2820_,
		_w2821_
	);
	LUT4 #(
		.INIT('h0777)
	) name2788 (
		_w85_,
		_w78_,
		_w47_,
		_w72_,
		_w2822_
	);
	LUT4 #(
		.INIT('h135f)
	) name2789 (
		_w38_,
		_w52_,
		_w43_,
		_w166_,
		_w2823_
	);
	LUT4 #(
		.INIT('h8000)
	) name2790 (
		_w677_,
		_w2125_,
		_w2822_,
		_w2823_,
		_w2824_
	);
	LUT4 #(
		.INIT('h0777)
	) name2791 (
		_w41_,
		_w43_,
		_w93_,
		_w259_,
		_w2825_
	);
	LUT4 #(
		.INIT('h135f)
	) name2792 (
		_w93_,
		_w44_,
		_w236_,
		_w166_,
		_w2826_
	);
	LUT4 #(
		.INIT('h8000)
	) name2793 (
		_w387_,
		_w1245_,
		_w2825_,
		_w2826_,
		_w2827_
	);
	LUT4 #(
		.INIT('h135f)
	) name2794 (
		_w122_,
		_w106_,
		_w56_,
		_w93_,
		_w2828_
	);
	LUT4 #(
		.INIT('h0777)
	) name2795 (
		_w43_,
		_w93_,
		_w46_,
		_w184_,
		_w2829_
	);
	LUT4 #(
		.INIT('h153f)
	) name2796 (
		_w38_,
		_w56_,
		_w236_,
		_w158_,
		_w2830_
	);
	LUT4 #(
		.INIT('h4000)
	) name2797 (
		_w458_,
		_w2829_,
		_w2830_,
		_w2828_,
		_w2831_
	);
	LUT4 #(
		.INIT('h8000)
	) name2798 (
		_w2821_,
		_w2824_,
		_w2827_,
		_w2831_,
		_w2832_
	);
	LUT4 #(
		.INIT('h8000)
	) name2799 (
		_w2805_,
		_w2813_,
		_w2819_,
		_w2832_,
		_w2833_
	);
	LUT2 #(
		.INIT('h8)
	) name2800 (
		_w2800_,
		_w2833_,
		_w2834_
	);
	LUT4 #(
		.INIT('h0777)
	) name2801 (
		_w2763_,
		_w2786_,
		_w2800_,
		_w2833_,
		_w2835_
	);
	LUT4 #(
		.INIT('h8000)
	) name2802 (
		_w2763_,
		_w2786_,
		_w2800_,
		_w2833_,
		_w2836_
	);
	LUT4 #(
		.INIT('h3220)
	) name2803 (
		\a[20] ,
		_w2753_,
		_w2787_,
		_w2834_,
		_w2837_
	);
	LUT4 #(
		.INIT('h044c)
	) name2804 (
		\a[20] ,
		_w2753_,
		_w2787_,
		_w2834_,
		_w2838_
	);
	LUT4 #(
		.INIT('h54ab)
	) name2805 (
		_w1052_,
		_w2339_,
		_w2340_,
		_w2342_,
		_w2839_
	);
	LUT3 #(
		.INIT('h2a)
	) name2806 (
		_w376_,
		_w1009_,
		_w1050_,
		_w2840_
	);
	LUT3 #(
		.INIT('h70)
	) name2807 (
		_w871_,
		_w927_,
		_w2527_,
		_w2841_
	);
	LUT3 #(
		.INIT('h70)
	) name2808 (
		_w763_,
		_w983_,
		_w2407_,
		_w2842_
	);
	LUT3 #(
		.INIT('h01)
	) name2809 (
		_w2841_,
		_w2842_,
		_w2840_,
		_w2843_
	);
	LUT4 #(
		.INIT('h1300)
	) name2810 (
		_w377_,
		_w2838_,
		_w2839_,
		_w2843_,
		_w2844_
	);
	LUT4 #(
		.INIT('h5551)
	) name2811 (
		_w2754_,
		_w2755_,
		_w2837_,
		_w2844_,
		_w2845_
	);
	LUT4 #(
		.INIT('h4c00)
	) name2812 (
		_w377_,
		_w2723_,
		_w2724_,
		_w2728_,
		_w2846_
	);
	LUT4 #(
		.INIT('h93cc)
	) name2813 (
		_w377_,
		_w2723_,
		_w2724_,
		_w2728_,
		_w2847_
	);
	LUT3 #(
		.INIT('h54)
	) name2814 (
		_w2729_,
		_w2845_,
		_w2846_,
		_w2848_
	);
	LUT4 #(
		.INIT('h3c39)
	) name2815 (
		\a[23] ,
		_w2483_,
		_w2711_,
		_w2712_,
		_w2849_
	);
	LUT2 #(
		.INIT('h9)
	) name2816 (
		_w2719_,
		_w2849_,
		_w2850_
	);
	LUT2 #(
		.INIT('h4)
	) name2817 (
		_w2848_,
		_w2850_,
		_w2851_
	);
	LUT2 #(
		.INIT('h2)
	) name2818 (
		_w2848_,
		_w2850_,
		_w2852_
	);
	LUT2 #(
		.INIT('h9)
	) name2819 (
		_w2848_,
		_w2850_,
		_w2853_
	);
	LUT4 #(
		.INIT('h6006)
	) name2820 (
		\a[26] ,
		\a[27] ,
		\a[28] ,
		\a[29] ,
		_w2854_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2821 (
		_w486_,
		_w487_,
		_w509_,
		_w2854_,
		_w2855_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2822 (
		_w587_,
		_w608_,
		_w624_,
		_w2549_,
		_w2856_
	);
	LUT3 #(
		.INIT('h70)
	) name2823 (
		_w544_,
		_w558_,
		_w2617_,
		_w2857_
	);
	LUT3 #(
		.INIT('h01)
	) name2824 (
		_w2855_,
		_w2856_,
		_w2857_,
		_w2858_
	);
	LUT4 #(
		.INIT('h95aa)
	) name2825 (
		\a[29] ,
		_w2526_,
		_w2550_,
		_w2858_,
		_w2859_
	);
	LUT4 #(
		.INIT('h20a2)
	) name2826 (
		_w2722_,
		_w2848_,
		_w2850_,
		_w2859_,
		_w2860_
	);
	LUT4 #(
		.INIT('he11e)
	) name2827 (
		_w2596_,
		_w2603_,
		_w2604_,
		_w2609_,
		_w2861_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2828 (
		_w486_,
		_w487_,
		_w509_,
		_w2549_,
		_w2862_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2829 (
		_w121_,
		_w418_,
		_w422_,
		_w2617_,
		_w2863_
	);
	LUT3 #(
		.INIT('h70)
	) name2830 (
		_w352_,
		_w373_,
		_w2854_,
		_w2864_
	);
	LUT3 #(
		.INIT('h01)
	) name2831 (
		_w2862_,
		_w2863_,
		_w2864_,
		_w2865_
	);
	LUT4 #(
		.INIT('h95aa)
	) name2832 (
		\a[29] ,
		_w2535_,
		_w2550_,
		_w2865_,
		_w2866_
	);
	LUT4 #(
		.INIT('h1f01)
	) name2833 (
		_w2721_,
		_w2860_,
		_w2861_,
		_w2866_,
		_w2867_
	);
	LUT2 #(
		.INIT('h9)
	) name2834 (
		_w2610_,
		_w2612_,
		_w2868_
	);
	LUT4 #(
		.INIT('h9a65)
	) name2835 (
		\a[29] ,
		_w2615_,
		_w2619_,
		_w2868_,
		_w2869_
	);
	LUT2 #(
		.INIT('h4)
	) name2836 (
		_w2867_,
		_w2869_,
		_w2870_
	);
	LUT2 #(
		.INIT('h2)
	) name2837 (
		_w2867_,
		_w2869_,
		_w2871_
	);
	LUT2 #(
		.INIT('h9)
	) name2838 (
		_w2867_,
		_w2869_,
		_w2872_
	);
	LUT2 #(
		.INIT('h9)
	) name2839 (
		\a[23] ,
		\a[24] ,
		_w2873_
	);
	LUT4 #(
		.INIT('h0180)
	) name2840 (
		\a[23] ,
		\a[24] ,
		\a[25] ,
		\a[26] ,
		_w2874_
	);
	LUT4 #(
		.INIT('h0660)
	) name2841 (
		\a[23] ,
		\a[24] ,
		\a[25] ,
		\a[26] ,
		_w2875_
	);
	LUT4 #(
		.INIT('h5150)
	) name2842 (
		_w374_,
		_w2361_,
		_w2874_,
		_w2875_,
		_w2876_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2843 (
		_w486_,
		_w487_,
		_w509_,
		_w2617_,
		_w2877_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2844 (
		_w121_,
		_w418_,
		_w422_,
		_w2854_,
		_w2878_
	);
	LUT3 #(
		.INIT('h70)
	) name2845 (
		_w544_,
		_w558_,
		_w2549_,
		_w2879_
	);
	LUT3 #(
		.INIT('h01)
	) name2846 (
		_w2877_,
		_w2878_,
		_w2879_,
		_w2880_
	);
	LUT4 #(
		.INIT('h6f00)
	) name2847 (
		_w2355_,
		_w2357_,
		_w2550_,
		_w2880_,
		_w2881_
	);
	LUT2 #(
		.INIT('h6)
	) name2848 (
		\a[29] ,
		_w2881_,
		_w2882_
	);
	LUT4 #(
		.INIT('h6665)
	) name2849 (
		_w2722_,
		_w2851_,
		_w2852_,
		_w2859_,
		_w2883_
	);
	LUT4 #(
		.INIT('h90f9)
	) name2850 (
		\a[26] ,
		_w2876_,
		_w2882_,
		_w2883_,
		_w2884_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name2851 (
		_w2721_,
		_w2860_,
		_w2861_,
		_w2866_,
		_w2885_
	);
	LUT2 #(
		.INIT('h4)
	) name2852 (
		_w2884_,
		_w2885_,
		_w2886_
	);
	LUT2 #(
		.INIT('h9)
	) name2853 (
		_w2853_,
		_w2859_,
		_w2887_
	);
	LUT3 #(
		.INIT('ha9)
	) name2854 (
		_w2755_,
		_w2837_,
		_w2844_,
		_w2888_
	);
	LUT3 #(
		.INIT('h2a)
	) name2855 (
		_w376_,
		_w763_,
		_w983_,
		_w2889_
	);
	LUT3 #(
		.INIT('h70)
	) name2856 (
		_w871_,
		_w927_,
		_w2407_,
		_w2890_
	);
	LUT3 #(
		.INIT('h70)
	) name2857 (
		_w801_,
		_w851_,
		_w2527_,
		_w2891_
	);
	LUT3 #(
		.INIT('h01)
	) name2858 (
		_w2890_,
		_w2891_,
		_w2889_,
		_w2892_
	);
	LUT4 #(
		.INIT('h7d00)
	) name2859 (
		_w377_,
		_w2343_,
		_w2345_,
		_w2892_,
		_w2893_
	);
	LUT4 #(
		.INIT('h00a9)
	) name2860 (
		_w2755_,
		_w2837_,
		_w2844_,
		_w2893_,
		_w2894_
	);
	LUT4 #(
		.INIT('h153f)
	) name2861 (
		_w56_,
		_w50_,
		_w176_,
		_w378_,
		_w2895_
	);
	LUT3 #(
		.INIT('h40)
	) name2862 (
		_w53_,
		_w1510_,
		_w2895_,
		_w2896_
	);
	LUT4 #(
		.INIT('h8000)
	) name2863 (
		_w772_,
		_w933_,
		_w1184_,
		_w1257_,
		_w2897_
	);
	LUT3 #(
		.INIT('h20)
	) name2864 (
		_w126_,
		_w86_,
		_w1373_,
		_w2898_
	);
	LUT3 #(
		.INIT('h40)
	) name2865 (
		_w74_,
		_w1334_,
		_w1359_,
		_w2899_
	);
	LUT4 #(
		.INIT('h8000)
	) name2866 (
		_w2896_,
		_w2898_,
		_w2899_,
		_w2897_,
		_w2900_
	);
	LUT4 #(
		.INIT('h135f)
	) name2867 (
		_w38_,
		_w85_,
		_w259_,
		_w378_,
		_w2901_
	);
	LUT2 #(
		.INIT('h4)
	) name2868 (
		_w457_,
		_w2901_,
		_w2902_
	);
	LUT4 #(
		.INIT('h0777)
	) name2869 (
		_w122_,
		_w56_,
		_w50_,
		_w236_,
		_w2903_
	);
	LUT4 #(
		.INIT('h135f)
	) name2870 (
		_w38_,
		_w55_,
		_w201_,
		_w166_,
		_w2904_
	);
	LUT3 #(
		.INIT('h80)
	) name2871 (
		_w2282_,
		_w2903_,
		_w2904_,
		_w2905_
	);
	LUT4 #(
		.INIT('h135f)
	) name2872 (
		_w106_,
		_w41_,
		_w93_,
		_w259_,
		_w2906_
	);
	LUT4 #(
		.INIT('h135f)
	) name2873 (
		_w106_,
		_w59_,
		_w50_,
		_w419_,
		_w2907_
	);
	LUT4 #(
		.INIT('h8000)
	) name2874 (
		_w116_,
		_w659_,
		_w2906_,
		_w2907_,
		_w2908_
	);
	LUT4 #(
		.INIT('h8000)
	) name2875 (
		_w879_,
		_w2902_,
		_w2905_,
		_w2908_,
		_w2909_
	);
	LUT2 #(
		.INIT('h8)
	) name2876 (
		_w2900_,
		_w2909_,
		_w2910_
	);
	LUT4 #(
		.INIT('h0777)
	) name2877 (
		_w106_,
		_w90_,
		_w65_,
		_w378_,
		_w2911_
	);
	LUT2 #(
		.INIT('h4)
	) name2878 (
		_w439_,
		_w2911_,
		_w2912_
	);
	LUT4 #(
		.INIT('h153f)
	) name2879 (
		_w52_,
		_w110_,
		_w184_,
		_w166_,
		_w2913_
	);
	LUT4 #(
		.INIT('h153f)
	) name2880 (
		_w90_,
		_w39_,
		_w46_,
		_w236_,
		_w2914_
	);
	LUT3 #(
		.INIT('h80)
	) name2881 (
		_w1166_,
		_w2913_,
		_w2914_,
		_w2915_
	);
	LUT2 #(
		.INIT('h8)
	) name2882 (
		_w2912_,
		_w2915_,
		_w2916_
	);
	LUT4 #(
		.INIT('h135f)
	) name2883 (
		_w90_,
		_w41_,
		_w43_,
		_w176_,
		_w2917_
	);
	LUT4 #(
		.INIT('h4000)
	) name2884 (
		_w410_,
		_w834_,
		_w835_,
		_w2917_,
		_w2918_
	);
	LUT4 #(
		.INIT('h4000)
	) name2885 (
		_w369_,
		_w997_,
		_w1438_,
		_w2422_,
		_w2919_
	);
	LUT4 #(
		.INIT('h153f)
	) name2886 (
		_w38_,
		_w122_,
		_w55_,
		_w43_,
		_w2920_
	);
	LUT4 #(
		.INIT('h153f)
	) name2887 (
		_w38_,
		_w47_,
		_w158_,
		_w419_,
		_w2921_
	);
	LUT4 #(
		.INIT('h8000)
	) name2888 (
		_w81_,
		_w1226_,
		_w2920_,
		_w2921_,
		_w2922_
	);
	LUT4 #(
		.INIT('h8000)
	) name2889 (
		_w95_,
		_w514_,
		_w1012_,
		_w1576_,
		_w2923_
	);
	LUT4 #(
		.INIT('h8000)
	) name2890 (
		_w2922_,
		_w2923_,
		_w2918_,
		_w2919_,
		_w2924_
	);
	LUT4 #(
		.INIT('h135f)
	) name2891 (
		_w90_,
		_w65_,
		_w201_,
		_w259_,
		_w2925_
	);
	LUT2 #(
		.INIT('h4)
	) name2892 (
		_w450_,
		_w2925_,
		_w2926_
	);
	LUT4 #(
		.INIT('h4000)
	) name2893 (
		_w276_,
		_w597_,
		_w598_,
		_w1337_,
		_w2927_
	);
	LUT4 #(
		.INIT('h135f)
	) name2894 (
		_w55_,
		_w59_,
		_w184_,
		_w166_,
		_w2928_
	);
	LUT4 #(
		.INIT('h135f)
	) name2895 (
		_w50_,
		_w46_,
		_w201_,
		_w158_,
		_w2929_
	);
	LUT4 #(
		.INIT('h8000)
	) name2896 (
		_w806_,
		_w1790_,
		_w2929_,
		_w2928_,
		_w2930_
	);
	LUT4 #(
		.INIT('h8000)
	) name2897 (
		_w1801_,
		_w2926_,
		_w2930_,
		_w2927_,
		_w2931_
	);
	LUT4 #(
		.INIT('h8000)
	) name2898 (
		_w540_,
		_w1020_,
		_w1957_,
		_w1958_,
		_w2932_
	);
	LUT4 #(
		.INIT('h8000)
	) name2899 (
		_w2916_,
		_w2924_,
		_w2931_,
		_w2932_,
		_w2933_
	);
	LUT4 #(
		.INIT('h0888)
	) name2900 (
		_w2763_,
		_w2786_,
		_w2910_,
		_w2933_,
		_w2934_
	);
	LUT4 #(
		.INIT('h8777)
	) name2901 (
		_w2763_,
		_w2786_,
		_w2910_,
		_w2933_,
		_w2935_
	);
	LUT4 #(
		.INIT('h54ab)
	) name2902 (
		_w1189_,
		_w2335_,
		_w2336_,
		_w2338_,
		_w2936_
	);
	LUT3 #(
		.INIT('h2a)
	) name2903 (
		_w376_,
		_w1136_,
		_w1187_,
		_w2937_
	);
	LUT3 #(
		.INIT('h70)
	) name2904 (
		_w1009_,
		_w1050_,
		_w2527_,
		_w2938_
	);
	LUT3 #(
		.INIT('h70)
	) name2905 (
		_w1071_,
		_w1102_,
		_w2407_,
		_w2939_
	);
	LUT3 #(
		.INIT('h01)
	) name2906 (
		_w2938_,
		_w2939_,
		_w2937_,
		_w2940_
	);
	LUT4 #(
		.INIT('h80cc)
	) name2907 (
		_w377_,
		_w2935_,
		_w2936_,
		_w2940_,
		_w2941_
	);
	LUT3 #(
		.INIT('ha9)
	) name2908 (
		\a[20] ,
		_w2835_,
		_w2836_,
		_w2942_
	);
	LUT3 #(
		.INIT('h2a)
	) name2909 (
		_w376_,
		_w1071_,
		_w1102_,
		_w2943_
	);
	LUT3 #(
		.INIT('h70)
	) name2910 (
		_w763_,
		_w983_,
		_w2527_,
		_w2944_
	);
	LUT3 #(
		.INIT('h70)
	) name2911 (
		_w1009_,
		_w1050_,
		_w2407_,
		_w2945_
	);
	LUT3 #(
		.INIT('h01)
	) name2912 (
		_w2944_,
		_w2945_,
		_w2943_,
		_w2946_
	);
	LUT4 #(
		.INIT('h7d00)
	) name2913 (
		_w377_,
		_w2339_,
		_w2341_,
		_w2946_,
		_w2947_
	);
	LUT4 #(
		.INIT('hf110)
	) name2914 (
		_w2934_,
		_w2941_,
		_w2942_,
		_w2947_,
		_w2948_
	);
	LUT4 #(
		.INIT('h3c39)
	) name2915 (
		\a[20] ,
		_w2753_,
		_w2835_,
		_w2836_,
		_w2949_
	);
	LUT4 #(
		.INIT('h708f)
	) name2916 (
		_w377_,
		_w2839_,
		_w2843_,
		_w2949_,
		_w2950_
	);
	LUT2 #(
		.INIT('h4)
	) name2917 (
		_w2948_,
		_w2950_,
		_w2951_
	);
	LUT2 #(
		.INIT('h2)
	) name2918 (
		_w2948_,
		_w2950_,
		_w2952_
	);
	LUT2 #(
		.INIT('h9)
	) name2919 (
		_w2948_,
		_w2950_,
		_w2953_
	);
	LUT3 #(
		.INIT('h70)
	) name2920 (
		_w725_,
		_w764_,
		_w2617_,
		_w2954_
	);
	LUT3 #(
		.INIT('h70)
	) name2921 (
		_w801_,
		_w851_,
		_w2549_,
		_w2955_
	);
	LUT3 #(
		.INIT('h70)
	) name2922 (
		_w666_,
		_w694_,
		_w2854_,
		_w2956_
	);
	LUT3 #(
		.INIT('h01)
	) name2923 (
		_w2955_,
		_w2956_,
		_w2954_,
		_w2957_
	);
	LUT4 #(
		.INIT('h6f00)
	) name2924 (
		_w2347_,
		_w2349_,
		_w2550_,
		_w2957_,
		_w2958_
	);
	LUT4 #(
		.INIT('h3132)
	) name2925 (
		\a[29] ,
		_w2951_,
		_w2952_,
		_w2958_,
		_w2959_
	);
	LUT4 #(
		.INIT('h5600)
	) name2926 (
		_w2755_,
		_w2837_,
		_w2844_,
		_w2893_,
		_w2960_
	);
	LUT4 #(
		.INIT('ha956)
	) name2927 (
		_w2755_,
		_w2837_,
		_w2844_,
		_w2893_,
		_w2961_
	);
	LUT2 #(
		.INIT('h9)
	) name2928 (
		_w2845_,
		_w2847_,
		_w2962_
	);
	LUT4 #(
		.INIT('h00d4)
	) name2929 (
		_w2888_,
		_w2893_,
		_w2959_,
		_w2962_,
		_w2963_
	);
	LUT4 #(
		.INIT('h2b00)
	) name2930 (
		_w2888_,
		_w2893_,
		_w2959_,
		_w2962_,
		_w2964_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2931 (
		_w587_,
		_w608_,
		_w624_,
		_w2617_,
		_w2965_
	);
	LUT3 #(
		.INIT('h70)
	) name2932 (
		_w666_,
		_w694_,
		_w2549_,
		_w2966_
	);
	LUT3 #(
		.INIT('h70)
	) name2933 (
		_w544_,
		_w558_,
		_w2854_,
		_w2967_
	);
	LUT3 #(
		.INIT('h01)
	) name2934 (
		_w2966_,
		_w2967_,
		_w2965_,
		_w2968_
	);
	LUT4 #(
		.INIT('h6f00)
	) name2935 (
		_w2351_,
		_w2353_,
		_w2550_,
		_w2968_,
		_w2969_
	);
	LUT2 #(
		.INIT('h6)
	) name2936 (
		\a[29] ,
		_w2969_,
		_w2970_
	);
	LUT3 #(
		.INIT('h45)
	) name2937 (
		_w2963_,
		_w2964_,
		_w2970_,
		_w2971_
	);
	LUT2 #(
		.INIT('h8)
	) name2938 (
		_w2887_,
		_w2971_,
		_w2972_
	);
	LUT4 #(
		.INIT('hf400)
	) name2939 (
		_w374_,
		_w2361_,
		_w2404_,
		_w2875_,
		_w2973_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2940 (
		_w121_,
		_w418_,
		_w422_,
		_w2874_,
		_w2974_
	);
	LUT3 #(
		.INIT('h18)
	) name2941 (
		\a[23] ,
		\a[24] ,
		\a[25] ,
		_w2975_
	);
	LUT3 #(
		.INIT('h70)
	) name2942 (
		_w352_,
		_w373_,
		_w2975_,
		_w2976_
	);
	LUT2 #(
		.INIT('h1)
	) name2943 (
		_w2974_,
		_w2976_,
		_w2977_
	);
	LUT3 #(
		.INIT('h9a)
	) name2944 (
		\a[26] ,
		_w2973_,
		_w2977_,
		_w2978_
	);
	LUT2 #(
		.INIT('h1)
	) name2945 (
		_w2887_,
		_w2971_,
		_w2979_
	);
	LUT2 #(
		.INIT('h6)
	) name2946 (
		_w2887_,
		_w2971_,
		_w2980_
	);
	LUT3 #(
		.INIT('h54)
	) name2947 (
		_w2972_,
		_w2978_,
		_w2979_,
		_w2981_
	);
	LUT4 #(
		.INIT('h9669)
	) name2948 (
		\a[26] ,
		_w2876_,
		_w2882_,
		_w2883_,
		_w2982_
	);
	LUT4 #(
		.INIT('h8e00)
	) name2949 (
		_w2887_,
		_w2971_,
		_w2978_,
		_w2982_,
		_w2983_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2950 (
		_w486_,
		_w487_,
		_w509_,
		_w2874_,
		_w2984_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2951 (
		_w121_,
		_w418_,
		_w422_,
		_w2975_,
		_w2985_
	);
	LUT4 #(
		.INIT('h6006)
	) name2952 (
		\a[23] ,
		\a[24] ,
		\a[25] ,
		\a[26] ,
		_w2986_
	);
	LUT3 #(
		.INIT('h70)
	) name2953 (
		_w352_,
		_w373_,
		_w2986_,
		_w2987_
	);
	LUT3 #(
		.INIT('h01)
	) name2954 (
		_w2984_,
		_w2985_,
		_w2987_,
		_w2988_
	);
	LUT4 #(
		.INIT('h95aa)
	) name2955 (
		\a[26] ,
		_w2535_,
		_w2875_,
		_w2988_,
		_w2989_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2956 (
		_w587_,
		_w608_,
		_w624_,
		_w2854_,
		_w2990_
	);
	LUT3 #(
		.INIT('h70)
	) name2957 (
		_w725_,
		_w764_,
		_w2549_,
		_w2991_
	);
	LUT3 #(
		.INIT('h70)
	) name2958 (
		_w666_,
		_w694_,
		_w2617_,
		_w2992_
	);
	LUT3 #(
		.INIT('h01)
	) name2959 (
		_w2991_,
		_w2992_,
		_w2990_,
		_w2993_
	);
	LUT4 #(
		.INIT('h95aa)
	) name2960 (
		\a[29] ,
		_w2550_,
		_w2598_,
		_w2993_,
		_w2994_
	);
	LUT3 #(
		.INIT('h60)
	) name2961 (
		_w2959_,
		_w2961_,
		_w2994_,
		_w2995_
	);
	LUT3 #(
		.INIT('h09)
	) name2962 (
		_w2959_,
		_w2961_,
		_w2994_,
		_w2996_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2963 (
		_w486_,
		_w487_,
		_w509_,
		_w2975_,
		_w2997_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2964 (
		_w121_,
		_w418_,
		_w422_,
		_w2986_,
		_w2998_
	);
	LUT3 #(
		.INIT('h70)
	) name2965 (
		_w544_,
		_w558_,
		_w2874_,
		_w2999_
	);
	LUT3 #(
		.INIT('h01)
	) name2966 (
		_w2997_,
		_w2998_,
		_w2999_,
		_w3000_
	);
	LUT4 #(
		.INIT('h6f00)
	) name2967 (
		_w2355_,
		_w2357_,
		_w2875_,
		_w3000_,
		_w3001_
	);
	LUT4 #(
		.INIT('h3231)
	) name2968 (
		\a[26] ,
		_w2995_,
		_w2996_,
		_w3001_,
		_w3002_
	);
	LUT4 #(
		.INIT('h54ab)
	) name2969 (
		_w2894_,
		_w2959_,
		_w2960_,
		_w2962_,
		_w3003_
	);
	LUT2 #(
		.INIT('h6)
	) name2970 (
		_w2970_,
		_w3003_,
		_w3004_
	);
	LUT3 #(
		.INIT('hb2)
	) name2971 (
		_w2989_,
		_w3002_,
		_w3004_,
		_w3005_
	);
	LUT2 #(
		.INIT('h9)
	) name2972 (
		_w2978_,
		_w2980_,
		_w3006_
	);
	LUT3 #(
		.INIT('h09)
	) name2973 (
		_w2978_,
		_w2980_,
		_w3005_,
		_w3007_
	);
	LUT3 #(
		.INIT('h96)
	) name2974 (
		_w2989_,
		_w3002_,
		_w3004_,
		_w3008_
	);
	LUT3 #(
		.INIT('h70)
	) name2975 (
		_w725_,
		_w764_,
		_w2854_,
		_w3009_
	);
	LUT3 #(
		.INIT('h70)
	) name2976 (
		_w801_,
		_w851_,
		_w2617_,
		_w3010_
	);
	LUT3 #(
		.INIT('h70)
	) name2977 (
		_w871_,
		_w927_,
		_w2549_,
		_w3011_
	);
	LUT3 #(
		.INIT('h01)
	) name2978 (
		_w3010_,
		_w3011_,
		_w3009_,
		_w3012_
	);
	LUT4 #(
		.INIT('h95aa)
	) name2979 (
		\a[29] ,
		_w2550_,
		_w2724_,
		_w3012_,
		_w3013_
	);
	LUT4 #(
		.INIT('he11e)
	) name2980 (
		_w2934_,
		_w2941_,
		_w2942_,
		_w2947_,
		_w3014_
	);
	LUT4 #(
		.INIT('h6c33)
	) name2981 (
		_w377_,
		_w2935_,
		_w2936_,
		_w2940_,
		_w3015_
	);
	LUT4 #(
		.INIT('h8000)
	) name2982 (
		_w391_,
		_w816_,
		_w980_,
		_w1012_,
		_w3016_
	);
	LUT4 #(
		.INIT('h135f)
	) name2983 (
		_w52_,
		_w67_,
		_w201_,
		_w236_,
		_w3017_
	);
	LUT2 #(
		.INIT('h8)
	) name2984 (
		_w1953_,
		_w3017_,
		_w3018_
	);
	LUT4 #(
		.INIT('h135f)
	) name2985 (
		_w110_,
		_w47_,
		_w43_,
		_w184_,
		_w3019_
	);
	LUT4 #(
		.INIT('h153f)
	) name2986 (
		_w47_,
		_w46_,
		_w166_,
		_w259_,
		_w3020_
	);
	LUT4 #(
		.INIT('h8000)
	) name2987 (
		_w1953_,
		_w3017_,
		_w3019_,
		_w3020_,
		_w3021_
	);
	LUT4 #(
		.INIT('h153f)
	) name2988 (
		_w67_,
		_w50_,
		_w201_,
		_w158_,
		_w3022_
	);
	LUT4 #(
		.INIT('h8000)
	) name2989 (
		_w1216_,
		_w1374_,
		_w1978_,
		_w3022_,
		_w3023_
	);
	LUT4 #(
		.INIT('h8000)
	) name2990 (
		_w891_,
		_w3023_,
		_w3016_,
		_w3021_,
		_w3024_
	);
	LUT4 #(
		.INIT('h8000)
	) name2991 (
		_w526_,
		_w1995_,
		_w2110_,
		_w3024_,
		_w3025_
	);
	LUT2 #(
		.INIT('h8)
	) name2992 (
		_w648_,
		_w3025_,
		_w3026_
	);
	LUT4 #(
		.INIT('h153f)
	) name2993 (
		_w110_,
		_w50_,
		_w201_,
		_w430_,
		_w3027_
	);
	LUT4 #(
		.INIT('h8000)
	) name2994 (
		_w584_,
		_w629_,
		_w670_,
		_w3027_,
		_w3028_
	);
	LUT4 #(
		.INIT('h135f)
	) name2995 (
		_w38_,
		_w59_,
		_w184_,
		_w158_,
		_w3029_
	);
	LUT4 #(
		.INIT('h4000)
	) name2996 (
		_w454_,
		_w662_,
		_w643_,
		_w3029_,
		_w3030_
	);
	LUT2 #(
		.INIT('h8)
	) name2997 (
		_w3028_,
		_w3030_,
		_w3031_
	);
	LUT4 #(
		.INIT('h8000)
	) name2998 (
		_w1138_,
		_w1649_,
		_w1682_,
		_w2913_,
		_w3032_
	);
	LUT4 #(
		.INIT('h135f)
	) name2999 (
		_w106_,
		_w52_,
		_w46_,
		_w236_,
		_w3033_
	);
	LUT3 #(
		.INIT('h80)
	) name3000 (
		_w1362_,
		_w1761_,
		_w3033_,
		_w3034_
	);
	LUT4 #(
		.INIT('h0777)
	) name3001 (
		_w78_,
		_w93_,
		_w65_,
		_w176_,
		_w3035_
	);
	LUT4 #(
		.INIT('h153f)
	) name3002 (
		_w59_,
		_w56_,
		_w259_,
		_w176_,
		_w3036_
	);
	LUT4 #(
		.INIT('h153f)
	) name3003 (
		_w67_,
		_w41_,
		_w72_,
		_w158_,
		_w3037_
	);
	LUT4 #(
		.INIT('h8000)
	) name3004 (
		_w1341_,
		_w3037_,
		_w3035_,
		_w3036_,
		_w3038_
	);
	LUT4 #(
		.INIT('h8000)
	) name3005 (
		_w1424_,
		_w3034_,
		_w3038_,
		_w3032_,
		_w3039_
	);
	LUT4 #(
		.INIT('h0777)
	) name3006 (
		_w50_,
		_w43_,
		_w46_,
		_w158_,
		_w3040_
	);
	LUT4 #(
		.INIT('h153f)
	) name3007 (
		_w56_,
		_w93_,
		_w378_,
		_w430_,
		_w3041_
	);
	LUT4 #(
		.INIT('h4000)
	) name3008 (
		_w186_,
		_w971_,
		_w3040_,
		_w3041_,
		_w3042_
	);
	LUT3 #(
		.INIT('h1f)
	) name3009 (
		_w85_,
		_w93_,
		_w176_,
		_w3043_
	);
	LUT2 #(
		.INIT('h8)
	) name3010 (
		_w966_,
		_w3043_,
		_w3044_
	);
	LUT4 #(
		.INIT('h0777)
	) name3011 (
		_w67_,
		_w72_,
		_w50_,
		_w419_,
		_w3045_
	);
	LUT2 #(
		.INIT('h8)
	) name3012 (
		_w899_,
		_w3045_,
		_w3046_
	);
	LUT4 #(
		.INIT('h8000)
	) name3013 (
		_w899_,
		_w966_,
		_w3043_,
		_w3045_,
		_w3047_
	);
	LUT2 #(
		.INIT('h8)
	) name3014 (
		_w3042_,
		_w3047_,
		_w3048_
	);
	LUT3 #(
		.INIT('h80)
	) name3015 (
		_w1580_,
		_w1634_,
		_w2015_,
		_w3049_
	);
	LUT4 #(
		.INIT('h8000)
	) name3016 (
		_w370_,
		_w1184_,
		_w1278_,
		_w1510_,
		_w3050_
	);
	LUT3 #(
		.INIT('h80)
	) name3017 (
		_w242_,
		_w3049_,
		_w3050_,
		_w3051_
	);
	LUT4 #(
		.INIT('h8000)
	) name3018 (
		_w3031_,
		_w3039_,
		_w3048_,
		_w3051_,
		_w3052_
	);
	LUT2 #(
		.INIT('h8)
	) name3019 (
		_w801_,
		_w3052_,
		_w3053_
	);
	LUT4 #(
		.INIT('h135f)
	) name3020 (
		_w648_,
		_w801_,
		_w3025_,
		_w3052_,
		_w3054_
	);
	LUT4 #(
		.INIT('h8000)
	) name3021 (
		_w648_,
		_w801_,
		_w3025_,
		_w3052_,
		_w3055_
	);
	LUT4 #(
		.INIT('h044c)
	) name3022 (
		\a[17] ,
		_w2787_,
		_w3026_,
		_w3053_,
		_w3056_
	);
	LUT4 #(
		.INIT('h3220)
	) name3023 (
		\a[17] ,
		_w2787_,
		_w3026_,
		_w3053_,
		_w3057_
	);
	LUT3 #(
		.INIT('h70)
	) name3024 (
		_w1136_,
		_w1187_,
		_w2407_,
		_w3058_
	);
	LUT3 #(
		.INIT('h70)
	) name3025 (
		_w1071_,
		_w1102_,
		_w2527_,
		_w3059_
	);
	LUT3 #(
		.INIT('h2a)
	) name3026 (
		_w376_,
		_w1202_,
		_w1233_,
		_w3060_
	);
	LUT3 #(
		.INIT('h01)
	) name3027 (
		_w3059_,
		_w3060_,
		_w3058_,
		_w3061_
	);
	LUT4 #(
		.INIT('h7d00)
	) name3028 (
		_w377_,
		_w2335_,
		_w2337_,
		_w3061_,
		_w3062_
	);
	LUT3 #(
		.INIT('h54)
	) name3029 (
		_w3056_,
		_w3057_,
		_w3062_,
		_w3063_
	);
	LUT2 #(
		.INIT('h2)
	) name3030 (
		_w3015_,
		_w3063_,
		_w3064_
	);
	LUT2 #(
		.INIT('h9)
	) name3031 (
		_w3015_,
		_w3063_,
		_w3065_
	);
	LUT3 #(
		.INIT('ha9)
	) name3032 (
		\a[17] ,
		_w3054_,
		_w3055_,
		_w3066_
	);
	LUT4 #(
		.INIT('h54ab)
	) name3033 (
		_w1296_,
		_w2331_,
		_w2332_,
		_w2334_,
		_w3067_
	);
	LUT3 #(
		.INIT('h70)
	) name3034 (
		_w1136_,
		_w1187_,
		_w2527_,
		_w3068_
	);
	LUT3 #(
		.INIT('h70)
	) name3035 (
		_w1202_,
		_w1233_,
		_w2407_,
		_w3069_
	);
	LUT3 #(
		.INIT('h2a)
	) name3036 (
		_w376_,
		_w1253_,
		_w1294_,
		_w3070_
	);
	LUT3 #(
		.INIT('h01)
	) name3037 (
		_w3069_,
		_w3070_,
		_w3068_,
		_w3071_
	);
	LUT4 #(
		.INIT('h2033)
	) name3038 (
		_w377_,
		_w3066_,
		_w3067_,
		_w3071_,
		_w3072_
	);
	LUT4 #(
		.INIT('h0777)
	) name3039 (
		_w67_,
		_w72_,
		_w46_,
		_w158_,
		_w3073_
	);
	LUT4 #(
		.INIT('h8000)
	) name3040 (
		_w1961_,
		_w2090_,
		_w2116_,
		_w3073_,
		_w3074_
	);
	LUT3 #(
		.INIT('h80)
	) name3041 (
		_w1011_,
		_w2052_,
		_w3074_,
		_w3075_
	);
	LUT4 #(
		.INIT('h135f)
	) name3042 (
		_w106_,
		_w67_,
		_w65_,
		_w158_,
		_w3076_
	);
	LUT4 #(
		.INIT('h135f)
	) name3043 (
		_w110_,
		_w44_,
		_w158_,
		_w430_,
		_w3077_
	);
	LUT4 #(
		.INIT('h8000)
	) name3044 (
		_w1448_,
		_w1761_,
		_w3076_,
		_w3077_,
		_w3078_
	);
	LUT3 #(
		.INIT('h80)
	) name3045 (
		_w2187_,
		_w2271_,
		_w3078_,
		_w3079_
	);
	LUT2 #(
		.INIT('h4)
	) name3046 (
		_w142_,
		_w1281_,
		_w3080_
	);
	LUT3 #(
		.INIT('h80)
	) name3047 (
		_w311_,
		_w876_,
		_w1114_,
		_w3081_
	);
	LUT3 #(
		.INIT('h80)
	) name3048 (
		_w2114_,
		_w3080_,
		_w3081_,
		_w3082_
	);
	LUT3 #(
		.INIT('h57)
	) name3049 (
		_w59_,
		_w72_,
		_w259_,
		_w3083_
	);
	LUT2 #(
		.INIT('h8)
	) name3050 (
		_w2126_,
		_w3083_,
		_w3084_
	);
	LUT4 #(
		.INIT('h135f)
	) name3051 (
		_w59_,
		_w90_,
		_w166_,
		_w176_,
		_w3085_
	);
	LUT4 #(
		.INIT('h8000)
	) name3052 (
		_w367_,
		_w553_,
		_w760_,
		_w3085_,
		_w3086_
	);
	LUT4 #(
		.INIT('h153f)
	) name3053 (
		_w52_,
		_w50_,
		_w158_,
		_w378_,
		_w3087_
	);
	LUT4 #(
		.INIT('h153f)
	) name3054 (
		_w110_,
		_w67_,
		_w419_,
		_w430_,
		_w3088_
	);
	LUT4 #(
		.INIT('h8000)
	) name3055 (
		_w1108_,
		_w1181_,
		_w3087_,
		_w3088_,
		_w3089_
	);
	LUT4 #(
		.INIT('h8000)
	) name3056 (
		_w1861_,
		_w3084_,
		_w3089_,
		_w3086_,
		_w3090_
	);
	LUT4 #(
		.INIT('h8000)
	) name3057 (
		_w3082_,
		_w3090_,
		_w3075_,
		_w3079_,
		_w3091_
	);
	LUT2 #(
		.INIT('h8)
	) name3058 (
		_w2421_,
		_w3091_,
		_w3092_
	);
	LUT4 #(
		.INIT('h20a0)
	) name3059 (
		_w648_,
		_w2421_,
		_w3025_,
		_w3091_,
		_w3093_
	);
	LUT4 #(
		.INIT('h935f)
	) name3060 (
		_w648_,
		_w2421_,
		_w3025_,
		_w3091_,
		_w3094_
	);
	LUT3 #(
		.INIT('h1f)
	) name3061 (
		_w90_,
		_w50_,
		_w184_,
		_w3095_
	);
	LUT4 #(
		.INIT('h4000)
	) name3062 (
		_w169_,
		_w668_,
		_w901_,
		_w3095_,
		_w3096_
	);
	LUT4 #(
		.INIT('h1000)
	) name3063 (
		_w282_,
		_w437_,
		_w1808_,
		_w2267_,
		_w3097_
	);
	LUT2 #(
		.INIT('h8)
	) name3064 (
		_w3096_,
		_w3097_,
		_w3098_
	);
	LUT3 #(
		.INIT('h57)
	) name3065 (
		_w93_,
		_w201_,
		_w419_,
		_w3099_
	);
	LUT4 #(
		.INIT('h8000)
	) name3066 (
		_w980_,
		_w986_,
		_w2427_,
		_w3099_,
		_w3100_
	);
	LUT4 #(
		.INIT('h0777)
	) name3067 (
		_w38_,
		_w78_,
		_w44_,
		_w184_,
		_w3101_
	);
	LUT3 #(
		.INIT('h80)
	) name3068 (
		_w1066_,
		_w1288_,
		_w3101_,
		_w3102_
	);
	LUT4 #(
		.INIT('h135f)
	) name3069 (
		_w65_,
		_w46_,
		_w176_,
		_w378_,
		_w3103_
	);
	LUT3 #(
		.INIT('h80)
	) name3070 (
		_w1184_,
		_w1472_,
		_w3103_,
		_w3104_
	);
	LUT3 #(
		.INIT('h80)
	) name3071 (
		_w3102_,
		_w3100_,
		_w3104_,
		_w3105_
	);
	LUT3 #(
		.INIT('h80)
	) name3072 (
		_w3082_,
		_w3098_,
		_w3105_,
		_w3106_
	);
	LUT4 #(
		.INIT('h135f)
	) name3073 (
		_w122_,
		_w55_,
		_w85_,
		_w236_,
		_w3107_
	);
	LUT2 #(
		.INIT('h8)
	) name3074 (
		_w1434_,
		_w3107_,
		_w3108_
	);
	LUT4 #(
		.INIT('h135f)
	) name3075 (
		_w38_,
		_w85_,
		_w166_,
		_w158_,
		_w3109_
	);
	LUT2 #(
		.INIT('h4)
	) name3076 (
		_w69_,
		_w3109_,
		_w3110_
	);
	LUT4 #(
		.INIT('h1000)
	) name3077 (
		_w69_,
		_w458_,
		_w1845_,
		_w3109_,
		_w3111_
	);
	LUT2 #(
		.INIT('h8)
	) name3078 (
		_w3108_,
		_w3111_,
		_w3112_
	);
	LUT4 #(
		.INIT('h153f)
	) name3079 (
		_w110_,
		_w78_,
		_w46_,
		_w184_,
		_w3113_
	);
	LUT3 #(
		.INIT('h80)
	) name3080 (
		_w296_,
		_w1518_,
		_w3113_,
		_w3114_
	);
	LUT4 #(
		.INIT('h0777)
	) name3081 (
		_w59_,
		_w39_,
		_w50_,
		_w176_,
		_w3115_
	);
	LUT4 #(
		.INIT('h0400)
	) name3082 (
		_w273_,
		_w348_,
		_w471_,
		_w3115_,
		_w3116_
	);
	LUT4 #(
		.INIT('h8000)
	) name3083 (
		_w841_,
		_w2189_,
		_w3114_,
		_w3116_,
		_w3117_
	);
	LUT2 #(
		.INIT('h8)
	) name3084 (
		_w3112_,
		_w3117_,
		_w3118_
	);
	LUT3 #(
		.INIT('h80)
	) name3085 (
		_w1628_,
		_w2903_,
		_w2929_,
		_w3119_
	);
	LUT2 #(
		.INIT('h4)
	) name3086 (
		_w379_,
		_w554_,
		_w3120_
	);
	LUT4 #(
		.INIT('h0777)
	) name3087 (
		_w122_,
		_w52_,
		_w59_,
		_w184_,
		_w3121_
	);
	LUT4 #(
		.INIT('h153f)
	) name3088 (
		_w90_,
		_w65_,
		_w201_,
		_w259_,
		_w3122_
	);
	LUT4 #(
		.INIT('h8000)
	) name3089 (
		_w322_,
		_w770_,
		_w3121_,
		_w3122_,
		_w3123_
	);
	LUT3 #(
		.INIT('h80)
	) name3090 (
		_w3120_,
		_w3119_,
		_w3123_,
		_w3124_
	);
	LUT4 #(
		.INIT('h153f)
	) name3091 (
		_w106_,
		_w78_,
		_w47_,
		_w50_,
		_w3125_
	);
	LUT2 #(
		.INIT('h4)
	) name3092 (
		_w429_,
		_w3125_,
		_w3126_
	);
	LUT4 #(
		.INIT('h153f)
	) name3093 (
		_w55_,
		_w67_,
		_w43_,
		_w166_,
		_w3127_
	);
	LUT4 #(
		.INIT('h4000)
	) name3094 (
		_w443_,
		_w1910_,
		_w2015_,
		_w3127_,
		_w3128_
	);
	LUT2 #(
		.INIT('h8)
	) name3095 (
		_w3126_,
		_w3128_,
		_w3129_
	);
	LUT4 #(
		.INIT('h153f)
	) name3096 (
		_w56_,
		_w41_,
		_w72_,
		_w39_,
		_w3130_
	);
	LUT4 #(
		.INIT('h8000)
	) name3097 (
		_w553_,
		_w649_,
		_w670_,
		_w3130_,
		_w3131_
	);
	LUT4 #(
		.INIT('h153f)
	) name3098 (
		_w38_,
		_w67_,
		_w39_,
		_w236_,
		_w3132_
	);
	LUT4 #(
		.INIT('h1000)
	) name3099 (
		_w339_,
		_w359_,
		_w1945_,
		_w3132_,
		_w3133_
	);
	LUT4 #(
		.INIT('h135f)
	) name3100 (
		_w59_,
		_w47_,
		_w166_,
		_w158_,
		_w3134_
	);
	LUT4 #(
		.INIT('h153f)
	) name3101 (
		_w85_,
		_w67_,
		_w78_,
		_w39_,
		_w3135_
	);
	LUT3 #(
		.INIT('h80)
	) name3102 (
		_w1888_,
		_w3135_,
		_w3134_,
		_w3136_
	);
	LUT4 #(
		.INIT('h8000)
	) name3103 (
		_w2781_,
		_w3136_,
		_w3131_,
		_w3133_,
		_w3137_
	);
	LUT3 #(
		.INIT('h80)
	) name3104 (
		_w3124_,
		_w3129_,
		_w3137_,
		_w3138_
	);
	LUT3 #(
		.INIT('h80)
	) name3105 (
		_w3106_,
		_w3118_,
		_w3138_,
		_w3139_
	);
	LUT3 #(
		.INIT('h80)
	) name3106 (
		_w1993_,
		_w2257_,
		_w2510_,
		_w3140_
	);
	LUT4 #(
		.INIT('h135f)
	) name3107 (
		_w90_,
		_w41_,
		_w201_,
		_w236_,
		_w3141_
	);
	LUT4 #(
		.INIT('h2000)
	) name3108 (
		_w309_,
		_w481_,
		_w1215_,
		_w3141_,
		_w3142_
	);
	LUT3 #(
		.INIT('h80)
	) name3109 (
		_w3044_,
		_w3140_,
		_w3142_,
		_w3143_
	);
	LUT3 #(
		.INIT('h57)
	) name3110 (
		_w56_,
		_w236_,
		_w259_,
		_w3144_
	);
	LUT3 #(
		.INIT('h80)
	) name3111 (
		_w1414_,
		_w1603_,
		_w3144_,
		_w3145_
	);
	LUT4 #(
		.INIT('h0777)
	) name3112 (
		_w106_,
		_w47_,
		_w50_,
		_w184_,
		_w3146_
	);
	LUT4 #(
		.INIT('h135f)
	) name3113 (
		_w55_,
		_w44_,
		_w259_,
		_w430_,
		_w3147_
	);
	LUT4 #(
		.INIT('h153f)
	) name3114 (
		_w72_,
		_w50_,
		_w43_,
		_w65_,
		_w3148_
	);
	LUT4 #(
		.INIT('h8000)
	) name3115 (
		_w990_,
		_w3148_,
		_w3146_,
		_w3147_,
		_w3149_
	);
	LUT3 #(
		.INIT('h80)
	) name3116 (
		_w3084_,
		_w3145_,
		_w3149_,
		_w3150_
	);
	LUT3 #(
		.INIT('h80)
	) name3117 (
		_w692_,
		_w3143_,
		_w3150_,
		_w3151_
	);
	LUT4 #(
		.INIT('h153f)
	) name3118 (
		_w38_,
		_w56_,
		_w184_,
		_w201_,
		_w3152_
	);
	LUT4 #(
		.INIT('h153f)
	) name3119 (
		_w38_,
		_w90_,
		_w419_,
		_w378_,
		_w3153_
	);
	LUT2 #(
		.INIT('h8)
	) name3120 (
		_w3152_,
		_w3153_,
		_w3154_
	);
	LUT4 #(
		.INIT('h0777)
	) name3121 (
		_w78_,
		_w56_,
		_w50_,
		_w201_,
		_w3155_
	);
	LUT4 #(
		.INIT('h8000)
	) name3122 (
		_w305_,
		_w408_,
		_w809_,
		_w3155_,
		_w3156_
	);
	LUT2 #(
		.INIT('h8)
	) name3123 (
		_w3154_,
		_w3156_,
		_w3157_
	);
	LUT4 #(
		.INIT('h0777)
	) name3124 (
		_w41_,
		_w43_,
		_w46_,
		_w236_,
		_w3158_
	);
	LUT3 #(
		.INIT('h80)
	) name3125 (
		_w1174_,
		_w1736_,
		_w3158_,
		_w3159_
	);
	LUT3 #(
		.INIT('h02)
	) name3126 (
		_w115_,
		_w77_,
		_w476_,
		_w3160_
	);
	LUT4 #(
		.INIT('h8000)
	) name3127 (
		_w2028_,
		_w2922_,
		_w3160_,
		_w3159_,
		_w3161_
	);
	LUT2 #(
		.INIT('h8)
	) name3128 (
		_w3157_,
		_w3161_,
		_w3162_
	);
	LUT4 #(
		.INIT('h153f)
	) name3129 (
		_w122_,
		_w78_,
		_w90_,
		_w65_,
		_w3163_
	);
	LUT4 #(
		.INIT('h4000)
	) name3130 (
		_w214_,
		_w1206_,
		_w1278_,
		_w3163_,
		_w3164_
	);
	LUT3 #(
		.INIT('h57)
	) name3131 (
		_w50_,
		_w166_,
		_w378_,
		_w3165_
	);
	LUT2 #(
		.INIT('h4)
	) name3132 (
		_w452_,
		_w3165_,
		_w3166_
	);
	LUT4 #(
		.INIT('h4000)
	) name3133 (
		_w346_,
		_w1350_,
		_w1351_,
		_w2046_,
		_w3167_
	);
	LUT3 #(
		.INIT('h80)
	) name3134 (
		_w3166_,
		_w3164_,
		_w3167_,
		_w3168_
	);
	LUT4 #(
		.INIT('h0777)
	) name3135 (
		_w106_,
		_w55_,
		_w90_,
		_w236_,
		_w3169_
	);
	LUT3 #(
		.INIT('h40)
	) name3136 (
		_w396_,
		_w1055_,
		_w3169_,
		_w3170_
	);
	LUT2 #(
		.INIT('h8)
	) name3137 (
		_w1670_,
		_w3170_,
		_w3171_
	);
	LUT2 #(
		.INIT('h8)
	) name3138 (
		_w1180_,
		_w1475_,
		_w3172_
	);
	LUT4 #(
		.INIT('h4000)
	) name3139 (
		_w203_,
		_w538_,
		_w663_,
		_w1245_,
		_w3173_
	);
	LUT3 #(
		.INIT('h80)
	) name3140 (
		_w704_,
		_w957_,
		_w2274_,
		_w3174_
	);
	LUT4 #(
		.INIT('h153f)
	) name3141 (
		_w56_,
		_w41_,
		_w259_,
		_w430_,
		_w3175_
	);
	LUT4 #(
		.INIT('h0800)
	) name3142 (
		_w139_,
		_w274_,
		_w444_,
		_w3175_,
		_w3176_
	);
	LUT4 #(
		.INIT('h8000)
	) name3143 (
		_w3172_,
		_w3174_,
		_w3176_,
		_w3173_,
		_w3177_
	);
	LUT3 #(
		.INIT('h80)
	) name3144 (
		_w3168_,
		_w3171_,
		_w3177_,
		_w3178_
	);
	LUT3 #(
		.INIT('h80)
	) name3145 (
		_w3162_,
		_w3151_,
		_w3178_,
		_w3179_
	);
	LUT4 #(
		.INIT('h044c)
	) name3146 (
		\a[14] ,
		_w3092_,
		_w3139_,
		_w3179_,
		_w3180_
	);
	LUT4 #(
		.INIT('h3220)
	) name3147 (
		\a[14] ,
		_w3092_,
		_w3139_,
		_w3179_,
		_w3181_
	);
	LUT4 #(
		.INIT('h54ab)
	) name3148 (
		_w1400_,
		_w2327_,
		_w2328_,
		_w2330_,
		_w3182_
	);
	LUT3 #(
		.INIT('h2a)
	) name3149 (
		_w376_,
		_w1381_,
		_w1398_,
		_w3183_
	);
	LUT3 #(
		.INIT('h70)
	) name3150 (
		_w1325_,
		_w1367_,
		_w2407_,
		_w3184_
	);
	LUT3 #(
		.INIT('h70)
	) name3151 (
		_w1253_,
		_w1294_,
		_w2527_,
		_w3185_
	);
	LUT3 #(
		.INIT('h01)
	) name3152 (
		_w3184_,
		_w3185_,
		_w3183_,
		_w3186_
	);
	LUT4 #(
		.INIT('h2033)
	) name3153 (
		_w377_,
		_w3181_,
		_w3182_,
		_w3186_,
		_w3187_
	);
	LUT4 #(
		.INIT('h1115)
	) name3154 (
		_w3093_,
		_w3094_,
		_w3180_,
		_w3187_,
		_w3188_
	);
	LUT4 #(
		.INIT('h4c00)
	) name3155 (
		_w377_,
		_w3066_,
		_w3067_,
		_w3071_,
		_w3189_
	);
	LUT4 #(
		.INIT('h93cc)
	) name3156 (
		_w377_,
		_w3066_,
		_w3067_,
		_w3071_,
		_w3190_
	);
	LUT3 #(
		.INIT('h54)
	) name3157 (
		_w3072_,
		_w3188_,
		_w3189_,
		_w3191_
	);
	LUT4 #(
		.INIT('h3c39)
	) name3158 (
		\a[17] ,
		_w2787_,
		_w3054_,
		_w3055_,
		_w3192_
	);
	LUT2 #(
		.INIT('h9)
	) name3159 (
		_w3062_,
		_w3192_,
		_w3193_
	);
	LUT2 #(
		.INIT('h4)
	) name3160 (
		_w3191_,
		_w3193_,
		_w3194_
	);
	LUT2 #(
		.INIT('h2)
	) name3161 (
		_w3191_,
		_w3193_,
		_w3195_
	);
	LUT2 #(
		.INIT('h9)
	) name3162 (
		_w3191_,
		_w3193_,
		_w3196_
	);
	LUT3 #(
		.INIT('h70)
	) name3163 (
		_w1009_,
		_w1050_,
		_w2549_,
		_w3197_
	);
	LUT3 #(
		.INIT('h70)
	) name3164 (
		_w871_,
		_w927_,
		_w2854_,
		_w3198_
	);
	LUT3 #(
		.INIT('h70)
	) name3165 (
		_w763_,
		_w983_,
		_w2617_,
		_w3199_
	);
	LUT3 #(
		.INIT('h01)
	) name3166 (
		_w3198_,
		_w3199_,
		_w3197_,
		_w3200_
	);
	LUT4 #(
		.INIT('h95aa)
	) name3167 (
		\a[29] ,
		_w2550_,
		_w2839_,
		_w3200_,
		_w3201_
	);
	LUT4 #(
		.INIT('h20a2)
	) name3168 (
		_w3065_,
		_w3191_,
		_w3193_,
		_w3201_,
		_w3202_
	);
	LUT4 #(
		.INIT('h222b)
	) name3169 (
		_w3013_,
		_w3014_,
		_w3064_,
		_w3202_,
		_w3203_
	);
	LUT3 #(
		.INIT('h69)
	) name3170 (
		\a[29] ,
		_w2953_,
		_w2958_,
		_w3204_
	);
	LUT2 #(
		.INIT('h4)
	) name3171 (
		_w3203_,
		_w3204_,
		_w3205_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3172 (
		_w486_,
		_w487_,
		_w509_,
		_w2986_,
		_w3206_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3173 (
		_w587_,
		_w608_,
		_w624_,
		_w2874_,
		_w3207_
	);
	LUT3 #(
		.INIT('h70)
	) name3174 (
		_w544_,
		_w558_,
		_w2975_,
		_w3208_
	);
	LUT3 #(
		.INIT('h01)
	) name3175 (
		_w3206_,
		_w3207_,
		_w3208_,
		_w3209_
	);
	LUT4 #(
		.INIT('h95aa)
	) name3176 (
		\a[26] ,
		_w2526_,
		_w2875_,
		_w3209_,
		_w3210_
	);
	LUT2 #(
		.INIT('h2)
	) name3177 (
		_w3203_,
		_w3204_,
		_w3211_
	);
	LUT2 #(
		.INIT('h9)
	) name3178 (
		_w3203_,
		_w3204_,
		_w3212_
	);
	LUT3 #(
		.INIT('h54)
	) name3179 (
		_w3205_,
		_w3210_,
		_w3211_,
		_w3213_
	);
	LUT4 #(
		.INIT('h0180)
	) name3180 (
		\a[20] ,
		\a[21] ,
		\a[22] ,
		\a[23] ,
		_w3214_
	);
	LUT4 #(
		.INIT('h2322)
	) name3181 (
		_w3214_,
		_w374_,
		_w2361_,
		_w37_,
		_w3215_
	);
	LUT3 #(
		.INIT('h96)
	) name3182 (
		_w2959_,
		_w2961_,
		_w2994_,
		_w3216_
	);
	LUT3 #(
		.INIT('h96)
	) name3183 (
		\a[26] ,
		_w3001_,
		_w3216_,
		_w3217_
	);
	LUT4 #(
		.INIT('h127b)
	) name3184 (
		\a[23] ,
		_w3213_,
		_w3215_,
		_w3217_,
		_w3218_
	);
	LUT2 #(
		.INIT('h8)
	) name3185 (
		_w3008_,
		_w3218_,
		_w3219_
	);
	LUT4 #(
		.INIT('h6669)
	) name3186 (
		_w3013_,
		_w3014_,
		_w3064_,
		_w3202_,
		_w3220_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3187 (
		_w587_,
		_w608_,
		_w624_,
		_w2975_,
		_w3221_
	);
	LUT3 #(
		.INIT('h70)
	) name3188 (
		_w666_,
		_w694_,
		_w2874_,
		_w3222_
	);
	LUT3 #(
		.INIT('h70)
	) name3189 (
		_w544_,
		_w558_,
		_w2986_,
		_w3223_
	);
	LUT3 #(
		.INIT('h01)
	) name3190 (
		_w3222_,
		_w3223_,
		_w3221_,
		_w3224_
	);
	LUT4 #(
		.INIT('h6f00)
	) name3191 (
		_w2351_,
		_w2353_,
		_w2875_,
		_w3224_,
		_w3225_
	);
	LUT3 #(
		.INIT('h84)
	) name3192 (
		\a[26] ,
		_w3220_,
		_w3225_,
		_w3226_
	);
	LUT4 #(
		.INIT('h6665)
	) name3193 (
		_w3065_,
		_w3194_,
		_w3195_,
		_w3201_,
		_w3227_
	);
	LUT3 #(
		.INIT('h70)
	) name3194 (
		_w763_,
		_w983_,
		_w2549_,
		_w3228_
	);
	LUT3 #(
		.INIT('h70)
	) name3195 (
		_w871_,
		_w927_,
		_w2617_,
		_w3229_
	);
	LUT3 #(
		.INIT('h70)
	) name3196 (
		_w801_,
		_w851_,
		_w2854_,
		_w3230_
	);
	LUT3 #(
		.INIT('h01)
	) name3197 (
		_w3229_,
		_w3230_,
		_w3228_,
		_w3231_
	);
	LUT4 #(
		.INIT('h6f00)
	) name3198 (
		_w2343_,
		_w2345_,
		_w2550_,
		_w3231_,
		_w3232_
	);
	LUT2 #(
		.INIT('h6)
	) name3199 (
		\a[29] ,
		_w3232_,
		_w3233_
	);
	LUT2 #(
		.INIT('h2)
	) name3200 (
		_w3227_,
		_w3233_,
		_w3234_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3201 (
		_w587_,
		_w608_,
		_w624_,
		_w2986_,
		_w3235_
	);
	LUT3 #(
		.INIT('h70)
	) name3202 (
		_w725_,
		_w764_,
		_w2874_,
		_w3236_
	);
	LUT3 #(
		.INIT('h70)
	) name3203 (
		_w666_,
		_w694_,
		_w2975_,
		_w3237_
	);
	LUT3 #(
		.INIT('h01)
	) name3204 (
		_w3236_,
		_w3237_,
		_w3235_,
		_w3238_
	);
	LUT4 #(
		.INIT('h95aa)
	) name3205 (
		\a[26] ,
		_w2598_,
		_w2875_,
		_w3238_,
		_w3239_
	);
	LUT2 #(
		.INIT('h4)
	) name3206 (
		_w3227_,
		_w3233_,
		_w3240_
	);
	LUT3 #(
		.INIT('h54)
	) name3207 (
		_w3234_,
		_w3239_,
		_w3240_,
		_w3241_
	);
	LUT3 #(
		.INIT('h12)
	) name3208 (
		\a[26] ,
		_w3220_,
		_w3225_,
		_w3242_
	);
	LUT3 #(
		.INIT('h69)
	) name3209 (
		\a[26] ,
		_w3220_,
		_w3225_,
		_w3243_
	);
	LUT3 #(
		.INIT('h54)
	) name3210 (
		_w3226_,
		_w3241_,
		_w3242_,
		_w3244_
	);
	LUT2 #(
		.INIT('h9)
	) name3211 (
		_w3210_,
		_w3212_,
		_w3245_
	);
	LUT2 #(
		.INIT('h4)
	) name3212 (
		_w3244_,
		_w3245_,
		_w3246_
	);
	LUT4 #(
		.INIT('hf400)
	) name3213 (
		_w374_,
		_w2361_,
		_w2404_,
		_w37_,
		_w3247_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name3214 (
		_w3214_,
		_w121_,
		_w418_,
		_w422_,
		_w3248_
	);
	LUT3 #(
		.INIT('h18)
	) name3215 (
		\a[20] ,
		\a[21] ,
		\a[22] ,
		_w3249_
	);
	LUT3 #(
		.INIT('h70)
	) name3216 (
		_w352_,
		_w373_,
		_w3249_,
		_w3250_
	);
	LUT2 #(
		.INIT('h1)
	) name3217 (
		_w3248_,
		_w3250_,
		_w3251_
	);
	LUT3 #(
		.INIT('h9a)
	) name3218 (
		\a[23] ,
		_w3247_,
		_w3251_,
		_w3252_
	);
	LUT2 #(
		.INIT('h2)
	) name3219 (
		_w3244_,
		_w3245_,
		_w3253_
	);
	LUT2 #(
		.INIT('h9)
	) name3220 (
		_w3244_,
		_w3245_,
		_w3254_
	);
	LUT3 #(
		.INIT('h54)
	) name3221 (
		_w3246_,
		_w3252_,
		_w3253_,
		_w3255_
	);
	LUT4 #(
		.INIT('h6996)
	) name3222 (
		\a[23] ,
		_w3213_,
		_w3215_,
		_w3217_,
		_w3256_
	);
	LUT4 #(
		.INIT('h4d00)
	) name3223 (
		_w3244_,
		_w3245_,
		_w3252_,
		_w3256_,
		_w3257_
	);
	LUT4 #(
		.INIT('h54ab)
	) name3224 (
		_w3246_,
		_w3252_,
		_w3253_,
		_w3256_,
		_w3258_
	);
	LUT2 #(
		.INIT('h9)
	) name3225 (
		_w3252_,
		_w3254_,
		_w3259_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name3226 (
		_w3214_,
		_w486_,
		_w487_,
		_w509_,
		_w3260_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3227 (
		_w121_,
		_w418_,
		_w422_,
		_w3249_,
		_w3261_
	);
	LUT4 #(
		.INIT('h6006)
	) name3228 (
		\a[20] ,
		\a[21] ,
		\a[22] ,
		\a[23] ,
		_w3262_
	);
	LUT3 #(
		.INIT('h70)
	) name3229 (
		_w352_,
		_w373_,
		_w3262_,
		_w3263_
	);
	LUT3 #(
		.INIT('h01)
	) name3230 (
		_w3260_,
		_w3261_,
		_w3263_,
		_w3264_
	);
	LUT4 #(
		.INIT('h95aa)
	) name3231 (
		\a[23] ,
		_w2535_,
		_w37_,
		_w3264_,
		_w3265_
	);
	LUT2 #(
		.INIT('h9)
	) name3232 (
		_w3227_,
		_w3233_,
		_w3266_
	);
	LUT2 #(
		.INIT('h9)
	) name3233 (
		_w3196_,
		_w3201_,
		_w3267_
	);
	LUT3 #(
		.INIT('h56)
	) name3234 (
		_w3094_,
		_w3180_,
		_w3187_,
		_w3268_
	);
	LUT3 #(
		.INIT('h70)
	) name3235 (
		_w1202_,
		_w1233_,
		_w2527_,
		_w3269_
	);
	LUT3 #(
		.INIT('h2a)
	) name3236 (
		_w376_,
		_w1325_,
		_w1367_,
		_w3270_
	);
	LUT3 #(
		.INIT('h70)
	) name3237 (
		_w1253_,
		_w1294_,
		_w2407_,
		_w3271_
	);
	LUT3 #(
		.INIT('h01)
	) name3238 (
		_w3270_,
		_w3271_,
		_w3269_,
		_w3272_
	);
	LUT4 #(
		.INIT('h7d00)
	) name3239 (
		_w377_,
		_w2331_,
		_w2333_,
		_w3272_,
		_w3273_
	);
	LUT4 #(
		.INIT('h0056)
	) name3240 (
		_w3094_,
		_w3180_,
		_w3187_,
		_w3273_,
		_w3274_
	);
	LUT3 #(
		.INIT('h70)
	) name3241 (
		_w1136_,
		_w1187_,
		_w2549_,
		_w3275_
	);
	LUT3 #(
		.INIT('h70)
	) name3242 (
		_w1009_,
		_w1050_,
		_w2854_,
		_w3276_
	);
	LUT3 #(
		.INIT('h70)
	) name3243 (
		_w1071_,
		_w1102_,
		_w2617_,
		_w3277_
	);
	LUT3 #(
		.INIT('h01)
	) name3244 (
		_w3276_,
		_w3277_,
		_w3275_,
		_w3278_
	);
	LUT4 #(
		.INIT('h95aa)
	) name3245 (
		\a[29] ,
		_w2550_,
		_w2936_,
		_w3278_,
		_w3279_
	);
	LUT4 #(
		.INIT('ha900)
	) name3246 (
		_w3094_,
		_w3180_,
		_w3187_,
		_w3273_,
		_w3280_
	);
	LUT4 #(
		.INIT('h56a9)
	) name3247 (
		_w3094_,
		_w3180_,
		_w3187_,
		_w3273_,
		_w3281_
	);
	LUT2 #(
		.INIT('h9)
	) name3248 (
		_w3188_,
		_w3190_,
		_w3282_
	);
	LUT4 #(
		.INIT('h2b00)
	) name3249 (
		_w3268_,
		_w3273_,
		_w3279_,
		_w3282_,
		_w3283_
	);
	LUT4 #(
		.INIT('h00d4)
	) name3250 (
		_w3268_,
		_w3273_,
		_w3279_,
		_w3282_,
		_w3284_
	);
	LUT3 #(
		.INIT('h70)
	) name3251 (
		_w1071_,
		_w1102_,
		_w2549_,
		_w3285_
	);
	LUT3 #(
		.INIT('h70)
	) name3252 (
		_w763_,
		_w983_,
		_w2854_,
		_w3286_
	);
	LUT3 #(
		.INIT('h70)
	) name3253 (
		_w1009_,
		_w1050_,
		_w2617_,
		_w3287_
	);
	LUT3 #(
		.INIT('h01)
	) name3254 (
		_w3286_,
		_w3287_,
		_w3285_,
		_w3288_
	);
	LUT4 #(
		.INIT('h6f00)
	) name3255 (
		_w2339_,
		_w2341_,
		_w2550_,
		_w3288_,
		_w3289_
	);
	LUT2 #(
		.INIT('h6)
	) name3256 (
		\a[29] ,
		_w3289_,
		_w3290_
	);
	LUT3 #(
		.INIT('h54)
	) name3257 (
		_w3283_,
		_w3284_,
		_w3290_,
		_w3291_
	);
	LUT3 #(
		.INIT('h70)
	) name3258 (
		_w725_,
		_w764_,
		_w2975_,
		_w3292_
	);
	LUT3 #(
		.INIT('h70)
	) name3259 (
		_w801_,
		_w851_,
		_w2874_,
		_w3293_
	);
	LUT3 #(
		.INIT('h70)
	) name3260 (
		_w666_,
		_w694_,
		_w2986_,
		_w3294_
	);
	LUT3 #(
		.INIT('h01)
	) name3261 (
		_w3293_,
		_w3294_,
		_w3292_,
		_w3295_
	);
	LUT4 #(
		.INIT('h6f00)
	) name3262 (
		_w2347_,
		_w2349_,
		_w2875_,
		_w3295_,
		_w3296_
	);
	LUT4 #(
		.INIT('h71b2)
	) name3263 (
		\a[26] ,
		_w3267_,
		_w3291_,
		_w3296_,
		_w3297_
	);
	LUT3 #(
		.INIT('h09)
	) name3264 (
		_w3239_,
		_w3266_,
		_w3297_,
		_w3298_
	);
	LUT3 #(
		.INIT('h60)
	) name3265 (
		_w3239_,
		_w3266_,
		_w3297_,
		_w3299_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3266 (
		_w486_,
		_w487_,
		_w509_,
		_w3249_,
		_w3300_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3267 (
		_w121_,
		_w418_,
		_w422_,
		_w3262_,
		_w3301_
	);
	LUT3 #(
		.INIT('h2a)
	) name3268 (
		_w3214_,
		_w544_,
		_w558_,
		_w3302_
	);
	LUT3 #(
		.INIT('h01)
	) name3269 (
		_w3300_,
		_w3301_,
		_w3302_,
		_w3303_
	);
	LUT4 #(
		.INIT('h6f00)
	) name3270 (
		_w2355_,
		_w2357_,
		_w37_,
		_w3303_,
		_w3304_
	);
	LUT4 #(
		.INIT('h3132)
	) name3271 (
		\a[23] ,
		_w3298_,
		_w3299_,
		_w3304_,
		_w3305_
	);
	LUT2 #(
		.INIT('h9)
	) name3272 (
		_w3241_,
		_w3243_,
		_w3306_
	);
	LUT3 #(
		.INIT('h8e)
	) name3273 (
		_w3265_,
		_w3305_,
		_w3306_,
		_w3307_
	);
	LUT3 #(
		.INIT('h09)
	) name3274 (
		_w3252_,
		_w3254_,
		_w3307_,
		_w3308_
	);
	LUT3 #(
		.INIT('h96)
	) name3275 (
		_w3265_,
		_w3305_,
		_w3306_,
		_w3309_
	);
	LUT2 #(
		.INIT('h9)
	) name3276 (
		\a[17] ,
		\a[18] ,
		_w3310_
	);
	LUT4 #(
		.INIT('h0180)
	) name3277 (
		\a[17] ,
		\a[18] ,
		\a[19] ,
		\a[20] ,
		_w3311_
	);
	LUT4 #(
		.INIT('h0660)
	) name3278 (
		\a[17] ,
		\a[18] ,
		\a[19] ,
		\a[20] ,
		_w3312_
	);
	LUT4 #(
		.INIT('h5150)
	) name3279 (
		_w374_,
		_w2361_,
		_w3311_,
		_w3312_,
		_w3313_
	);
	LUT3 #(
		.INIT('h70)
	) name3280 (
		_w725_,
		_w764_,
		_w2986_,
		_w3314_
	);
	LUT3 #(
		.INIT('h70)
	) name3281 (
		_w801_,
		_w851_,
		_w2975_,
		_w3315_
	);
	LUT3 #(
		.INIT('h70)
	) name3282 (
		_w871_,
		_w927_,
		_w2874_,
		_w3316_
	);
	LUT3 #(
		.INIT('h01)
	) name3283 (
		_w3315_,
		_w3316_,
		_w3314_,
		_w3317_
	);
	LUT4 #(
		.INIT('h95aa)
	) name3284 (
		\a[26] ,
		_w2724_,
		_w2875_,
		_w3317_,
		_w3318_
	);
	LUT4 #(
		.INIT('h54ab)
	) name3285 (
		_w3274_,
		_w3279_,
		_w3280_,
		_w3282_,
		_w3319_
	);
	LUT2 #(
		.INIT('h9)
	) name3286 (
		_w3290_,
		_w3319_,
		_w3320_
	);
	LUT4 #(
		.INIT('h135f)
	) name3287 (
		_w78_,
		_w56_,
		_w41_,
		_w39_,
		_w3321_
	);
	LUT3 #(
		.INIT('h40)
	) name3288 (
		_w441_,
		_w2082_,
		_w3321_,
		_w3322_
	);
	LUT3 #(
		.INIT('h80)
	) name3289 (
		_w168_,
		_w806_,
		_w2169_,
		_w3323_
	);
	LUT4 #(
		.INIT('h135f)
	) name3290 (
		_w85_,
		_w67_,
		_w184_,
		_w236_,
		_w3324_
	);
	LUT4 #(
		.INIT('h153f)
	) name3291 (
		_w41_,
		_w50_,
		_w259_,
		_w176_,
		_w3325_
	);
	LUT4 #(
		.INIT('h4000)
	) name3292 (
		_w398_,
		_w492_,
		_w3324_,
		_w3325_,
		_w3326_
	);
	LUT3 #(
		.INIT('h80)
	) name3293 (
		_w3322_,
		_w3323_,
		_w3326_,
		_w3327_
	);
	LUT4 #(
		.INIT('h135f)
	) name3294 (
		_w72_,
		_w43_,
		_w65_,
		_w44_,
		_w3328_
	);
	LUT3 #(
		.INIT('h57)
	) name3295 (
		_w122_,
		_w59_,
		_w47_,
		_w3329_
	);
	LUT4 #(
		.INIT('h4000)
	) name3296 (
		_w137_,
		_w803_,
		_w3329_,
		_w3328_,
		_w3330_
	);
	LUT2 #(
		.INIT('h8)
	) name3297 (
		_w719_,
		_w3330_,
		_w3331_
	);
	LUT4 #(
		.INIT('h135f)
	) name3298 (
		_w50_,
		_w93_,
		_w236_,
		_w176_,
		_w3332_
	);
	LUT4 #(
		.INIT('h153f)
	) name3299 (
		_w90_,
		_w65_,
		_w419_,
		_w430_,
		_w3333_
	);
	LUT4 #(
		.INIT('h8000)
	) name3300 (
		_w1143_,
		_w2745_,
		_w3332_,
		_w3333_,
		_w3334_
	);
	LUT4 #(
		.INIT('h153f)
	) name3301 (
		_w65_,
		_w46_,
		_w236_,
		_w158_,
		_w3335_
	);
	LUT4 #(
		.INIT('h153f)
	) name3302 (
		_w59_,
		_w56_,
		_w201_,
		_w259_,
		_w3336_
	);
	LUT4 #(
		.INIT('h8000)
	) name3303 (
		_w997_,
		_w2125_,
		_w3335_,
		_w3336_,
		_w3337_
	);
	LUT3 #(
		.INIT('h80)
	) name3304 (
		_w1836_,
		_w3334_,
		_w3337_,
		_w3338_
	);
	LUT3 #(
		.INIT('h80)
	) name3305 (
		_w3327_,
		_w3331_,
		_w3338_,
		_w3339_
	);
	LUT4 #(
		.INIT('h8000)
	) name3306 (
		_w292_,
		_w643_,
		_w687_,
		_w1222_,
		_w3340_
	);
	LUT4 #(
		.INIT('h153f)
	) name3307 (
		_w59_,
		_w67_,
		_w72_,
		_w39_,
		_w3341_
	);
	LUT4 #(
		.INIT('h153f)
	) name3308 (
		_w85_,
		_w56_,
		_w43_,
		_w176_,
		_w3342_
	);
	LUT4 #(
		.INIT('h8000)
	) name3309 (
		_w132_,
		_w776_,
		_w3341_,
		_w3342_,
		_w3343_
	);
	LUT2 #(
		.INIT('h8)
	) name3310 (
		_w3340_,
		_w3343_,
		_w3344_
	);
	LUT3 #(
		.INIT('h40)
	) name3311 (
		_w142_,
		_w902_,
		_w940_,
		_w3345_
	);
	LUT4 #(
		.INIT('h153f)
	) name3312 (
		_w47_,
		_w41_,
		_w236_,
		_w259_,
		_w3346_
	);
	LUT4 #(
		.INIT('h8000)
	) name3313 (
		_w1726_,
		_w2625_,
		_w3022_,
		_w3346_,
		_w3347_
	);
	LUT3 #(
		.INIT('h80)
	) name3314 (
		_w932_,
		_w3345_,
		_w3347_,
		_w3348_
	);
	LUT3 #(
		.INIT('h20)
	) name3315 (
		_w150_,
		_w170_,
		_w2510_,
		_w3349_
	);
	LUT4 #(
		.INIT('h135f)
	) name3316 (
		_w122_,
		_w59_,
		_w56_,
		_w158_,
		_w3350_
	);
	LUT3 #(
		.INIT('h80)
	) name3317 (
		_w2468_,
		_w2560_,
		_w3350_,
		_w3351_
	);
	LUT4 #(
		.INIT('h153f)
	) name3318 (
		_w55_,
		_w65_,
		_w378_,
		_w430_,
		_w3352_
	);
	LUT4 #(
		.INIT('h8000)
	) name3319 (
		_w427_,
		_w962_,
		_w1456_,
		_w3352_,
		_w3353_
	);
	LUT3 #(
		.INIT('h80)
	) name3320 (
		_w3349_,
		_w3351_,
		_w3353_,
		_w3354_
	);
	LUT4 #(
		.INIT('h4000)
	) name3321 (
		_w468_,
		_w882_,
		_w2502_,
		_w2503_,
		_w3355_
	);
	LUT4 #(
		.INIT('h8000)
	) name3322 (
		_w2580_,
		_w2583_,
		_w2756_,
		_w3355_,
		_w3356_
	);
	LUT2 #(
		.INIT('h8)
	) name3323 (
		_w3354_,
		_w3356_,
		_w3357_
	);
	LUT4 #(
		.INIT('h8000)
	) name3324 (
		_w3344_,
		_w3348_,
		_w3354_,
		_w3356_,
		_w3358_
	);
	LUT2 #(
		.INIT('h8)
	) name3325 (
		_w3339_,
		_w3358_,
		_w3359_
	);
	LUT2 #(
		.INIT('h2)
	) name3326 (
		_w3139_,
		_w3359_,
		_w3360_
	);
	LUT2 #(
		.INIT('h9)
	) name3327 (
		_w3139_,
		_w3359_,
		_w3361_
	);
	LUT4 #(
		.INIT('h54ab)
	) name3328 (
		_w1547_,
		_w2323_,
		_w2324_,
		_w2326_,
		_w3362_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3329 (
		_w1454_,
		_w1426_,
		_w1478_,
		_w2407_,
		_w3363_
	);
	LUT3 #(
		.INIT('h70)
	) name3330 (
		_w1381_,
		_w1398_,
		_w2527_,
		_w3364_
	);
	LUT3 #(
		.INIT('h2a)
	) name3331 (
		_w376_,
		_w1501_,
		_w1545_,
		_w3365_
	);
	LUT3 #(
		.INIT('h01)
	) name3332 (
		_w3364_,
		_w3365_,
		_w3363_,
		_w3366_
	);
	LUT4 #(
		.INIT('h80cc)
	) name3333 (
		_w377_,
		_w3361_,
		_w3362_,
		_w3366_,
		_w3367_
	);
	LUT3 #(
		.INIT('h96)
	) name3334 (
		\a[14] ,
		_w3139_,
		_w3179_,
		_w3368_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name3335 (
		_w376_,
		_w1454_,
		_w1426_,
		_w1478_,
		_w3369_
	);
	LUT3 #(
		.INIT('h70)
	) name3336 (
		_w1325_,
		_w1367_,
		_w2527_,
		_w3370_
	);
	LUT3 #(
		.INIT('h70)
	) name3337 (
		_w1381_,
		_w1398_,
		_w2407_,
		_w3371_
	);
	LUT3 #(
		.INIT('h01)
	) name3338 (
		_w3370_,
		_w3371_,
		_w3369_,
		_w3372_
	);
	LUT4 #(
		.INIT('h7d00)
	) name3339 (
		_w377_,
		_w2327_,
		_w2329_,
		_w3372_,
		_w3373_
	);
	LUT4 #(
		.INIT('hf110)
	) name3340 (
		_w3360_,
		_w3367_,
		_w3368_,
		_w3373_,
		_w3374_
	);
	LUT4 #(
		.INIT('hc993)
	) name3341 (
		\a[14] ,
		_w3092_,
		_w3139_,
		_w3179_,
		_w3375_
	);
	LUT4 #(
		.INIT('h708f)
	) name3342 (
		_w377_,
		_w3182_,
		_w3186_,
		_w3375_,
		_w3376_
	);
	LUT2 #(
		.INIT('h4)
	) name3343 (
		_w3374_,
		_w3376_,
		_w3377_
	);
	LUT2 #(
		.INIT('h2)
	) name3344 (
		_w3374_,
		_w3376_,
		_w3378_
	);
	LUT2 #(
		.INIT('h9)
	) name3345 (
		_w3374_,
		_w3376_,
		_w3379_
	);
	LUT3 #(
		.INIT('h70)
	) name3346 (
		_w1136_,
		_w1187_,
		_w2617_,
		_w3380_
	);
	LUT3 #(
		.INIT('h70)
	) name3347 (
		_w1071_,
		_w1102_,
		_w2854_,
		_w3381_
	);
	LUT3 #(
		.INIT('h70)
	) name3348 (
		_w1202_,
		_w1233_,
		_w2549_,
		_w3382_
	);
	LUT3 #(
		.INIT('h01)
	) name3349 (
		_w3381_,
		_w3382_,
		_w3380_,
		_w3383_
	);
	LUT4 #(
		.INIT('h6f00)
	) name3350 (
		_w2335_,
		_w2337_,
		_w2550_,
		_w3383_,
		_w3384_
	);
	LUT4 #(
		.INIT('h3132)
	) name3351 (
		\a[29] ,
		_w3377_,
		_w3378_,
		_w3384_,
		_w3385_
	);
	LUT3 #(
		.INIT('h09)
	) name3352 (
		_w3279_,
		_w3281_,
		_w3385_,
		_w3386_
	);
	LUT3 #(
		.INIT('h60)
	) name3353 (
		_w3279_,
		_w3281_,
		_w3385_,
		_w3387_
	);
	LUT3 #(
		.INIT('h70)
	) name3354 (
		_w763_,
		_w983_,
		_w2874_,
		_w3388_
	);
	LUT3 #(
		.INIT('h70)
	) name3355 (
		_w871_,
		_w927_,
		_w2975_,
		_w3389_
	);
	LUT3 #(
		.INIT('h70)
	) name3356 (
		_w801_,
		_w851_,
		_w2986_,
		_w3390_
	);
	LUT3 #(
		.INIT('h01)
	) name3357 (
		_w3389_,
		_w3390_,
		_w3388_,
		_w3391_
	);
	LUT4 #(
		.INIT('h6f00)
	) name3358 (
		_w2343_,
		_w2345_,
		_w2875_,
		_w3391_,
		_w3392_
	);
	LUT4 #(
		.INIT('h3132)
	) name3359 (
		\a[26] ,
		_w3386_,
		_w3387_,
		_w3392_,
		_w3393_
	);
	LUT3 #(
		.INIT('hb2)
	) name3360 (
		_w3318_,
		_w3320_,
		_w3393_,
		_w3394_
	);
	LUT4 #(
		.INIT('h6996)
	) name3361 (
		\a[26] ,
		_w3267_,
		_w3291_,
		_w3296_,
		_w3395_
	);
	LUT2 #(
		.INIT('h4)
	) name3362 (
		_w3394_,
		_w3395_,
		_w3396_
	);
	LUT2 #(
		.INIT('h2)
	) name3363 (
		_w3394_,
		_w3395_,
		_w3397_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3364 (
		_w486_,
		_w487_,
		_w509_,
		_w3262_,
		_w3398_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name3365 (
		_w3214_,
		_w587_,
		_w608_,
		_w624_,
		_w3399_
	);
	LUT3 #(
		.INIT('h70)
	) name3366 (
		_w544_,
		_w558_,
		_w3249_,
		_w3400_
	);
	LUT3 #(
		.INIT('h01)
	) name3367 (
		_w3398_,
		_w3399_,
		_w3400_,
		_w3401_
	);
	LUT4 #(
		.INIT('h95aa)
	) name3368 (
		\a[23] ,
		_w2526_,
		_w37_,
		_w3401_,
		_w3402_
	);
	LUT3 #(
		.INIT('h54)
	) name3369 (
		_w3396_,
		_w3397_,
		_w3402_,
		_w3403_
	);
	LUT3 #(
		.INIT('h96)
	) name3370 (
		_w3239_,
		_w3266_,
		_w3297_,
		_w3404_
	);
	LUT3 #(
		.INIT('h69)
	) name3371 (
		\a[23] ,
		_w3304_,
		_w3404_,
		_w3405_
	);
	LUT4 #(
		.INIT('h90f9)
	) name3372 (
		\a[20] ,
		_w3313_,
		_w3403_,
		_w3405_,
		_w3406_
	);
	LUT2 #(
		.INIT('h2)
	) name3373 (
		_w3309_,
		_w3406_,
		_w3407_
	);
	LUT2 #(
		.INIT('h4)
	) name3374 (
		_w3309_,
		_w3406_,
		_w3408_
	);
	LUT2 #(
		.INIT('h9)
	) name3375 (
		_w3309_,
		_w3406_,
		_w3409_
	);
	LUT4 #(
		.INIT('h9669)
	) name3376 (
		\a[20] ,
		_w3313_,
		_w3403_,
		_w3405_,
		_w3410_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3377 (
		_w587_,
		_w608_,
		_w624_,
		_w3249_,
		_w3411_
	);
	LUT3 #(
		.INIT('h2a)
	) name3378 (
		_w3214_,
		_w666_,
		_w694_,
		_w3412_
	);
	LUT3 #(
		.INIT('h70)
	) name3379 (
		_w544_,
		_w558_,
		_w3262_,
		_w3413_
	);
	LUT3 #(
		.INIT('h01)
	) name3380 (
		_w3412_,
		_w3413_,
		_w3411_,
		_w3414_
	);
	LUT4 #(
		.INIT('h6f00)
	) name3381 (
		_w2351_,
		_w2353_,
		_w37_,
		_w3414_,
		_w3415_
	);
	LUT3 #(
		.INIT('h96)
	) name3382 (
		_w3318_,
		_w3320_,
		_w3393_,
		_w3416_
	);
	LUT3 #(
		.INIT('h90)
	) name3383 (
		\a[23] ,
		_w3415_,
		_w3416_,
		_w3417_
	);
	LUT3 #(
		.INIT('h06)
	) name3384 (
		\a[23] ,
		_w3415_,
		_w3416_,
		_w3418_
	);
	LUT3 #(
		.INIT('h69)
	) name3385 (
		\a[23] ,
		_w3415_,
		_w3416_,
		_w3419_
	);
	LUT3 #(
		.INIT('h96)
	) name3386 (
		_w3279_,
		_w3281_,
		_w3385_,
		_w3420_
	);
	LUT3 #(
		.INIT('h69)
	) name3387 (
		\a[26] ,
		_w3392_,
		_w3420_,
		_w3421_
	);
	LUT3 #(
		.INIT('h70)
	) name3388 (
		_w1202_,
		_w1233_,
		_w2617_,
		_w3422_
	);
	LUT3 #(
		.INIT('h70)
	) name3389 (
		_w1253_,
		_w1294_,
		_w2549_,
		_w3423_
	);
	LUT3 #(
		.INIT('h70)
	) name3390 (
		_w1136_,
		_w1187_,
		_w2854_,
		_w3424_
	);
	LUT3 #(
		.INIT('h01)
	) name3391 (
		_w3423_,
		_w3424_,
		_w3422_,
		_w3425_
	);
	LUT4 #(
		.INIT('h95aa)
	) name3392 (
		\a[29] ,
		_w2550_,
		_w3067_,
		_w3425_,
		_w3426_
	);
	LUT4 #(
		.INIT('he11e)
	) name3393 (
		_w3360_,
		_w3367_,
		_w3368_,
		_w3373_,
		_w3427_
	);
	LUT4 #(
		.INIT('h6c33)
	) name3394 (
		_w377_,
		_w3361_,
		_w3362_,
		_w3366_,
		_w3428_
	);
	LUT3 #(
		.INIT('h20)
	) name3395 (
		_w384_,
		_w461_,
		_w2517_,
		_w3429_
	);
	LUT4 #(
		.INIT('h153f)
	) name3396 (
		_w106_,
		_w50_,
		_w43_,
		_w46_,
		_w3430_
	);
	LUT4 #(
		.INIT('h8000)
	) name3397 (
		_w1138_,
		_w2369_,
		_w2826_,
		_w3430_,
		_w3431_
	);
	LUT4 #(
		.INIT('h0777)
	) name3398 (
		_w47_,
		_w72_,
		_w39_,
		_w65_,
		_w3432_
	);
	LUT4 #(
		.INIT('h153f)
	) name3399 (
		_w38_,
		_w122_,
		_w47_,
		_w166_,
		_w3433_
	);
	LUT4 #(
		.INIT('h1000)
	) name3400 (
		_w190_,
		_w457_,
		_w3432_,
		_w3433_,
		_w3434_
	);
	LUT3 #(
		.INIT('h80)
	) name3401 (
		_w3429_,
		_w3431_,
		_w3434_,
		_w3435_
	);
	LUT4 #(
		.INIT('h8000)
	) name3402 (
		_w1623_,
		_w1626_,
		_w3126_,
		_w3128_,
		_w3436_
	);
	LUT4 #(
		.INIT('h153f)
	) name3403 (
		_w41_,
		_w50_,
		_w236_,
		_w419_,
		_w3437_
	);
	LUT4 #(
		.INIT('h4000)
	) name3404 (
		_w45_,
		_w707_,
		_w1427_,
		_w3437_,
		_w3438_
	);
	LUT4 #(
		.INIT('h153f)
	) name3405 (
		_w52_,
		_w110_,
		_w39_,
		_w158_,
		_w3439_
	);
	LUT4 #(
		.INIT('h1000)
	) name3406 (
		_w295_,
		_w286_,
		_w1762_,
		_w3439_,
		_w3440_
	);
	LUT4 #(
		.INIT('h153f)
	) name3407 (
		_w67_,
		_w65_,
		_w201_,
		_w176_,
		_w3441_
	);
	LUT3 #(
		.INIT('h37)
	) name3408 (
		_w38_,
		_w72_,
		_w44_,
		_w3442_
	);
	LUT4 #(
		.INIT('h8000)
	) name3409 (
		_w1687_,
		_w1865_,
		_w3442_,
		_w3441_,
		_w3443_
	);
	LUT4 #(
		.INIT('h135f)
	) name3410 (
		_w38_,
		_w85_,
		_w184_,
		_w158_,
		_w3444_
	);
	LUT4 #(
		.INIT('h8000)
	) name3411 (
		_w1046_,
		_w1137_,
		_w2706_,
		_w3444_,
		_w3445_
	);
	LUT4 #(
		.INIT('h8000)
	) name3412 (
		_w3443_,
		_w3445_,
		_w3438_,
		_w3440_,
		_w3446_
	);
	LUT4 #(
		.INIT('h135f)
	) name3413 (
		_w47_,
		_w93_,
		_w166_,
		_w176_,
		_w3447_
	);
	LUT4 #(
		.INIT('h8000)
	) name3414 (
		_w676_,
		_w1472_,
		_w2135_,
		_w3447_,
		_w3448_
	);
	LUT4 #(
		.INIT('h153f)
	) name3415 (
		_w59_,
		_w78_,
		_w90_,
		_w430_,
		_w3449_
	);
	LUT2 #(
		.INIT('h8)
	) name3416 (
		_w522_,
		_w3449_,
		_w3450_
	);
	LUT4 #(
		.INIT('h135f)
	) name3417 (
		_w59_,
		_w90_,
		_w72_,
		_w184_,
		_w3451_
	);
	LUT4 #(
		.INIT('h153f)
	) name3418 (
		_w55_,
		_w93_,
		_w158_,
		_w176_,
		_w3452_
	);
	LUT4 #(
		.INIT('h8000)
	) name3419 (
		_w252_,
		_w344_,
		_w3451_,
		_w3452_,
		_w3453_
	);
	LUT3 #(
		.INIT('h80)
	) name3420 (
		_w3450_,
		_w3448_,
		_w3453_,
		_w3454_
	);
	LUT4 #(
		.INIT('h8000)
	) name3421 (
		_w3446_,
		_w3454_,
		_w3435_,
		_w3436_,
		_w3455_
	);
	LUT2 #(
		.INIT('h8)
	) name3422 (
		_w871_,
		_w3455_,
		_w3456_
	);
	LUT4 #(
		.INIT('h153f)
	) name3423 (
		_w59_,
		_w110_,
		_w78_,
		_w158_,
		_w3457_
	);
	LUT4 #(
		.INIT('h4000)
	) name3424 (
		_w481_,
		_w2758_,
		_w3113_,
		_w3457_,
		_w3458_
	);
	LUT4 #(
		.INIT('h135f)
	) name3425 (
		_w122_,
		_w106_,
		_w47_,
		_w46_,
		_w3459_
	);
	LUT4 #(
		.INIT('h153f)
	) name3426 (
		_w38_,
		_w90_,
		_w419_,
		_w430_,
		_w3460_
	);
	LUT4 #(
		.INIT('h8000)
	) name3427 (
		_w1079_,
		_w1190_,
		_w3459_,
		_w3460_,
		_w3461_
	);
	LUT2 #(
		.INIT('h8)
	) name3428 (
		_w3458_,
		_w3461_,
		_w3462_
	);
	LUT4 #(
		.INIT('h8000)
	) name3429 (
		_w403_,
		_w1278_,
		_w1423_,
		_w1664_,
		_w3463_
	);
	LUT4 #(
		.INIT('h135f)
	) name3430 (
		_w38_,
		_w65_,
		_w184_,
		_w236_,
		_w3464_
	);
	LUT2 #(
		.INIT('h4)
	) name3431 (
		_w436_,
		_w3464_,
		_w3465_
	);
	LUT4 #(
		.INIT('h153f)
	) name3432 (
		_w110_,
		_w72_,
		_w44_,
		_w176_,
		_w3466_
	);
	LUT4 #(
		.INIT('h153f)
	) name3433 (
		_w55_,
		_w59_,
		_w176_,
		_w419_,
		_w3467_
	);
	LUT4 #(
		.INIT('h4000)
	) name3434 (
		_w436_,
		_w3464_,
		_w3466_,
		_w3467_,
		_w3468_
	);
	LUT4 #(
		.INIT('h153f)
	) name3435 (
		_w90_,
		_w41_,
		_w236_,
		_w430_,
		_w3469_
	);
	LUT4 #(
		.INIT('h8000)
	) name3436 (
		_w1683_,
		_w1738_,
		_w2392_,
		_w3469_,
		_w3470_
	);
	LUT4 #(
		.INIT('h8000)
	) name3437 (
		_w1062_,
		_w3470_,
		_w3463_,
		_w3468_,
		_w3471_
	);
	LUT2 #(
		.INIT('h8)
	) name3438 (
		_w3462_,
		_w3471_,
		_w3472_
	);
	LUT4 #(
		.INIT('h135f)
	) name3439 (
		_w38_,
		_w85_,
		_w78_,
		_w166_,
		_w3473_
	);
	LUT4 #(
		.INIT('h0777)
	) name3440 (
		_w38_,
		_w106_,
		_w67_,
		_w39_,
		_w3474_
	);
	LUT4 #(
		.INIT('h2000)
	) name3441 (
		_w260_,
		_w365_,
		_w3474_,
		_w3473_,
		_w3475_
	);
	LUT4 #(
		.INIT('h8000)
	) name3442 (
		_w112_,
		_w283_,
		_w1301_,
		_w2379_,
		_w3476_
	);
	LUT4 #(
		.INIT('h8000)
	) name3443 (
		_w1137_,
		_w1173_,
		_w1257_,
		_w3103_,
		_w3477_
	);
	LUT4 #(
		.INIT('h8000)
	) name3444 (
		_w564_,
		_w663_,
		_w820_,
		_w906_,
		_w3478_
	);
	LUT4 #(
		.INIT('h8000)
	) name3445 (
		_w3477_,
		_w3478_,
		_w3475_,
		_w3476_,
		_w3479_
	);
	LUT4 #(
		.INIT('h8000)
	) name3446 (
		_w2631_,
		_w2773_,
		_w3454_,
		_w3479_,
		_w3480_
	);
	LUT2 #(
		.INIT('h8)
	) name3447 (
		_w3472_,
		_w3480_,
		_w3481_
	);
	LUT4 #(
		.INIT('h0777)
	) name3448 (
		_w871_,
		_w3455_,
		_w3472_,
		_w3480_,
		_w3482_
	);
	LUT4 #(
		.INIT('h8000)
	) name3449 (
		_w871_,
		_w3455_,
		_w3472_,
		_w3480_,
		_w3483_
	);
	LUT4 #(
		.INIT('h044c)
	) name3450 (
		\a[11] ,
		_w3139_,
		_w3456_,
		_w3481_,
		_w3484_
	);
	LUT4 #(
		.INIT('h3220)
	) name3451 (
		\a[11] ,
		_w3139_,
		_w3456_,
		_w3481_,
		_w3485_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3452 (
		_w1454_,
		_w1426_,
		_w1478_,
		_w2527_,
		_w3486_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name3453 (
		_w376_,
		_w1584_,
		_w1569_,
		_w1606_,
		_w3487_
	);
	LUT3 #(
		.INIT('h70)
	) name3454 (
		_w1501_,
		_w1545_,
		_w2407_,
		_w3488_
	);
	LUT3 #(
		.INIT('h01)
	) name3455 (
		_w3487_,
		_w3488_,
		_w3486_,
		_w3489_
	);
	LUT4 #(
		.INIT('h7d00)
	) name3456 (
		_w377_,
		_w2323_,
		_w2325_,
		_w3489_,
		_w3490_
	);
	LUT3 #(
		.INIT('h54)
	) name3457 (
		_w3484_,
		_w3485_,
		_w3490_,
		_w3491_
	);
	LUT2 #(
		.INIT('h2)
	) name3458 (
		_w3428_,
		_w3491_,
		_w3492_
	);
	LUT2 #(
		.INIT('h9)
	) name3459 (
		_w3428_,
		_w3491_,
		_w3493_
	);
	LUT3 #(
		.INIT('ha9)
	) name3460 (
		\a[11] ,
		_w3482_,
		_w3483_,
		_w3494_
	);
	LUT4 #(
		.INIT('h54ab)
	) name3461 (
		_w1663_,
		_w2319_,
		_w2320_,
		_w2322_,
		_w3495_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3462 (
		_w1584_,
		_w1569_,
		_w1606_,
		_w2407_,
		_w3496_
	);
	LUT3 #(
		.INIT('h70)
	) name3463 (
		_w1501_,
		_w1545_,
		_w2527_,
		_w3497_
	);
	LUT3 #(
		.INIT('h2a)
	) name3464 (
		_w376_,
		_w1620_,
		_w1661_,
		_w3498_
	);
	LUT3 #(
		.INIT('h01)
	) name3465 (
		_w3496_,
		_w3497_,
		_w3498_,
		_w3499_
	);
	LUT4 #(
		.INIT('h2033)
	) name3466 (
		_w377_,
		_w3494_,
		_w3495_,
		_w3499_,
		_w3500_
	);
	LUT4 #(
		.INIT('h153f)
	) name3467 (
		_w52_,
		_w78_,
		_w90_,
		_w158_,
		_w3501_
	);
	LUT4 #(
		.INIT('h4000)
	) name3468 (
		_w461_,
		_w1208_,
		_w1209_,
		_w3501_,
		_w3502_
	);
	LUT4 #(
		.INIT('h135f)
	) name3469 (
		_w56_,
		_w50_,
		_w43_,
		_w419_,
		_w3503_
	);
	LUT3 #(
		.INIT('h57)
	) name3470 (
		_w106_,
		_w52_,
		_w90_,
		_w3504_
	);
	LUT2 #(
		.INIT('h8)
	) name3471 (
		_w1576_,
		_w3504_,
		_w3505_
	);
	LUT4 #(
		.INIT('h8000)
	) name3472 (
		_w1427_,
		_w1576_,
		_w3503_,
		_w3504_,
		_w3506_
	);
	LUT4 #(
		.INIT('h135f)
	) name3473 (
		_w59_,
		_w56_,
		_w39_,
		_w184_,
		_w3507_
	);
	LUT4 #(
		.INIT('h135f)
	) name3474 (
		_w55_,
		_w67_,
		_w78_,
		_w419_,
		_w3508_
	);
	LUT3 #(
		.INIT('h80)
	) name3475 (
		_w1374_,
		_w3507_,
		_w3508_,
		_w3509_
	);
	LUT4 #(
		.INIT('h153f)
	) name3476 (
		_w38_,
		_w122_,
		_w110_,
		_w72_,
		_w3510_
	);
	LUT4 #(
		.INIT('h8000)
	) name3477 (
		_w1837_,
		_w1858_,
		_w2117_,
		_w3510_,
		_w3511_
	);
	LUT4 #(
		.INIT('h8000)
	) name3478 (
		_w3509_,
		_w3511_,
		_w3502_,
		_w3506_,
		_w3512_
	);
	LUT3 #(
		.INIT('h80)
	) name3479 (
		_w1612_,
		_w2646_,
		_w3512_,
		_w3513_
	);
	LUT3 #(
		.INIT('h80)
	) name3480 (
		_w1136_,
		_w1642_,
		_w3513_,
		_w3514_
	);
	LUT2 #(
		.INIT('h2)
	) name3481 (
		_w3456_,
		_w3514_,
		_w3515_
	);
	LUT2 #(
		.INIT('h4)
	) name3482 (
		_w3456_,
		_w3514_,
		_w3516_
	);
	LUT2 #(
		.INIT('h9)
	) name3483 (
		_w3456_,
		_w3514_,
		_w3517_
	);
	LUT4 #(
		.INIT('h135f)
	) name3484 (
		_w67_,
		_w46_,
		_w236_,
		_w166_,
		_w3518_
	);
	LUT4 #(
		.INIT('h4000)
	) name3485 (
		_w315_,
		_w2072_,
		_w3346_,
		_w3518_,
		_w3519_
	);
	LUT4 #(
		.INIT('h0777)
	) name3486 (
		_w59_,
		_w78_,
		_w46_,
		_w419_,
		_w3520_
	);
	LUT4 #(
		.INIT('h153f)
	) name3487 (
		_w110_,
		_w44_,
		_w166_,
		_w378_,
		_w3521_
	);
	LUT3 #(
		.INIT('h80)
	) name3488 (
		_w1447_,
		_w3521_,
		_w3520_,
		_w3522_
	);
	LUT3 #(
		.INIT('h80)
	) name3489 (
		_w1768_,
		_w3519_,
		_w3522_,
		_w3523_
	);
	LUT4 #(
		.INIT('h153f)
	) name3490 (
		_w110_,
		_w72_,
		_w44_,
		_w184_,
		_w3524_
	);
	LUT2 #(
		.INIT('h4)
	) name3491 (
		_w398_,
		_w3524_,
		_w3525_
	);
	LUT3 #(
		.INIT('h80)
	) name3492 (
		_w191_,
		_w1700_,
		_w2624_,
		_w3526_
	);
	LUT2 #(
		.INIT('h8)
	) name3493 (
		_w3525_,
		_w3526_,
		_w3527_
	);
	LUT4 #(
		.INIT('h4000)
	) name3494 (
		_w86_,
		_w908_,
		_w985_,
		_w1078_,
		_w3528_
	);
	LUT4 #(
		.INIT('h8000)
	) name3495 (
		_w284_,
		_w290_,
		_w3465_,
		_w3528_,
		_w3529_
	);
	LUT3 #(
		.INIT('h80)
	) name3496 (
		_w3527_,
		_w3523_,
		_w3529_,
		_w3530_
	);
	LUT4 #(
		.INIT('h135f)
	) name3497 (
		_w78_,
		_w93_,
		_w65_,
		_w259_,
		_w3531_
	);
	LUT3 #(
		.INIT('h57)
	) name3498 (
		_w110_,
		_w72_,
		_w43_,
		_w3532_
	);
	LUT4 #(
		.INIT('h153f)
	) name3499 (
		_w110_,
		_w43_,
		_w46_,
		_w201_,
		_w3533_
	);
	LUT4 #(
		.INIT('h4000)
	) name3500 (
		_w482_,
		_w3532_,
		_w3533_,
		_w3531_,
		_w3534_
	);
	LUT4 #(
		.INIT('h1000)
	) name3501 (
		_w379_,
		_w473_,
		_w554_,
		_w1356_,
		_w3535_
	);
	LUT3 #(
		.INIT('h80)
	) name3502 (
		_w211_,
		_w619_,
		_w802_,
		_w3536_
	);
	LUT4 #(
		.INIT('h8000)
	) name3503 (
		_w1267_,
		_w3536_,
		_w3534_,
		_w3535_,
		_w3537_
	);
	LUT4 #(
		.INIT('h0777)
	) name3504 (
		_w122_,
		_w55_,
		_w78_,
		_w90_,
		_w3538_
	);
	LUT4 #(
		.INIT('h153f)
	) name3505 (
		_w38_,
		_w85_,
		_w43_,
		_w176_,
		_w3539_
	);
	LUT3 #(
		.INIT('h80)
	) name3506 (
		_w3073_,
		_w3538_,
		_w3539_,
		_w3540_
	);
	LUT2 #(
		.INIT('h8)
	) name3507 (
		_w1964_,
		_w3540_,
		_w3541_
	);
	LUT4 #(
		.INIT('h153f)
	) name3508 (
		_w41_,
		_w65_,
		_w259_,
		_w430_,
		_w3542_
	);
	LUT4 #(
		.INIT('h153f)
	) name3509 (
		_w38_,
		_w93_,
		_w419_,
		_w430_,
		_w3543_
	);
	LUT4 #(
		.INIT('h153f)
	) name3510 (
		_w122_,
		_w106_,
		_w67_,
		_w65_,
		_w3544_
	);
	LUT4 #(
		.INIT('h135f)
	) name3511 (
		_w52_,
		_w59_,
		_w78_,
		_w236_,
		_w3545_
	);
	LUT4 #(
		.INIT('h8000)
	) name3512 (
		_w3544_,
		_w3545_,
		_w3542_,
		_w3543_,
		_w3546_
	);
	LUT2 #(
		.INIT('h8)
	) name3513 (
		_w2670_,
		_w3546_,
		_w3547_
	);
	LUT4 #(
		.INIT('h8000)
	) name3514 (
		_w1964_,
		_w2670_,
		_w3540_,
		_w3546_,
		_w3548_
	);
	LUT4 #(
		.INIT('h135f)
	) name3515 (
		_w55_,
		_w65_,
		_w158_,
		_w419_,
		_w3549_
	);
	LUT2 #(
		.INIT('h8)
	) name3516 (
		_w1359_,
		_w3549_,
		_w3550_
	);
	LUT4 #(
		.INIT('h8000)
	) name3517 (
		_w1013_,
		_w1191_,
		_w1982_,
		_w1983_,
		_w3551_
	);
	LUT3 #(
		.INIT('h80)
	) name3518 (
		_w2118_,
		_w2275_,
		_w2706_,
		_w3552_
	);
	LUT4 #(
		.INIT('h153f)
	) name3519 (
		_w59_,
		_w47_,
		_w43_,
		_w184_,
		_w3553_
	);
	LUT4 #(
		.INIT('h153f)
	) name3520 (
		_w56_,
		_w65_,
		_w166_,
		_w259_,
		_w3554_
	);
	LUT4 #(
		.INIT('h8000)
	) name3521 (
		_w403_,
		_w1067_,
		_w3553_,
		_w3554_,
		_w3555_
	);
	LUT4 #(
		.INIT('h8000)
	) name3522 (
		_w3550_,
		_w3552_,
		_w3555_,
		_w3551_,
		_w3556_
	);
	LUT4 #(
		.INIT('h8000)
	) name3523 (
		_w3171_,
		_w3537_,
		_w3548_,
		_w3556_,
		_w3557_
	);
	LUT2 #(
		.INIT('h8)
	) name3524 (
		_w3530_,
		_w3557_,
		_w3558_
	);
	LUT4 #(
		.INIT('h135f)
	) name3525 (
		_w106_,
		_w78_,
		_w93_,
		_w44_,
		_w3559_
	);
	LUT4 #(
		.INIT('h8000)
	) name3526 (
		_w611_,
		_w908_,
		_w2502_,
		_w3559_,
		_w3560_
	);
	LUT4 #(
		.INIT('h153f)
	) name3527 (
		_w65_,
		_w44_,
		_w176_,
		_w419_,
		_w3561_
	);
	LUT4 #(
		.INIT('h8000)
	) name3528 (
		_w802_,
		_w1079_,
		_w1280_,
		_w3561_,
		_w3562_
	);
	LUT3 #(
		.INIT('h80)
	) name3529 (
		_w2899_,
		_w3560_,
		_w3562_,
		_w3563_
	);
	LUT3 #(
		.INIT('h80)
	) name3530 (
		_w609_,
		_w768_,
		_w2073_,
		_w3564_
	);
	LUT3 #(
		.INIT('h1f)
	) name3531 (
		_w38_,
		_w90_,
		_w378_,
		_w3565_
	);
	LUT4 #(
		.INIT('h135f)
	) name3532 (
		_w67_,
		_w46_,
		_w419_,
		_w430_,
		_w3566_
	);
	LUT3 #(
		.INIT('h37)
	) name3533 (
		_w106_,
		_w110_,
		_w43_,
		_w3567_
	);
	LUT4 #(
		.INIT('h135f)
	) name3534 (
		_w122_,
		_w56_,
		_w46_,
		_w201_,
		_w3568_
	);
	LUT4 #(
		.INIT('h8000)
	) name3535 (
		_w3567_,
		_w3568_,
		_w3565_,
		_w3566_,
		_w3569_
	);
	LUT4 #(
		.INIT('h135f)
	) name3536 (
		_w110_,
		_w90_,
		_w39_,
		_w176_,
		_w3570_
	);
	LUT4 #(
		.INIT('h153f)
	) name3537 (
		_w59_,
		_w44_,
		_w378_,
		_w430_,
		_w3571_
	);
	LUT4 #(
		.INIT('h8000)
	) name3538 (
		_w343_,
		_w660_,
		_w3570_,
		_w3571_,
		_w3572_
	);
	LUT4 #(
		.INIT('h0777)
	) name3539 (
		_w106_,
		_w52_,
		_w93_,
		_w184_,
		_w3573_
	);
	LUT4 #(
		.INIT('h8000)
	) name3540 (
		_w54_,
		_w597_,
		_w598_,
		_w3573_,
		_w3574_
	);
	LUT4 #(
		.INIT('h8000)
	) name3541 (
		_w3564_,
		_w3569_,
		_w3572_,
		_w3574_,
		_w3575_
	);
	LUT2 #(
		.INIT('h8)
	) name3542 (
		_w3563_,
		_w3575_,
		_w3576_
	);
	LUT3 #(
		.INIT('h1f)
	) name3543 (
		_w38_,
		_w55_,
		_w259_,
		_w3577_
	);
	LUT4 #(
		.INIT('h135f)
	) name3544 (
		_w106_,
		_w55_,
		_w44_,
		_w419_,
		_w3578_
	);
	LUT4 #(
		.INIT('h8000)
	) name3545 (
		_w491_,
		_w675_,
		_w3577_,
		_w3578_,
		_w3579_
	);
	LUT4 #(
		.INIT('h8000)
	) name3546 (
		_w809_,
		_w829_,
		_w935_,
		_w2222_,
		_w3580_
	);
	LUT4 #(
		.INIT('h8000)
	) name3547 (
		_w2197_,
		_w2898_,
		_w3580_,
		_w3579_,
		_w3581_
	);
	LUT3 #(
		.INIT('h57)
	) name3548 (
		_w59_,
		_w39_,
		_w43_,
		_w3582_
	);
	LUT4 #(
		.INIT('h0777)
	) name3549 (
		_w90_,
		_w72_,
		_w50_,
		_w236_,
		_w3583_
	);
	LUT2 #(
		.INIT('h8)
	) name3550 (
		_w3582_,
		_w3583_,
		_w3584_
	);
	LUT4 #(
		.INIT('h135f)
	) name3551 (
		_w85_,
		_w46_,
		_w176_,
		_w378_,
		_w3585_
	);
	LUT3 #(
		.INIT('h80)
	) name3552 (
		_w198_,
		_w3158_,
		_w3585_,
		_w3586_
	);
	LUT4 #(
		.INIT('h135f)
	) name3553 (
		_w85_,
		_w90_,
		_w39_,
		_w184_,
		_w3587_
	);
	LUT4 #(
		.INIT('h8000)
	) name3554 (
		_w605_,
		_w1297_,
		_w1625_,
		_w3587_,
		_w3588_
	);
	LUT4 #(
		.INIT('h153f)
	) name3555 (
		_w55_,
		_w56_,
		_w184_,
		_w158_,
		_w3589_
	);
	LUT4 #(
		.INIT('h135f)
	) name3556 (
		_w59_,
		_w110_,
		_w176_,
		_w430_,
		_w3590_
	);
	LUT4 #(
		.INIT('h2000)
	) name3557 (
		_w148_,
		_w325_,
		_w3589_,
		_w3590_,
		_w3591_
	);
	LUT4 #(
		.INIT('h8000)
	) name3558 (
		_w3584_,
		_w3586_,
		_w3588_,
		_w3591_,
		_w3592_
	);
	LUT4 #(
		.INIT('h8000)
	) name3559 (
		_w2916_,
		_w2924_,
		_w3581_,
		_w3592_,
		_w3593_
	);
	LUT2 #(
		.INIT('h8)
	) name3560 (
		_w3576_,
		_w3593_,
		_w3594_
	);
	LUT4 #(
		.INIT('h0777)
	) name3561 (
		_w3530_,
		_w3557_,
		_w3576_,
		_w3593_,
		_w3595_
	);
	LUT4 #(
		.INIT('h8000)
	) name3562 (
		_w3530_,
		_w3557_,
		_w3576_,
		_w3593_,
		_w3596_
	);
	LUT4 #(
		.INIT('h044c)
	) name3563 (
		\a[8] ,
		_w3456_,
		_w3558_,
		_w3594_,
		_w3597_
	);
	LUT4 #(
		.INIT('h3220)
	) name3564 (
		\a[8] ,
		_w3456_,
		_w3558_,
		_w3594_,
		_w3598_
	);
	LUT4 #(
		.INIT('h54ab)
	) name3565 (
		_w1773_,
		_w2315_,
		_w2316_,
		_w2318_,
		_w3599_
	);
	LUT3 #(
		.INIT('h70)
	) name3566 (
		_w1692_,
		_w1723_,
		_w2407_,
		_w3600_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name3567 (
		_w376_,
		_w1751_,
		_w1742_,
		_w1771_,
		_w3601_
	);
	LUT3 #(
		.INIT('h70)
	) name3568 (
		_w1620_,
		_w1661_,
		_w2527_,
		_w3602_
	);
	LUT3 #(
		.INIT('h01)
	) name3569 (
		_w3601_,
		_w3602_,
		_w3600_,
		_w3603_
	);
	LUT4 #(
		.INIT('h2033)
	) name3570 (
		_w377_,
		_w3598_,
		_w3599_,
		_w3603_,
		_w3604_
	);
	LUT4 #(
		.INIT('h4445)
	) name3571 (
		_w3515_,
		_w3516_,
		_w3597_,
		_w3604_,
		_w3605_
	);
	LUT4 #(
		.INIT('h4c00)
	) name3572 (
		_w377_,
		_w3494_,
		_w3495_,
		_w3499_,
		_w3606_
	);
	LUT4 #(
		.INIT('h93cc)
	) name3573 (
		_w377_,
		_w3494_,
		_w3495_,
		_w3499_,
		_w3607_
	);
	LUT3 #(
		.INIT('h54)
	) name3574 (
		_w3500_,
		_w3605_,
		_w3606_,
		_w3608_
	);
	LUT4 #(
		.INIT('h3c39)
	) name3575 (
		\a[11] ,
		_w3139_,
		_w3482_,
		_w3483_,
		_w3609_
	);
	LUT2 #(
		.INIT('h9)
	) name3576 (
		_w3490_,
		_w3609_,
		_w3610_
	);
	LUT2 #(
		.INIT('h4)
	) name3577 (
		_w3608_,
		_w3610_,
		_w3611_
	);
	LUT2 #(
		.INIT('h2)
	) name3578 (
		_w3608_,
		_w3610_,
		_w3612_
	);
	LUT2 #(
		.INIT('h9)
	) name3579 (
		_w3608_,
		_w3610_,
		_w3613_
	);
	LUT3 #(
		.INIT('h70)
	) name3580 (
		_w1381_,
		_w1398_,
		_w2549_,
		_w3614_
	);
	LUT3 #(
		.INIT('h70)
	) name3581 (
		_w1325_,
		_w1367_,
		_w2617_,
		_w3615_
	);
	LUT3 #(
		.INIT('h70)
	) name3582 (
		_w1253_,
		_w1294_,
		_w2854_,
		_w3616_
	);
	LUT3 #(
		.INIT('h01)
	) name3583 (
		_w3615_,
		_w3616_,
		_w3614_,
		_w3617_
	);
	LUT4 #(
		.INIT('h95aa)
	) name3584 (
		\a[29] ,
		_w2550_,
		_w3182_,
		_w3617_,
		_w3618_
	);
	LUT4 #(
		.INIT('h20a2)
	) name3585 (
		_w3493_,
		_w3608_,
		_w3610_,
		_w3618_,
		_w3619_
	);
	LUT4 #(
		.INIT('h222b)
	) name3586 (
		_w3426_,
		_w3427_,
		_w3492_,
		_w3619_,
		_w3620_
	);
	LUT3 #(
		.INIT('h69)
	) name3587 (
		\a[29] ,
		_w3379_,
		_w3384_,
		_w3621_
	);
	LUT2 #(
		.INIT('h4)
	) name3588 (
		_w3620_,
		_w3621_,
		_w3622_
	);
	LUT2 #(
		.INIT('h2)
	) name3589 (
		_w3620_,
		_w3621_,
		_w3623_
	);
	LUT3 #(
		.INIT('h70)
	) name3590 (
		_w1009_,
		_w1050_,
		_w2874_,
		_w3624_
	);
	LUT3 #(
		.INIT('h70)
	) name3591 (
		_w871_,
		_w927_,
		_w2986_,
		_w3625_
	);
	LUT3 #(
		.INIT('h70)
	) name3592 (
		_w763_,
		_w983_,
		_w2975_,
		_w3626_
	);
	LUT3 #(
		.INIT('h01)
	) name3593 (
		_w3625_,
		_w3626_,
		_w3624_,
		_w3627_
	);
	LUT4 #(
		.INIT('h95aa)
	) name3594 (
		\a[26] ,
		_w2839_,
		_w2875_,
		_w3627_,
		_w3628_
	);
	LUT3 #(
		.INIT('h54)
	) name3595 (
		_w3622_,
		_w3623_,
		_w3628_,
		_w3629_
	);
	LUT2 #(
		.INIT('h2)
	) name3596 (
		_w3421_,
		_w3629_,
		_w3630_
	);
	LUT2 #(
		.INIT('h4)
	) name3597 (
		_w3421_,
		_w3629_,
		_w3631_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3598 (
		_w587_,
		_w608_,
		_w624_,
		_w3262_,
		_w3632_
	);
	LUT3 #(
		.INIT('h2a)
	) name3599 (
		_w3214_,
		_w725_,
		_w764_,
		_w3633_
	);
	LUT3 #(
		.INIT('h70)
	) name3600 (
		_w666_,
		_w694_,
		_w3249_,
		_w3634_
	);
	LUT3 #(
		.INIT('h01)
	) name3601 (
		_w3633_,
		_w3634_,
		_w3632_,
		_w3635_
	);
	LUT4 #(
		.INIT('h95aa)
	) name3602 (
		\a[23] ,
		_w2598_,
		_w37_,
		_w3635_,
		_w3636_
	);
	LUT3 #(
		.INIT('h54)
	) name3603 (
		_w3630_,
		_w3631_,
		_w3636_,
		_w3637_
	);
	LUT3 #(
		.INIT('h54)
	) name3604 (
		_w3417_,
		_w3418_,
		_w3637_,
		_w3638_
	);
	LUT2 #(
		.INIT('h9)
	) name3605 (
		_w3394_,
		_w3395_,
		_w3639_
	);
	LUT2 #(
		.INIT('h6)
	) name3606 (
		_w3402_,
		_w3639_,
		_w3640_
	);
	LUT2 #(
		.INIT('h1)
	) name3607 (
		_w3638_,
		_w3640_,
		_w3641_
	);
	LUT2 #(
		.INIT('h8)
	) name3608 (
		_w3638_,
		_w3640_,
		_w3642_
	);
	LUT4 #(
		.INIT('hf400)
	) name3609 (
		_w374_,
		_w2361_,
		_w2404_,
		_w3312_,
		_w3643_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3610 (
		_w121_,
		_w418_,
		_w422_,
		_w3311_,
		_w3644_
	);
	LUT3 #(
		.INIT('h18)
	) name3611 (
		\a[17] ,
		\a[18] ,
		\a[19] ,
		_w3645_
	);
	LUT3 #(
		.INIT('h70)
	) name3612 (
		_w352_,
		_w373_,
		_w3645_,
		_w3646_
	);
	LUT2 #(
		.INIT('h1)
	) name3613 (
		_w3644_,
		_w3646_,
		_w3647_
	);
	LUT3 #(
		.INIT('h9a)
	) name3614 (
		\a[20] ,
		_w3643_,
		_w3647_,
		_w3648_
	);
	LUT3 #(
		.INIT('h54)
	) name3615 (
		_w3641_,
		_w3642_,
		_w3648_,
		_w3649_
	);
	LUT4 #(
		.INIT('h022a)
	) name3616 (
		_w3410_,
		_w3638_,
		_w3640_,
		_w3648_,
		_w3650_
	);
	LUT4 #(
		.INIT('h6665)
	) name3617 (
		_w3410_,
		_w3641_,
		_w3642_,
		_w3648_,
		_w3651_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3618 (
		_w486_,
		_w487_,
		_w509_,
		_w3311_,
		_w3652_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3619 (
		_w121_,
		_w418_,
		_w422_,
		_w3645_,
		_w3653_
	);
	LUT4 #(
		.INIT('h6006)
	) name3620 (
		\a[17] ,
		\a[18] ,
		\a[19] ,
		\a[20] ,
		_w3654_
	);
	LUT3 #(
		.INIT('h70)
	) name3621 (
		_w352_,
		_w373_,
		_w3654_,
		_w3655_
	);
	LUT3 #(
		.INIT('h01)
	) name3622 (
		_w3652_,
		_w3653_,
		_w3655_,
		_w3656_
	);
	LUT4 #(
		.INIT('h95aa)
	) name3623 (
		\a[20] ,
		_w2535_,
		_w3312_,
		_w3656_,
		_w3657_
	);
	LUT2 #(
		.INIT('h9)
	) name3624 (
		_w3421_,
		_w3629_,
		_w3658_
	);
	LUT4 #(
		.INIT('h6669)
	) name3625 (
		_w3426_,
		_w3427_,
		_w3492_,
		_w3619_,
		_w3659_
	);
	LUT3 #(
		.INIT('h70)
	) name3626 (
		_w1071_,
		_w1102_,
		_w2874_,
		_w3660_
	);
	LUT3 #(
		.INIT('h70)
	) name3627 (
		_w763_,
		_w983_,
		_w2986_,
		_w3661_
	);
	LUT3 #(
		.INIT('h70)
	) name3628 (
		_w1009_,
		_w1050_,
		_w2975_,
		_w3662_
	);
	LUT3 #(
		.INIT('h01)
	) name3629 (
		_w3661_,
		_w3662_,
		_w3660_,
		_w3663_
	);
	LUT4 #(
		.INIT('h6f00)
	) name3630 (
		_w2339_,
		_w2341_,
		_w2875_,
		_w3663_,
		_w3664_
	);
	LUT3 #(
		.INIT('h84)
	) name3631 (
		\a[26] ,
		_w3659_,
		_w3664_,
		_w3665_
	);
	LUT3 #(
		.INIT('h12)
	) name3632 (
		\a[26] ,
		_w3659_,
		_w3664_,
		_w3666_
	);
	LUT3 #(
		.INIT('h69)
	) name3633 (
		\a[26] ,
		_w3659_,
		_w3664_,
		_w3667_
	);
	LUT4 #(
		.INIT('h6665)
	) name3634 (
		_w3493_,
		_w3611_,
		_w3612_,
		_w3618_,
		_w3668_
	);
	LUT3 #(
		.INIT('h70)
	) name3635 (
		_w1202_,
		_w1233_,
		_w2854_,
		_w3669_
	);
	LUT3 #(
		.INIT('h70)
	) name3636 (
		_w1325_,
		_w1367_,
		_w2549_,
		_w3670_
	);
	LUT3 #(
		.INIT('h70)
	) name3637 (
		_w1253_,
		_w1294_,
		_w2617_,
		_w3671_
	);
	LUT3 #(
		.INIT('h01)
	) name3638 (
		_w3670_,
		_w3671_,
		_w3669_,
		_w3672_
	);
	LUT4 #(
		.INIT('h6f00)
	) name3639 (
		_w2331_,
		_w2333_,
		_w2550_,
		_w3672_,
		_w3673_
	);
	LUT2 #(
		.INIT('h6)
	) name3640 (
		\a[29] ,
		_w3673_,
		_w3674_
	);
	LUT2 #(
		.INIT('h2)
	) name3641 (
		_w3668_,
		_w3674_,
		_w3675_
	);
	LUT3 #(
		.INIT('h70)
	) name3642 (
		_w1136_,
		_w1187_,
		_w2874_,
		_w3676_
	);
	LUT3 #(
		.INIT('h70)
	) name3643 (
		_w1009_,
		_w1050_,
		_w2986_,
		_w3677_
	);
	LUT3 #(
		.INIT('h70)
	) name3644 (
		_w1071_,
		_w1102_,
		_w2975_,
		_w3678_
	);
	LUT3 #(
		.INIT('h01)
	) name3645 (
		_w3677_,
		_w3678_,
		_w3676_,
		_w3679_
	);
	LUT4 #(
		.INIT('h95aa)
	) name3646 (
		\a[26] ,
		_w2875_,
		_w2936_,
		_w3679_,
		_w3680_
	);
	LUT2 #(
		.INIT('h4)
	) name3647 (
		_w3668_,
		_w3674_,
		_w3681_
	);
	LUT3 #(
		.INIT('h54)
	) name3648 (
		_w3675_,
		_w3680_,
		_w3681_,
		_w3682_
	);
	LUT3 #(
		.INIT('h54)
	) name3649 (
		_w3665_,
		_w3666_,
		_w3682_,
		_w3683_
	);
	LUT2 #(
		.INIT('h9)
	) name3650 (
		_w3620_,
		_w3621_,
		_w3684_
	);
	LUT2 #(
		.INIT('h9)
	) name3651 (
		_w3628_,
		_w3684_,
		_w3685_
	);
	LUT3 #(
		.INIT('h70)
	) name3652 (
		_w725_,
		_w764_,
		_w3249_,
		_w3686_
	);
	LUT3 #(
		.INIT('h2a)
	) name3653 (
		_w3214_,
		_w801_,
		_w851_,
		_w3687_
	);
	LUT3 #(
		.INIT('h70)
	) name3654 (
		_w666_,
		_w694_,
		_w3262_,
		_w3688_
	);
	LUT3 #(
		.INIT('h01)
	) name3655 (
		_w3687_,
		_w3688_,
		_w3686_,
		_w3689_
	);
	LUT4 #(
		.INIT('h6f00)
	) name3656 (
		_w2347_,
		_w2349_,
		_w37_,
		_w3689_,
		_w3690_
	);
	LUT4 #(
		.INIT('h4d8e)
	) name3657 (
		\a[23] ,
		_w3683_,
		_w3685_,
		_w3690_,
		_w3691_
	);
	LUT3 #(
		.INIT('h09)
	) name3658 (
		_w3636_,
		_w3658_,
		_w3691_,
		_w3692_
	);
	LUT3 #(
		.INIT('h60)
	) name3659 (
		_w3636_,
		_w3658_,
		_w3691_,
		_w3693_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3660 (
		_w486_,
		_w487_,
		_w509_,
		_w3645_,
		_w3694_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3661 (
		_w121_,
		_w418_,
		_w422_,
		_w3654_,
		_w3695_
	);
	LUT3 #(
		.INIT('h70)
	) name3662 (
		_w544_,
		_w558_,
		_w3311_,
		_w3696_
	);
	LUT3 #(
		.INIT('h01)
	) name3663 (
		_w3694_,
		_w3695_,
		_w3696_,
		_w3697_
	);
	LUT4 #(
		.INIT('h6f00)
	) name3664 (
		_w2355_,
		_w2357_,
		_w3312_,
		_w3697_,
		_w3698_
	);
	LUT4 #(
		.INIT('h3132)
	) name3665 (
		\a[20] ,
		_w3692_,
		_w3693_,
		_w3698_,
		_w3699_
	);
	LUT2 #(
		.INIT('h9)
	) name3666 (
		_w3419_,
		_w3637_,
		_w3700_
	);
	LUT3 #(
		.INIT('h8e)
	) name3667 (
		_w3657_,
		_w3699_,
		_w3700_,
		_w3701_
	);
	LUT2 #(
		.INIT('h6)
	) name3668 (
		_w3638_,
		_w3640_,
		_w3702_
	);
	LUT2 #(
		.INIT('h9)
	) name3669 (
		_w3648_,
		_w3702_,
		_w3703_
	);
	LUT3 #(
		.INIT('h21)
	) name3670 (
		_w3648_,
		_w3701_,
		_w3702_,
		_w3704_
	);
	LUT3 #(
		.INIT('h48)
	) name3671 (
		_w3648_,
		_w3701_,
		_w3702_,
		_w3705_
	);
	LUT3 #(
		.INIT('h96)
	) name3672 (
		_w3648_,
		_w3701_,
		_w3702_,
		_w3706_
	);
	LUT3 #(
		.INIT('h96)
	) name3673 (
		_w3657_,
		_w3699_,
		_w3700_,
		_w3707_
	);
	LUT2 #(
		.INIT('h9)
	) name3674 (
		\a[14] ,
		\a[15] ,
		_w3708_
	);
	LUT4 #(
		.INIT('h0180)
	) name3675 (
		\a[14] ,
		\a[15] ,
		\a[16] ,
		\a[17] ,
		_w3709_
	);
	LUT4 #(
		.INIT('h0660)
	) name3676 (
		\a[14] ,
		\a[15] ,
		\a[16] ,
		\a[17] ,
		_w3710_
	);
	LUT4 #(
		.INIT('h5150)
	) name3677 (
		_w374_,
		_w2361_,
		_w3709_,
		_w3710_,
		_w3711_
	);
	LUT3 #(
		.INIT('h70)
	) name3678 (
		_w725_,
		_w764_,
		_w3262_,
		_w3712_
	);
	LUT3 #(
		.INIT('h70)
	) name3679 (
		_w801_,
		_w851_,
		_w3249_,
		_w3713_
	);
	LUT3 #(
		.INIT('h2a)
	) name3680 (
		_w3214_,
		_w871_,
		_w927_,
		_w3714_
	);
	LUT3 #(
		.INIT('h01)
	) name3681 (
		_w3713_,
		_w3714_,
		_w3712_,
		_w3715_
	);
	LUT4 #(
		.INIT('h95aa)
	) name3682 (
		\a[23] ,
		_w2724_,
		_w37_,
		_w3715_,
		_w3716_
	);
	LUT2 #(
		.INIT('h9)
	) name3683 (
		_w3667_,
		_w3682_,
		_w3717_
	);
	LUT2 #(
		.INIT('h9)
	) name3684 (
		_w3668_,
		_w3674_,
		_w3718_
	);
	LUT2 #(
		.INIT('h9)
	) name3685 (
		_w3613_,
		_w3618_,
		_w3719_
	);
	LUT3 #(
		.INIT('h56)
	) name3686 (
		_w3517_,
		_w3597_,
		_w3604_,
		_w3720_
	);
	LUT3 #(
		.INIT('h2a)
	) name3687 (
		_w376_,
		_w1692_,
		_w1723_,
		_w3721_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3688 (
		_w1584_,
		_w1569_,
		_w1606_,
		_w2527_,
		_w3722_
	);
	LUT3 #(
		.INIT('h70)
	) name3689 (
		_w1620_,
		_w1661_,
		_w2407_,
		_w3723_
	);
	LUT3 #(
		.INIT('h01)
	) name3690 (
		_w3722_,
		_w3723_,
		_w3721_,
		_w3724_
	);
	LUT4 #(
		.INIT('h7d00)
	) name3691 (
		_w377_,
		_w2319_,
		_w2321_,
		_w3724_,
		_w3725_
	);
	LUT4 #(
		.INIT('h0056)
	) name3692 (
		_w3517_,
		_w3597_,
		_w3604_,
		_w3725_,
		_w3726_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3693 (
		_w1454_,
		_w1426_,
		_w1478_,
		_w2617_,
		_w3727_
	);
	LUT3 #(
		.INIT('h70)
	) name3694 (
		_w1381_,
		_w1398_,
		_w2854_,
		_w3728_
	);
	LUT3 #(
		.INIT('h70)
	) name3695 (
		_w1501_,
		_w1545_,
		_w2549_,
		_w3729_
	);
	LUT3 #(
		.INIT('h01)
	) name3696 (
		_w3728_,
		_w3729_,
		_w3727_,
		_w3730_
	);
	LUT4 #(
		.INIT('h95aa)
	) name3697 (
		\a[29] ,
		_w2550_,
		_w3362_,
		_w3730_,
		_w3731_
	);
	LUT4 #(
		.INIT('ha900)
	) name3698 (
		_w3517_,
		_w3597_,
		_w3604_,
		_w3725_,
		_w3732_
	);
	LUT4 #(
		.INIT('h56a9)
	) name3699 (
		_w3517_,
		_w3597_,
		_w3604_,
		_w3725_,
		_w3733_
	);
	LUT2 #(
		.INIT('h9)
	) name3700 (
		_w3605_,
		_w3607_,
		_w3734_
	);
	LUT4 #(
		.INIT('h2b00)
	) name3701 (
		_w3720_,
		_w3725_,
		_w3731_,
		_w3734_,
		_w3735_
	);
	LUT4 #(
		.INIT('h00d4)
	) name3702 (
		_w3720_,
		_w3725_,
		_w3731_,
		_w3734_,
		_w3736_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3703 (
		_w1454_,
		_w1426_,
		_w1478_,
		_w2549_,
		_w3737_
	);
	LUT3 #(
		.INIT('h70)
	) name3704 (
		_w1325_,
		_w1367_,
		_w2854_,
		_w3738_
	);
	LUT3 #(
		.INIT('h70)
	) name3705 (
		_w1381_,
		_w1398_,
		_w2617_,
		_w3739_
	);
	LUT3 #(
		.INIT('h01)
	) name3706 (
		_w3738_,
		_w3739_,
		_w3737_,
		_w3740_
	);
	LUT4 #(
		.INIT('h6f00)
	) name3707 (
		_w2327_,
		_w2329_,
		_w2550_,
		_w3740_,
		_w3741_
	);
	LUT2 #(
		.INIT('h6)
	) name3708 (
		\a[29] ,
		_w3741_,
		_w3742_
	);
	LUT3 #(
		.INIT('h54)
	) name3709 (
		_w3735_,
		_w3736_,
		_w3742_,
		_w3743_
	);
	LUT3 #(
		.INIT('h70)
	) name3710 (
		_w1136_,
		_w1187_,
		_w2975_,
		_w3744_
	);
	LUT3 #(
		.INIT('h70)
	) name3711 (
		_w1071_,
		_w1102_,
		_w2986_,
		_w3745_
	);
	LUT3 #(
		.INIT('h70)
	) name3712 (
		_w1202_,
		_w1233_,
		_w2874_,
		_w3746_
	);
	LUT3 #(
		.INIT('h01)
	) name3713 (
		_w3745_,
		_w3746_,
		_w3744_,
		_w3747_
	);
	LUT4 #(
		.INIT('h6f00)
	) name3714 (
		_w2335_,
		_w2337_,
		_w2875_,
		_w3747_,
		_w3748_
	);
	LUT4 #(
		.INIT('h71b2)
	) name3715 (
		\a[26] ,
		_w3719_,
		_w3743_,
		_w3748_,
		_w3749_
	);
	LUT3 #(
		.INIT('h09)
	) name3716 (
		_w3680_,
		_w3718_,
		_w3749_,
		_w3750_
	);
	LUT3 #(
		.INIT('h60)
	) name3717 (
		_w3680_,
		_w3718_,
		_w3749_,
		_w3751_
	);
	LUT3 #(
		.INIT('h2a)
	) name3718 (
		_w3214_,
		_w763_,
		_w983_,
		_w3752_
	);
	LUT3 #(
		.INIT('h70)
	) name3719 (
		_w871_,
		_w927_,
		_w3249_,
		_w3753_
	);
	LUT3 #(
		.INIT('h70)
	) name3720 (
		_w801_,
		_w851_,
		_w3262_,
		_w3754_
	);
	LUT3 #(
		.INIT('h01)
	) name3721 (
		_w3753_,
		_w3754_,
		_w3752_,
		_w3755_
	);
	LUT4 #(
		.INIT('h6f00)
	) name3722 (
		_w2343_,
		_w2345_,
		_w37_,
		_w3755_,
		_w3756_
	);
	LUT4 #(
		.INIT('h3132)
	) name3723 (
		\a[23] ,
		_w3750_,
		_w3751_,
		_w3756_,
		_w3757_
	);
	LUT3 #(
		.INIT('hb2)
	) name3724 (
		_w3716_,
		_w3717_,
		_w3757_,
		_w3758_
	);
	LUT4 #(
		.INIT('h9669)
	) name3725 (
		\a[23] ,
		_w3683_,
		_w3685_,
		_w3690_,
		_w3759_
	);
	LUT2 #(
		.INIT('h1)
	) name3726 (
		_w3758_,
		_w3759_,
		_w3760_
	);
	LUT2 #(
		.INIT('h8)
	) name3727 (
		_w3758_,
		_w3759_,
		_w3761_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3728 (
		_w486_,
		_w487_,
		_w509_,
		_w3654_,
		_w3762_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3729 (
		_w587_,
		_w608_,
		_w624_,
		_w3311_,
		_w3763_
	);
	LUT3 #(
		.INIT('h70)
	) name3730 (
		_w544_,
		_w558_,
		_w3645_,
		_w3764_
	);
	LUT3 #(
		.INIT('h01)
	) name3731 (
		_w3762_,
		_w3763_,
		_w3764_,
		_w3765_
	);
	LUT4 #(
		.INIT('h95aa)
	) name3732 (
		\a[20] ,
		_w2526_,
		_w3312_,
		_w3765_,
		_w3766_
	);
	LUT3 #(
		.INIT('h54)
	) name3733 (
		_w3760_,
		_w3761_,
		_w3766_,
		_w3767_
	);
	LUT3 #(
		.INIT('h96)
	) name3734 (
		_w3636_,
		_w3658_,
		_w3691_,
		_w3768_
	);
	LUT3 #(
		.INIT('h69)
	) name3735 (
		\a[20] ,
		_w3698_,
		_w3768_,
		_w3769_
	);
	LUT4 #(
		.INIT('h90f9)
	) name3736 (
		\a[17] ,
		_w3711_,
		_w3767_,
		_w3769_,
		_w3770_
	);
	LUT2 #(
		.INIT('h2)
	) name3737 (
		_w3707_,
		_w3770_,
		_w3771_
	);
	LUT4 #(
		.INIT('h9669)
	) name3738 (
		\a[17] ,
		_w3711_,
		_w3767_,
		_w3769_,
		_w3772_
	);
	LUT3 #(
		.INIT('h96)
	) name3739 (
		_w3716_,
		_w3717_,
		_w3757_,
		_w3773_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3740 (
		_w587_,
		_w608_,
		_w624_,
		_w3645_,
		_w3774_
	);
	LUT3 #(
		.INIT('h70)
	) name3741 (
		_w666_,
		_w694_,
		_w3311_,
		_w3775_
	);
	LUT3 #(
		.INIT('h70)
	) name3742 (
		_w544_,
		_w558_,
		_w3654_,
		_w3776_
	);
	LUT3 #(
		.INIT('h01)
	) name3743 (
		_w3775_,
		_w3776_,
		_w3774_,
		_w3777_
	);
	LUT4 #(
		.INIT('h6f00)
	) name3744 (
		_w2351_,
		_w2353_,
		_w3312_,
		_w3777_,
		_w3778_
	);
	LUT3 #(
		.INIT('h84)
	) name3745 (
		\a[20] ,
		_w3773_,
		_w3778_,
		_w3779_
	);
	LUT3 #(
		.INIT('h12)
	) name3746 (
		\a[20] ,
		_w3773_,
		_w3778_,
		_w3780_
	);
	LUT3 #(
		.INIT('h69)
	) name3747 (
		\a[20] ,
		_w3773_,
		_w3778_,
		_w3781_
	);
	LUT3 #(
		.INIT('h96)
	) name3748 (
		_w3680_,
		_w3718_,
		_w3749_,
		_w3782_
	);
	LUT3 #(
		.INIT('h69)
	) name3749 (
		\a[23] ,
		_w3756_,
		_w3782_,
		_w3783_
	);
	LUT3 #(
		.INIT('h70)
	) name3750 (
		_w1202_,
		_w1233_,
		_w2975_,
		_w3784_
	);
	LUT3 #(
		.INIT('h70)
	) name3751 (
		_w1253_,
		_w1294_,
		_w2874_,
		_w3785_
	);
	LUT3 #(
		.INIT('h70)
	) name3752 (
		_w1136_,
		_w1187_,
		_w2986_,
		_w3786_
	);
	LUT3 #(
		.INIT('h01)
	) name3753 (
		_w3785_,
		_w3786_,
		_w3784_,
		_w3787_
	);
	LUT4 #(
		.INIT('h95aa)
	) name3754 (
		\a[26] ,
		_w2875_,
		_w3067_,
		_w3787_,
		_w3788_
	);
	LUT4 #(
		.INIT('h54ab)
	) name3755 (
		_w3726_,
		_w3731_,
		_w3732_,
		_w3734_,
		_w3789_
	);
	LUT2 #(
		.INIT('h9)
	) name3756 (
		_w3742_,
		_w3789_,
		_w3790_
	);
	LUT3 #(
		.INIT('h57)
	) name3757 (
		_w55_,
		_w158_,
		_w378_,
		_w3791_
	);
	LUT2 #(
		.INIT('h4)
	) name3758 (
		_w462_,
		_w3791_,
		_w3792_
	);
	LUT4 #(
		.INIT('h135f)
	) name3759 (
		_w122_,
		_w52_,
		_w47_,
		_w201_,
		_w3793_
	);
	LUT4 #(
		.INIT('h135f)
	) name3760 (
		_w90_,
		_w41_,
		_w158_,
		_w259_,
		_w3794_
	);
	LUT4 #(
		.INIT('h8000)
	) name3761 (
		_w806_,
		_w950_,
		_w3793_,
		_w3794_,
		_w3795_
	);
	LUT3 #(
		.INIT('h57)
	) name3762 (
		_w78_,
		_w56_,
		_w65_,
		_w3796_
	);
	LUT4 #(
		.INIT('h8000)
	) name3763 (
		_w1061_,
		_w1196_,
		_w3088_,
		_w3796_,
		_w3797_
	);
	LUT4 #(
		.INIT('h8000)
	) name3764 (
		_w3560_,
		_w3792_,
		_w3797_,
		_w3795_,
		_w3798_
	);
	LUT3 #(
		.INIT('h37)
	) name3765 (
		_w122_,
		_w110_,
		_w176_,
		_w3799_
	);
	LUT4 #(
		.INIT('h4000)
	) name3766 (
		_w451_,
		_w720_,
		_w721_,
		_w3799_,
		_w3800_
	);
	LUT4 #(
		.INIT('h4000)
	) name3767 (
		_w142_,
		_w1281_,
		_w1514_,
		_w2649_,
		_w3801_
	);
	LUT3 #(
		.INIT('h20)
	) name3768 (
		_w68_,
		_w334_,
		_w843_,
		_w3802_
	);
	LUT4 #(
		.INIT('h8000)
	) name3769 (
		_w1372_,
		_w1480_,
		_w2809_,
		_w3561_,
		_w3803_
	);
	LUT4 #(
		.INIT('h8000)
	) name3770 (
		_w3802_,
		_w3803_,
		_w3800_,
		_w3801_,
		_w3804_
	);
	LUT4 #(
		.INIT('h8000)
	) name3771 (
		_w1146_,
		_w3527_,
		_w3804_,
		_w3798_,
		_w3805_
	);
	LUT2 #(
		.INIT('h8)
	) name3772 (
		_w2800_,
		_w3805_,
		_w3806_
	);
	LUT4 #(
		.INIT('h153f)
	) name3773 (
		_w110_,
		_w50_,
		_w259_,
		_w378_,
		_w3807_
	);
	LUT4 #(
		.INIT('h0777)
	) name3774 (
		_w106_,
		_w59_,
		_w43_,
		_w46_,
		_w3808_
	);
	LUT4 #(
		.INIT('h4000)
	) name3775 (
		_w478_,
		_w555_,
		_w3808_,
		_w3807_,
		_w3809_
	);
	LUT4 #(
		.INIT('h1000)
	) name3776 (
		_w295_,
		_w407_,
		_w951_,
		_w2570_,
		_w3810_
	);
	LUT4 #(
		.INIT('h135f)
	) name3777 (
		_w65_,
		_w46_,
		_w236_,
		_w259_,
		_w3811_
	);
	LUT3 #(
		.INIT('h80)
	) name3778 (
		_w834_,
		_w2561_,
		_w3811_,
		_w3812_
	);
	LUT4 #(
		.INIT('h8000)
	) name3779 (
		_w911_,
		_w3812_,
		_w3809_,
		_w3810_,
		_w3813_
	);
	LUT4 #(
		.INIT('h135f)
	) name3780 (
		_w85_,
		_w78_,
		_w72_,
		_w46_,
		_w3814_
	);
	LUT2 #(
		.INIT('h4)
	) name3781 (
		_w458_,
		_w3814_,
		_w3815_
	);
	LUT3 #(
		.INIT('h80)
	) name3782 (
		_w844_,
		_w1562_,
		_w1585_,
		_w3816_
	);
	LUT4 #(
		.INIT('h8000)
	) name3783 (
		_w875_,
		_w880_,
		_w3815_,
		_w3816_,
		_w3817_
	);
	LUT4 #(
		.INIT('h8000)
	) name3784 (
		_w2456_,
		_w2464_,
		_w3813_,
		_w3817_,
		_w3818_
	);
	LUT4 #(
		.INIT('he888)
	) name3785 (
		\a[2] ,
		\a[5] ,
		_w3151_,
		_w3818_,
		_w3819_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3786 (
		_w1817_,
		_w1799_,
		_w1840_,
		_w2407_,
		_w3820_
	);
	LUT3 #(
		.INIT('h70)
	) name3787 (
		_w1795_,
		_w1796_,
		_w2527_,
		_w3821_
	);
	LUT3 #(
		.INIT('h2a)
	) name3788 (
		_w376_,
		_w1863_,
		_w1875_,
		_w3822_
	);
	LUT3 #(
		.INIT('h01)
	) name3789 (
		_w3821_,
		_w3822_,
		_w3820_,
		_w3823_
	);
	LUT4 #(
		.INIT('h7d00)
	) name3790 (
		_w377_,
		_w2311_,
		_w2313_,
		_w3823_,
		_w3824_
	);
	LUT4 #(
		.INIT('hd554)
	) name3791 (
		_w3558_,
		_w3806_,
		_w3819_,
		_w3824_,
		_w3825_
	);
	LUT3 #(
		.INIT('ha9)
	) name3792 (
		\a[8] ,
		_w3595_,
		_w3596_,
		_w3826_
	);
	LUT3 #(
		.INIT('h70)
	) name3793 (
		_w1692_,
		_w1723_,
		_w2527_,
		_w3827_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3794 (
		_w1751_,
		_w1742_,
		_w1771_,
		_w2407_,
		_w3828_
	);
	LUT3 #(
		.INIT('h2a)
	) name3795 (
		_w376_,
		_w1795_,
		_w1796_,
		_w3829_
	);
	LUT3 #(
		.INIT('h01)
	) name3796 (
		_w3828_,
		_w3829_,
		_w3827_,
		_w3830_
	);
	LUT4 #(
		.INIT('h7d00)
	) name3797 (
		_w377_,
		_w2315_,
		_w2317_,
		_w3830_,
		_w3831_
	);
	LUT3 #(
		.INIT('he8)
	) name3798 (
		_w3825_,
		_w3826_,
		_w3831_,
		_w3832_
	);
	LUT4 #(
		.INIT('h3c39)
	) name3799 (
		\a[8] ,
		_w3456_,
		_w3595_,
		_w3596_,
		_w3833_
	);
	LUT4 #(
		.INIT('h708f)
	) name3800 (
		_w377_,
		_w3599_,
		_w3603_,
		_w3833_,
		_w3834_
	);
	LUT2 #(
		.INIT('h4)
	) name3801 (
		_w3832_,
		_w3834_,
		_w3835_
	);
	LUT2 #(
		.INIT('h2)
	) name3802 (
		_w3832_,
		_w3834_,
		_w3836_
	);
	LUT2 #(
		.INIT('h9)
	) name3803 (
		_w3832_,
		_w3834_,
		_w3837_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3804 (
		_w1454_,
		_w1426_,
		_w1478_,
		_w2854_,
		_w3838_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3805 (
		_w1584_,
		_w1569_,
		_w1606_,
		_w2549_,
		_w3839_
	);
	LUT3 #(
		.INIT('h70)
	) name3806 (
		_w1501_,
		_w1545_,
		_w2617_,
		_w3840_
	);
	LUT3 #(
		.INIT('h01)
	) name3807 (
		_w3839_,
		_w3840_,
		_w3838_,
		_w3841_
	);
	LUT4 #(
		.INIT('h6f00)
	) name3808 (
		_w2323_,
		_w2325_,
		_w2550_,
		_w3841_,
		_w3842_
	);
	LUT4 #(
		.INIT('h3132)
	) name3809 (
		\a[29] ,
		_w3835_,
		_w3836_,
		_w3842_,
		_w3843_
	);
	LUT3 #(
		.INIT('h09)
	) name3810 (
		_w3731_,
		_w3733_,
		_w3843_,
		_w3844_
	);
	LUT3 #(
		.INIT('h60)
	) name3811 (
		_w3731_,
		_w3733_,
		_w3843_,
		_w3845_
	);
	LUT3 #(
		.INIT('h70)
	) name3812 (
		_w1202_,
		_w1233_,
		_w2986_,
		_w3846_
	);
	LUT3 #(
		.INIT('h70)
	) name3813 (
		_w1325_,
		_w1367_,
		_w2874_,
		_w3847_
	);
	LUT3 #(
		.INIT('h70)
	) name3814 (
		_w1253_,
		_w1294_,
		_w2975_,
		_w3848_
	);
	LUT3 #(
		.INIT('h01)
	) name3815 (
		_w3847_,
		_w3848_,
		_w3846_,
		_w3849_
	);
	LUT4 #(
		.INIT('h6f00)
	) name3816 (
		_w2331_,
		_w2333_,
		_w2875_,
		_w3849_,
		_w3850_
	);
	LUT4 #(
		.INIT('h3132)
	) name3817 (
		\a[26] ,
		_w3844_,
		_w3845_,
		_w3850_,
		_w3851_
	);
	LUT3 #(
		.INIT('hb2)
	) name3818 (
		_w3788_,
		_w3790_,
		_w3851_,
		_w3852_
	);
	LUT4 #(
		.INIT('h6996)
	) name3819 (
		\a[26] ,
		_w3719_,
		_w3743_,
		_w3748_,
		_w3853_
	);
	LUT2 #(
		.INIT('h4)
	) name3820 (
		_w3852_,
		_w3853_,
		_w3854_
	);
	LUT2 #(
		.INIT('h2)
	) name3821 (
		_w3852_,
		_w3853_,
		_w3855_
	);
	LUT3 #(
		.INIT('h2a)
	) name3822 (
		_w3214_,
		_w1009_,
		_w1050_,
		_w3856_
	);
	LUT3 #(
		.INIT('h70)
	) name3823 (
		_w871_,
		_w927_,
		_w3262_,
		_w3857_
	);
	LUT3 #(
		.INIT('h70)
	) name3824 (
		_w763_,
		_w983_,
		_w3249_,
		_w3858_
	);
	LUT3 #(
		.INIT('h01)
	) name3825 (
		_w3857_,
		_w3858_,
		_w3856_,
		_w3859_
	);
	LUT4 #(
		.INIT('h95aa)
	) name3826 (
		\a[23] ,
		_w2839_,
		_w37_,
		_w3859_,
		_w3860_
	);
	LUT3 #(
		.INIT('h54)
	) name3827 (
		_w3854_,
		_w3855_,
		_w3860_,
		_w3861_
	);
	LUT2 #(
		.INIT('h2)
	) name3828 (
		_w3783_,
		_w3861_,
		_w3862_
	);
	LUT2 #(
		.INIT('h4)
	) name3829 (
		_w3783_,
		_w3861_,
		_w3863_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3830 (
		_w587_,
		_w608_,
		_w624_,
		_w3654_,
		_w3864_
	);
	LUT3 #(
		.INIT('h70)
	) name3831 (
		_w725_,
		_w764_,
		_w3311_,
		_w3865_
	);
	LUT3 #(
		.INIT('h70)
	) name3832 (
		_w666_,
		_w694_,
		_w3645_,
		_w3866_
	);
	LUT3 #(
		.INIT('h01)
	) name3833 (
		_w3865_,
		_w3866_,
		_w3864_,
		_w3867_
	);
	LUT4 #(
		.INIT('h95aa)
	) name3834 (
		\a[20] ,
		_w2598_,
		_w3312_,
		_w3867_,
		_w3868_
	);
	LUT3 #(
		.INIT('h54)
	) name3835 (
		_w3862_,
		_w3863_,
		_w3868_,
		_w3869_
	);
	LUT3 #(
		.INIT('h54)
	) name3836 (
		_w3779_,
		_w3780_,
		_w3869_,
		_w3870_
	);
	LUT2 #(
		.INIT('h6)
	) name3837 (
		_w3758_,
		_w3759_,
		_w3871_
	);
	LUT2 #(
		.INIT('h9)
	) name3838 (
		_w3766_,
		_w3871_,
		_w3872_
	);
	LUT2 #(
		.INIT('h4)
	) name3839 (
		_w3870_,
		_w3872_,
		_w3873_
	);
	LUT2 #(
		.INIT('h2)
	) name3840 (
		_w3870_,
		_w3872_,
		_w3874_
	);
	LUT4 #(
		.INIT('hf400)
	) name3841 (
		_w374_,
		_w2361_,
		_w2404_,
		_w3710_,
		_w3875_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3842 (
		_w121_,
		_w418_,
		_w422_,
		_w3709_,
		_w3876_
	);
	LUT3 #(
		.INIT('h18)
	) name3843 (
		\a[14] ,
		\a[15] ,
		\a[16] ,
		_w3877_
	);
	LUT3 #(
		.INIT('h70)
	) name3844 (
		_w352_,
		_w373_,
		_w3877_,
		_w3878_
	);
	LUT2 #(
		.INIT('h1)
	) name3845 (
		_w3876_,
		_w3878_,
		_w3879_
	);
	LUT3 #(
		.INIT('h9a)
	) name3846 (
		\a[17] ,
		_w3875_,
		_w3879_,
		_w3880_
	);
	LUT3 #(
		.INIT('h54)
	) name3847 (
		_w3873_,
		_w3874_,
		_w3880_,
		_w3881_
	);
	LUT4 #(
		.INIT('h20a2)
	) name3848 (
		_w3772_,
		_w3870_,
		_w3872_,
		_w3880_,
		_w3882_
	);
	LUT4 #(
		.INIT('h6665)
	) name3849 (
		_w3772_,
		_w3873_,
		_w3874_,
		_w3880_,
		_w3883_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3850 (
		_w486_,
		_w487_,
		_w509_,
		_w3709_,
		_w3884_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3851 (
		_w121_,
		_w418_,
		_w422_,
		_w3877_,
		_w3885_
	);
	LUT4 #(
		.INIT('h6006)
	) name3852 (
		\a[14] ,
		\a[15] ,
		\a[16] ,
		\a[17] ,
		_w3886_
	);
	LUT3 #(
		.INIT('h70)
	) name3853 (
		_w352_,
		_w373_,
		_w3886_,
		_w3887_
	);
	LUT3 #(
		.INIT('h01)
	) name3854 (
		_w3884_,
		_w3885_,
		_w3887_,
		_w3888_
	);
	LUT4 #(
		.INIT('h95aa)
	) name3855 (
		\a[17] ,
		_w2535_,
		_w3710_,
		_w3888_,
		_w3889_
	);
	LUT2 #(
		.INIT('h9)
	) name3856 (
		_w3783_,
		_w3861_,
		_w3890_
	);
	LUT3 #(
		.INIT('h2a)
	) name3857 (
		_w3214_,
		_w1071_,
		_w1102_,
		_w3891_
	);
	LUT3 #(
		.INIT('h70)
	) name3858 (
		_w763_,
		_w983_,
		_w3262_,
		_w3892_
	);
	LUT3 #(
		.INIT('h70)
	) name3859 (
		_w1009_,
		_w1050_,
		_w3249_,
		_w3893_
	);
	LUT3 #(
		.INIT('h01)
	) name3860 (
		_w3892_,
		_w3893_,
		_w3891_,
		_w3894_
	);
	LUT4 #(
		.INIT('h6f00)
	) name3861 (
		_w2339_,
		_w2341_,
		_w37_,
		_w3894_,
		_w3895_
	);
	LUT3 #(
		.INIT('h96)
	) name3862 (
		_w3788_,
		_w3790_,
		_w3851_,
		_w3896_
	);
	LUT3 #(
		.INIT('h90)
	) name3863 (
		\a[23] ,
		_w3895_,
		_w3896_,
		_w3897_
	);
	LUT3 #(
		.INIT('h06)
	) name3864 (
		\a[23] ,
		_w3895_,
		_w3896_,
		_w3898_
	);
	LUT3 #(
		.INIT('h69)
	) name3865 (
		\a[23] ,
		_w3895_,
		_w3896_,
		_w3899_
	);
	LUT3 #(
		.INIT('h96)
	) name3866 (
		_w3731_,
		_w3733_,
		_w3843_,
		_w3900_
	);
	LUT3 #(
		.INIT('h69)
	) name3867 (
		\a[26] ,
		_w3850_,
		_w3900_,
		_w3901_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3868 (
		_w1584_,
		_w1569_,
		_w1606_,
		_w2617_,
		_w3902_
	);
	LUT3 #(
		.INIT('h70)
	) name3869 (
		_w1501_,
		_w1545_,
		_w2854_,
		_w3903_
	);
	LUT3 #(
		.INIT('h70)
	) name3870 (
		_w1620_,
		_w1661_,
		_w2549_,
		_w3904_
	);
	LUT3 #(
		.INIT('h01)
	) name3871 (
		_w3902_,
		_w3903_,
		_w3904_,
		_w3905_
	);
	LUT4 #(
		.INIT('h95aa)
	) name3872 (
		\a[29] ,
		_w2550_,
		_w3495_,
		_w3905_,
		_w3906_
	);
	LUT3 #(
		.INIT('h69)
	) name3873 (
		_w3825_,
		_w3826_,
		_w3831_,
		_w3907_
	);
	LUT4 #(
		.INIT('h9336)
	) name3874 (
		_w3558_,
		_w3806_,
		_w3819_,
		_w3824_,
		_w3908_
	);
	LUT4 #(
		.INIT('h54ab)
	) name3875 (
		_w1842_,
		_w2311_,
		_w2312_,
		_w2314_,
		_w3909_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3876 (
		_w1751_,
		_w1742_,
		_w1771_,
		_w2527_,
		_w3910_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name3877 (
		_w376_,
		_w1817_,
		_w1799_,
		_w1840_,
		_w3911_
	);
	LUT3 #(
		.INIT('h70)
	) name3878 (
		_w1795_,
		_w1796_,
		_w2407_,
		_w3912_
	);
	LUT3 #(
		.INIT('h01)
	) name3879 (
		_w3911_,
		_w3912_,
		_w3910_,
		_w3913_
	);
	LUT3 #(
		.INIT('h70)
	) name3880 (
		_w377_,
		_w3909_,
		_w3913_,
		_w3914_
	);
	LUT2 #(
		.INIT('h2)
	) name3881 (
		_w3908_,
		_w3914_,
		_w3915_
	);
	LUT2 #(
		.INIT('h9)
	) name3882 (
		_w3558_,
		_w3819_,
		_w3916_
	);
	LUT2 #(
		.INIT('h9)
	) name3883 (
		_w3824_,
		_w3916_,
		_w3917_
	);
	LUT4 #(
		.INIT('h153f)
	) name3884 (
		_w47_,
		_w93_,
		_w176_,
		_w378_,
		_w3918_
	);
	LUT4 #(
		.INIT('h4000)
	) name3885 (
		_w396_,
		_w673_,
		_w1905_,
		_w3918_,
		_w3919_
	);
	LUT3 #(
		.INIT('h80)
	) name3886 (
		_w2468_,
		_w2576_,
		_w3134_,
		_w3920_
	);
	LUT3 #(
		.INIT('h80)
	) name3887 (
		_w1327_,
		_w3919_,
		_w3920_,
		_w3921_
	);
	LUT4 #(
		.INIT('h153f)
	) name3888 (
		_w55_,
		_w85_,
		_w78_,
		_w236_,
		_w3922_
	);
	LUT2 #(
		.INIT('h4)
	) name3889 (
		_w412_,
		_w3922_,
		_w3923_
	);
	LUT4 #(
		.INIT('h8000)
	) name3890 (
		_w87_,
		_w583_,
		_w714_,
		_w2282_,
		_w3924_
	);
	LUT4 #(
		.INIT('h0777)
	) name3891 (
		_w106_,
		_w59_,
		_w72_,
		_w50_,
		_w3925_
	);
	LUT4 #(
		.INIT('h2000)
	) name3892 (
		_w479_,
		_w439_,
		_w832_,
		_w3925_,
		_w3926_
	);
	LUT4 #(
		.INIT('h8000)
	) name3893 (
		_w1427_,
		_w3459_,
		_w3460_,
		_w3503_,
		_w3927_
	);
	LUT4 #(
		.INIT('h8000)
	) name3894 (
		_w3923_,
		_w3924_,
		_w3926_,
		_w3927_,
		_w3928_
	);
	LUT3 #(
		.INIT('h80)
	) name3895 (
		_w328_,
		_w3921_,
		_w3928_,
		_w3929_
	);
	LUT4 #(
		.INIT('h8000)
	) name3896 (
		_w1918_,
		_w1927_,
		_w2062_,
		_w2075_,
		_w3930_
	);
	LUT2 #(
		.INIT('h8)
	) name3897 (
		_w3929_,
		_w3930_,
		_w3931_
	);
	LUT4 #(
		.INIT('h135f)
	) name3898 (
		_w122_,
		_w67_,
		_w56_,
		_w72_,
		_w3932_
	);
	LUT3 #(
		.INIT('h80)
	) name3899 (
		_w2669_,
		_w3336_,
		_w3932_,
		_w3933_
	);
	LUT2 #(
		.INIT('h4)
	) name3900 (
		_w478_,
		_w1091_,
		_w3934_
	);
	LUT4 #(
		.INIT('h1000)
	) name3901 (
		_w477_,
		_w478_,
		_w1091_,
		_w2625_,
		_w3935_
	);
	LUT4 #(
		.INIT('h8000)
	) name3902 (
		_w862_,
		_w3100_,
		_w3935_,
		_w3933_,
		_w3936_
	);
	LUT4 #(
		.INIT('h0777)
	) name3903 (
		_w43_,
		_w93_,
		_w44_,
		_w201_,
		_w3937_
	);
	LUT4 #(
		.INIT('h0777)
	) name3904 (
		_w122_,
		_w41_,
		_w50_,
		_w259_,
		_w3938_
	);
	LUT4 #(
		.INIT('h8000)
	) name3905 (
		_w265_,
		_w1506_,
		_w3937_,
		_w3938_,
		_w3939_
	);
	LUT3 #(
		.INIT('h80)
	) name3906 (
		_w752_,
		_w997_,
		_w1438_,
		_w3940_
	);
	LUT4 #(
		.INIT('h8000)
	) name3907 (
		_w2473_,
		_w2476_,
		_w3939_,
		_w3940_,
		_w3941_
	);
	LUT3 #(
		.INIT('h80)
	) name3908 (
		_w968_,
		_w3936_,
		_w3941_,
		_w3942_
	);
	LUT2 #(
		.INIT('h8)
	) name3909 (
		_w2183_,
		_w3942_,
		_w3943_
	);
	LUT4 #(
		.INIT('h1000)
	) name3910 (
		_w353_,
		_w439_,
		_w832_,
		_w1810_,
		_w3944_
	);
	LUT2 #(
		.INIT('h8)
	) name3911 (
		_w3505_,
		_w3944_,
		_w3945_
	);
	LUT4 #(
		.INIT('h8000)
	) name3912 (
		_w384_,
		_w804_,
		_w1785_,
		_w2118_,
		_w3946_
	);
	LUT3 #(
		.INIT('h57)
	) name3913 (
		_w67_,
		_w201_,
		_w158_,
		_w3947_
	);
	LUT4 #(
		.INIT('h0777)
	) name3914 (
		_w90_,
		_w43_,
		_w93_,
		_w236_,
		_w3948_
	);
	LUT4 #(
		.INIT('h2000)
	) name3915 (
		_w370_,
		_w386_,
		_w3948_,
		_w3947_,
		_w3949_
	);
	LUT3 #(
		.INIT('h80)
	) name3916 (
		_w3519_,
		_w3946_,
		_w3949_,
		_w3950_
	);
	LUT2 #(
		.INIT('h8)
	) name3917 (
		_w3945_,
		_w3950_,
		_w3951_
	);
	LUT4 #(
		.INIT('h0777)
	) name3918 (
		_w52_,
		_w72_,
		_w50_,
		_w43_,
		_w3952_
	);
	LUT4 #(
		.INIT('h8000)
	) name3919 (
		_w940_,
		_w1961_,
		_w2257_,
		_w3952_,
		_w3953_
	);
	LUT3 #(
		.INIT('h37)
	) name3920 (
		_w67_,
		_w78_,
		_w50_,
		_w3954_
	);
	LUT4 #(
		.INIT('h4000)
	) name3921 (
		_w301_,
		_w2210_,
		_w2803_,
		_w3954_,
		_w3955_
	);
	LUT3 #(
		.INIT('h80)
	) name3922 (
		_w2468_,
		_w3099_,
		_w3341_,
		_w3956_
	);
	LUT4 #(
		.INIT('h8000)
	) name3923 (
		_w2511_,
		_w3955_,
		_w3956_,
		_w3953_,
		_w3957_
	);
	LUT4 #(
		.INIT('h8000)
	) name3924 (
		_w2236_,
		_w2240_,
		_w2486_,
		_w2487_,
		_w3958_
	);
	LUT4 #(
		.INIT('h8000)
	) name3925 (
		_w3945_,
		_w3950_,
		_w3957_,
		_w3958_,
		_w3959_
	);
	LUT2 #(
		.INIT('h8)
	) name3926 (
		_w1426_,
		_w3959_,
		_w3960_
	);
	LUT3 #(
		.INIT('h95)
	) name3927 (
		\a[2] ,
		_w1426_,
		_w3959_,
		_w3961_
	);
	LUT3 #(
		.INIT('h70)
	) name3928 (
		_w1973_,
		_w1997_,
		_w2407_,
		_w3962_
	);
	LUT3 #(
		.INIT('h70)
	) name3929 (
		_w1501_,
		_w1949_,
		_w2527_,
		_w3963_
	);
	LUT3 #(
		.INIT('h2a)
	) name3930 (
		_w376_,
		_w2023_,
		_w2055_,
		_w3964_
	);
	LUT3 #(
		.INIT('h01)
	) name3931 (
		_w3963_,
		_w3964_,
		_w3962_,
		_w3965_
	);
	LUT4 #(
		.INIT('h7d00)
	) name3932 (
		_w377_,
		_w2303_,
		_w2305_,
		_w3965_,
		_w3966_
	);
	LUT4 #(
		.INIT('hd554)
	) name3933 (
		\a[2] ,
		_w3943_,
		_w3960_,
		_w3966_,
		_w3967_
	);
	LUT3 #(
		.INIT('h95)
	) name3934 (
		\a[2] ,
		_w3929_,
		_w3930_,
		_w3968_
	);
	LUT4 #(
		.INIT('h6999)
	) name3935 (
		\a[2] ,
		\a[5] ,
		_w3151_,
		_w3818_,
		_w3969_
	);
	LUT4 #(
		.INIT('h2b00)
	) name3936 (
		\a[2] ,
		_w3931_,
		_w3967_,
		_w3969_,
		_w3970_
	);
	LUT4 #(
		.INIT('h00d4)
	) name3937 (
		\a[2] ,
		_w3931_,
		_w3967_,
		_w3969_,
		_w3971_
	);
	LUT4 #(
		.INIT('h54ab)
	) name3938 (
		_w1930_,
		_w2307_,
		_w2308_,
		_w2310_,
		_w3972_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3939 (
		_w1817_,
		_w1799_,
		_w1840_,
		_w2527_,
		_w3973_
	);
	LUT3 #(
		.INIT('h2a)
	) name3940 (
		_w376_,
		_w1898_,
		_w1928_,
		_w3974_
	);
	LUT3 #(
		.INIT('h70)
	) name3941 (
		_w1863_,
		_w1875_,
		_w2407_,
		_w3975_
	);
	LUT3 #(
		.INIT('h01)
	) name3942 (
		_w3974_,
		_w3975_,
		_w3973_,
		_w3976_
	);
	LUT3 #(
		.INIT('h70)
	) name3943 (
		_w377_,
		_w3972_,
		_w3976_,
		_w3977_
	);
	LUT3 #(
		.INIT('h54)
	) name3944 (
		_w3970_,
		_w3971_,
		_w3977_,
		_w3978_
	);
	LUT2 #(
		.INIT('h2)
	) name3945 (
		_w3917_,
		_w3978_,
		_w3979_
	);
	LUT2 #(
		.INIT('h4)
	) name3946 (
		_w3917_,
		_w3978_,
		_w3980_
	);
	LUT2 #(
		.INIT('h9)
	) name3947 (
		_w3917_,
		_w3978_,
		_w3981_
	);
	LUT3 #(
		.INIT('h70)
	) name3948 (
		_w1692_,
		_w1723_,
		_w2617_,
		_w3982_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3949 (
		_w1751_,
		_w1742_,
		_w1771_,
		_w2549_,
		_w3983_
	);
	LUT3 #(
		.INIT('h70)
	) name3950 (
		_w1620_,
		_w1661_,
		_w2854_,
		_w3984_
	);
	LUT3 #(
		.INIT('h01)
	) name3951 (
		_w3983_,
		_w3984_,
		_w3982_,
		_w3985_
	);
	LUT4 #(
		.INIT('h95aa)
	) name3952 (
		\a[29] ,
		_w2550_,
		_w3599_,
		_w3985_,
		_w3986_
	);
	LUT2 #(
		.INIT('h9)
	) name3953 (
		_w3908_,
		_w3914_,
		_w3987_
	);
	LUT4 #(
		.INIT('h2b00)
	) name3954 (
		_w3917_,
		_w3978_,
		_w3986_,
		_w3987_,
		_w3988_
	);
	LUT4 #(
		.INIT('h222b)
	) name3955 (
		_w3906_,
		_w3907_,
		_w3915_,
		_w3988_,
		_w3989_
	);
	LUT3 #(
		.INIT('h69)
	) name3956 (
		\a[29] ,
		_w3837_,
		_w3842_,
		_w3990_
	);
	LUT2 #(
		.INIT('h4)
	) name3957 (
		_w3989_,
		_w3990_,
		_w3991_
	);
	LUT2 #(
		.INIT('h2)
	) name3958 (
		_w3989_,
		_w3990_,
		_w3992_
	);
	LUT3 #(
		.INIT('h70)
	) name3959 (
		_w1381_,
		_w1398_,
		_w2874_,
		_w3993_
	);
	LUT3 #(
		.INIT('h70)
	) name3960 (
		_w1325_,
		_w1367_,
		_w2975_,
		_w3994_
	);
	LUT3 #(
		.INIT('h70)
	) name3961 (
		_w1253_,
		_w1294_,
		_w2986_,
		_w3995_
	);
	LUT3 #(
		.INIT('h01)
	) name3962 (
		_w3994_,
		_w3995_,
		_w3993_,
		_w3996_
	);
	LUT4 #(
		.INIT('h95aa)
	) name3963 (
		\a[26] ,
		_w2875_,
		_w3182_,
		_w3996_,
		_w3997_
	);
	LUT3 #(
		.INIT('h54)
	) name3964 (
		_w3991_,
		_w3992_,
		_w3997_,
		_w3998_
	);
	LUT2 #(
		.INIT('h2)
	) name3965 (
		_w3901_,
		_w3998_,
		_w3999_
	);
	LUT2 #(
		.INIT('h4)
	) name3966 (
		_w3901_,
		_w3998_,
		_w4000_
	);
	LUT3 #(
		.INIT('h2a)
	) name3967 (
		_w3214_,
		_w1136_,
		_w1187_,
		_w4001_
	);
	LUT3 #(
		.INIT('h70)
	) name3968 (
		_w1009_,
		_w1050_,
		_w3262_,
		_w4002_
	);
	LUT3 #(
		.INIT('h70)
	) name3969 (
		_w1071_,
		_w1102_,
		_w3249_,
		_w4003_
	);
	LUT3 #(
		.INIT('h01)
	) name3970 (
		_w4002_,
		_w4003_,
		_w4001_,
		_w4004_
	);
	LUT4 #(
		.INIT('h95aa)
	) name3971 (
		\a[23] ,
		_w2936_,
		_w37_,
		_w4004_,
		_w4005_
	);
	LUT3 #(
		.INIT('h54)
	) name3972 (
		_w3999_,
		_w4000_,
		_w4005_,
		_w4006_
	);
	LUT3 #(
		.INIT('h54)
	) name3973 (
		_w3897_,
		_w3898_,
		_w4006_,
		_w4007_
	);
	LUT2 #(
		.INIT('h9)
	) name3974 (
		_w3852_,
		_w3853_,
		_w4008_
	);
	LUT2 #(
		.INIT('h6)
	) name3975 (
		_w3860_,
		_w4008_,
		_w4009_
	);
	LUT3 #(
		.INIT('h70)
	) name3976 (
		_w725_,
		_w764_,
		_w3645_,
		_w4010_
	);
	LUT3 #(
		.INIT('h70)
	) name3977 (
		_w801_,
		_w851_,
		_w3311_,
		_w4011_
	);
	LUT3 #(
		.INIT('h70)
	) name3978 (
		_w666_,
		_w694_,
		_w3654_,
		_w4012_
	);
	LUT3 #(
		.INIT('h01)
	) name3979 (
		_w4011_,
		_w4012_,
		_w4010_,
		_w4013_
	);
	LUT4 #(
		.INIT('h6f00)
	) name3980 (
		_w2347_,
		_w2349_,
		_w3312_,
		_w4013_,
		_w4014_
	);
	LUT4 #(
		.INIT('hd4e8)
	) name3981 (
		\a[20] ,
		_w4007_,
		_w4009_,
		_w4014_,
		_w4015_
	);
	LUT3 #(
		.INIT('h09)
	) name3982 (
		_w3868_,
		_w3890_,
		_w4015_,
		_w4016_
	);
	LUT3 #(
		.INIT('h60)
	) name3983 (
		_w3868_,
		_w3890_,
		_w4015_,
		_w4017_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3984 (
		_w486_,
		_w487_,
		_w509_,
		_w3877_,
		_w4018_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3985 (
		_w121_,
		_w418_,
		_w422_,
		_w3886_,
		_w4019_
	);
	LUT3 #(
		.INIT('h70)
	) name3986 (
		_w544_,
		_w558_,
		_w3709_,
		_w4020_
	);
	LUT3 #(
		.INIT('h01)
	) name3987 (
		_w4018_,
		_w4019_,
		_w4020_,
		_w4021_
	);
	LUT4 #(
		.INIT('h6f00)
	) name3988 (
		_w2355_,
		_w2357_,
		_w3710_,
		_w4021_,
		_w4022_
	);
	LUT4 #(
		.INIT('h3132)
	) name3989 (
		\a[17] ,
		_w4016_,
		_w4017_,
		_w4022_,
		_w4023_
	);
	LUT2 #(
		.INIT('h9)
	) name3990 (
		_w3781_,
		_w3869_,
		_w4024_
	);
	LUT3 #(
		.INIT('h8e)
	) name3991 (
		_w3889_,
		_w4023_,
		_w4024_,
		_w4025_
	);
	LUT2 #(
		.INIT('h9)
	) name3992 (
		_w3870_,
		_w3872_,
		_w4026_
	);
	LUT2 #(
		.INIT('h6)
	) name3993 (
		_w3880_,
		_w4026_,
		_w4027_
	);
	LUT3 #(
		.INIT('h21)
	) name3994 (
		_w3880_,
		_w4025_,
		_w4026_,
		_w4028_
	);
	LUT3 #(
		.INIT('h48)
	) name3995 (
		_w3880_,
		_w4025_,
		_w4026_,
		_w4029_
	);
	LUT3 #(
		.INIT('h96)
	) name3996 (
		_w3880_,
		_w4025_,
		_w4026_,
		_w4030_
	);
	LUT3 #(
		.INIT('h96)
	) name3997 (
		_w3889_,
		_w4023_,
		_w4024_,
		_w4031_
	);
	LUT2 #(
		.INIT('h9)
	) name3998 (
		\a[11] ,
		\a[12] ,
		_w4032_
	);
	LUT4 #(
		.INIT('h0180)
	) name3999 (
		\a[11] ,
		\a[12] ,
		\a[13] ,
		\a[14] ,
		_w4033_
	);
	LUT4 #(
		.INIT('h0660)
	) name4000 (
		\a[11] ,
		\a[12] ,
		\a[13] ,
		\a[14] ,
		_w4034_
	);
	LUT4 #(
		.INIT('h5150)
	) name4001 (
		_w374_,
		_w2361_,
		_w4033_,
		_w4034_,
		_w4035_
	);
	LUT2 #(
		.INIT('h9)
	) name4002 (
		_w3899_,
		_w4006_,
		_w4036_
	);
	LUT3 #(
		.INIT('h70)
	) name4003 (
		_w725_,
		_w764_,
		_w3654_,
		_w4037_
	);
	LUT3 #(
		.INIT('h70)
	) name4004 (
		_w801_,
		_w851_,
		_w3645_,
		_w4038_
	);
	LUT3 #(
		.INIT('h70)
	) name4005 (
		_w871_,
		_w927_,
		_w3311_,
		_w4039_
	);
	LUT3 #(
		.INIT('h01)
	) name4006 (
		_w4038_,
		_w4039_,
		_w4037_,
		_w4040_
	);
	LUT4 #(
		.INIT('h95aa)
	) name4007 (
		\a[20] ,
		_w2724_,
		_w3312_,
		_w4040_,
		_w4041_
	);
	LUT2 #(
		.INIT('h9)
	) name4008 (
		_w3901_,
		_w3998_,
		_w4042_
	);
	LUT4 #(
		.INIT('h6669)
	) name4009 (
		_w3906_,
		_w3907_,
		_w3915_,
		_w3988_,
		_w4043_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4010 (
		_w1454_,
		_w1426_,
		_w1478_,
		_w2874_,
		_w4044_
	);
	LUT3 #(
		.INIT('h70)
	) name4011 (
		_w1325_,
		_w1367_,
		_w2986_,
		_w4045_
	);
	LUT3 #(
		.INIT('h70)
	) name4012 (
		_w1381_,
		_w1398_,
		_w2975_,
		_w4046_
	);
	LUT3 #(
		.INIT('h01)
	) name4013 (
		_w4045_,
		_w4046_,
		_w4044_,
		_w4047_
	);
	LUT4 #(
		.INIT('h6f00)
	) name4014 (
		_w2327_,
		_w2329_,
		_w2875_,
		_w4047_,
		_w4048_
	);
	LUT3 #(
		.INIT('h84)
	) name4015 (
		\a[26] ,
		_w4043_,
		_w4048_,
		_w4049_
	);
	LUT3 #(
		.INIT('h12)
	) name4016 (
		\a[26] ,
		_w4043_,
		_w4048_,
		_w4050_
	);
	LUT3 #(
		.INIT('h69)
	) name4017 (
		\a[26] ,
		_w4043_,
		_w4048_,
		_w4051_
	);
	LUT3 #(
		.INIT('h70)
	) name4018 (
		_w1692_,
		_w1723_,
		_w2549_,
		_w4052_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4019 (
		_w1584_,
		_w1569_,
		_w1606_,
		_w2854_,
		_w4053_
	);
	LUT3 #(
		.INIT('h70)
	) name4020 (
		_w1620_,
		_w1661_,
		_w2617_,
		_w4054_
	);
	LUT3 #(
		.INIT('h01)
	) name4021 (
		_w4053_,
		_w4054_,
		_w4052_,
		_w4055_
	);
	LUT4 #(
		.INIT('h6f00)
	) name4022 (
		_w2319_,
		_w2321_,
		_w2550_,
		_w4055_,
		_w4056_
	);
	LUT2 #(
		.INIT('h6)
	) name4023 (
		\a[29] ,
		_w4056_,
		_w4057_
	);
	LUT4 #(
		.INIT('h54ab)
	) name4024 (
		_w3979_,
		_w3980_,
		_w3986_,
		_w3987_,
		_w4058_
	);
	LUT2 #(
		.INIT('h4)
	) name4025 (
		_w4057_,
		_w4058_,
		_w4059_
	);
	LUT2 #(
		.INIT('h2)
	) name4026 (
		_w4057_,
		_w4058_,
		_w4060_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4027 (
		_w1454_,
		_w1426_,
		_w1478_,
		_w2975_,
		_w4061_
	);
	LUT3 #(
		.INIT('h70)
	) name4028 (
		_w1381_,
		_w1398_,
		_w2986_,
		_w4062_
	);
	LUT3 #(
		.INIT('h70)
	) name4029 (
		_w1501_,
		_w1545_,
		_w2874_,
		_w4063_
	);
	LUT3 #(
		.INIT('h01)
	) name4030 (
		_w4062_,
		_w4063_,
		_w4061_,
		_w4064_
	);
	LUT4 #(
		.INIT('h95aa)
	) name4031 (
		\a[26] ,
		_w2875_,
		_w3362_,
		_w4064_,
		_w4065_
	);
	LUT3 #(
		.INIT('h54)
	) name4032 (
		_w4059_,
		_w4060_,
		_w4065_,
		_w4066_
	);
	LUT3 #(
		.INIT('h54)
	) name4033 (
		_w4049_,
		_w4050_,
		_w4066_,
		_w4067_
	);
	LUT2 #(
		.INIT('h9)
	) name4034 (
		_w3989_,
		_w3990_,
		_w4068_
	);
	LUT2 #(
		.INIT('h9)
	) name4035 (
		_w3997_,
		_w4068_,
		_w4069_
	);
	LUT3 #(
		.INIT('h70)
	) name4036 (
		_w1136_,
		_w1187_,
		_w3249_,
		_w4070_
	);
	LUT3 #(
		.INIT('h70)
	) name4037 (
		_w1071_,
		_w1102_,
		_w3262_,
		_w4071_
	);
	LUT3 #(
		.INIT('h2a)
	) name4038 (
		_w3214_,
		_w1202_,
		_w1233_,
		_w4072_
	);
	LUT3 #(
		.INIT('h01)
	) name4039 (
		_w4071_,
		_w4072_,
		_w4070_,
		_w4073_
	);
	LUT4 #(
		.INIT('h6f00)
	) name4040 (
		_w2335_,
		_w2337_,
		_w37_,
		_w4073_,
		_w4074_
	);
	LUT4 #(
		.INIT('h4d8e)
	) name4041 (
		\a[23] ,
		_w4067_,
		_w4069_,
		_w4074_,
		_w4075_
	);
	LUT3 #(
		.INIT('h09)
	) name4042 (
		_w4005_,
		_w4042_,
		_w4075_,
		_w4076_
	);
	LUT3 #(
		.INIT('h60)
	) name4043 (
		_w4005_,
		_w4042_,
		_w4075_,
		_w4077_
	);
	LUT3 #(
		.INIT('h70)
	) name4044 (
		_w763_,
		_w983_,
		_w3311_,
		_w4078_
	);
	LUT3 #(
		.INIT('h70)
	) name4045 (
		_w871_,
		_w927_,
		_w3645_,
		_w4079_
	);
	LUT3 #(
		.INIT('h70)
	) name4046 (
		_w801_,
		_w851_,
		_w3654_,
		_w4080_
	);
	LUT3 #(
		.INIT('h01)
	) name4047 (
		_w4079_,
		_w4080_,
		_w4078_,
		_w4081_
	);
	LUT4 #(
		.INIT('h6f00)
	) name4048 (
		_w2343_,
		_w2345_,
		_w3312_,
		_w4081_,
		_w4082_
	);
	LUT4 #(
		.INIT('h3132)
	) name4049 (
		\a[20] ,
		_w4076_,
		_w4077_,
		_w4082_,
		_w4083_
	);
	LUT3 #(
		.INIT('hd4)
	) name4050 (
		_w4036_,
		_w4041_,
		_w4083_,
		_w4084_
	);
	LUT4 #(
		.INIT('h9669)
	) name4051 (
		\a[20] ,
		_w4007_,
		_w4009_,
		_w4014_,
		_w4085_
	);
	LUT2 #(
		.INIT('h4)
	) name4052 (
		_w4084_,
		_w4085_,
		_w4086_
	);
	LUT2 #(
		.INIT('h2)
	) name4053 (
		_w4084_,
		_w4085_,
		_w4087_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4054 (
		_w486_,
		_w487_,
		_w509_,
		_w3886_,
		_w4088_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4055 (
		_w587_,
		_w608_,
		_w624_,
		_w3709_,
		_w4089_
	);
	LUT3 #(
		.INIT('h70)
	) name4056 (
		_w544_,
		_w558_,
		_w3877_,
		_w4090_
	);
	LUT3 #(
		.INIT('h01)
	) name4057 (
		_w4088_,
		_w4089_,
		_w4090_,
		_w4091_
	);
	LUT4 #(
		.INIT('h95aa)
	) name4058 (
		\a[17] ,
		_w2526_,
		_w3710_,
		_w4091_,
		_w4092_
	);
	LUT3 #(
		.INIT('h54)
	) name4059 (
		_w4086_,
		_w4087_,
		_w4092_,
		_w4093_
	);
	LUT3 #(
		.INIT('h96)
	) name4060 (
		_w3868_,
		_w3890_,
		_w4015_,
		_w4094_
	);
	LUT3 #(
		.INIT('h69)
	) name4061 (
		\a[17] ,
		_w4022_,
		_w4094_,
		_w4095_
	);
	LUT4 #(
		.INIT('h90f9)
	) name4062 (
		\a[14] ,
		_w4035_,
		_w4093_,
		_w4095_,
		_w4096_
	);
	LUT2 #(
		.INIT('h2)
	) name4063 (
		_w4031_,
		_w4096_,
		_w4097_
	);
	LUT2 #(
		.INIT('h4)
	) name4064 (
		_w4031_,
		_w4096_,
		_w4098_
	);
	LUT2 #(
		.INIT('h9)
	) name4065 (
		_w4031_,
		_w4096_,
		_w4099_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4066 (
		_w587_,
		_w608_,
		_w624_,
		_w3877_,
		_w4100_
	);
	LUT3 #(
		.INIT('h70)
	) name4067 (
		_w666_,
		_w694_,
		_w3709_,
		_w4101_
	);
	LUT3 #(
		.INIT('h70)
	) name4068 (
		_w544_,
		_w558_,
		_w3886_,
		_w4102_
	);
	LUT3 #(
		.INIT('h01)
	) name4069 (
		_w4101_,
		_w4102_,
		_w4100_,
		_w4103_
	);
	LUT4 #(
		.INIT('h6f00)
	) name4070 (
		_w2351_,
		_w2353_,
		_w3710_,
		_w4103_,
		_w4104_
	);
	LUT3 #(
		.INIT('h96)
	) name4071 (
		_w4036_,
		_w4041_,
		_w4083_,
		_w4105_
	);
	LUT3 #(
		.INIT('h90)
	) name4072 (
		\a[17] ,
		_w4104_,
		_w4105_,
		_w4106_
	);
	LUT3 #(
		.INIT('h06)
	) name4073 (
		\a[17] ,
		_w4104_,
		_w4105_,
		_w4107_
	);
	LUT3 #(
		.INIT('h69)
	) name4074 (
		\a[17] ,
		_w4104_,
		_w4105_,
		_w4108_
	);
	LUT3 #(
		.INIT('h96)
	) name4075 (
		_w4005_,
		_w4042_,
		_w4075_,
		_w4109_
	);
	LUT3 #(
		.INIT('h69)
	) name4076 (
		\a[20] ,
		_w4082_,
		_w4109_,
		_w4110_
	);
	LUT3 #(
		.INIT('h70)
	) name4077 (
		_w1202_,
		_w1233_,
		_w3249_,
		_w4111_
	);
	LUT3 #(
		.INIT('h2a)
	) name4078 (
		_w3214_,
		_w1253_,
		_w1294_,
		_w4112_
	);
	LUT3 #(
		.INIT('h70)
	) name4079 (
		_w1136_,
		_w1187_,
		_w3262_,
		_w4113_
	);
	LUT3 #(
		.INIT('h01)
	) name4080 (
		_w4112_,
		_w4113_,
		_w4111_,
		_w4114_
	);
	LUT4 #(
		.INIT('h95aa)
	) name4081 (
		\a[23] ,
		_w3067_,
		_w37_,
		_w4114_,
		_w4115_
	);
	LUT2 #(
		.INIT('h9)
	) name4082 (
		_w4051_,
		_w4066_,
		_w4116_
	);
	LUT2 #(
		.INIT('h9)
	) name4083 (
		_w4057_,
		_w4058_,
		_w4117_
	);
	LUT2 #(
		.INIT('h9)
	) name4084 (
		_w3981_,
		_w3986_,
		_w4118_
	);
	LUT3 #(
		.INIT('h70)
	) name4085 (
		_w1898_,
		_w1928_,
		_w2407_,
		_w4119_
	);
	LUT3 #(
		.INIT('h2a)
	) name4086 (
		_w376_,
		_w1501_,
		_w1949_,
		_w4120_
	);
	LUT3 #(
		.INIT('h70)
	) name4087 (
		_w1863_,
		_w1875_,
		_w2527_,
		_w4121_
	);
	LUT3 #(
		.INIT('h01)
	) name4088 (
		_w4120_,
		_w4121_,
		_w4119_,
		_w4122_
	);
	LUT4 #(
		.INIT('h7d00)
	) name4089 (
		_w377_,
		_w2307_,
		_w2309_,
		_w4122_,
		_w4123_
	);
	LUT3 #(
		.INIT('h09)
	) name4090 (
		_w3967_,
		_w3968_,
		_w4123_,
		_w4124_
	);
	LUT4 #(
		.INIT('h9336)
	) name4091 (
		\a[2] ,
		_w3943_,
		_w3960_,
		_w3966_,
		_w4125_
	);
	LUT4 #(
		.INIT('h54ab)
	) name4092 (
		_w1999_,
		_w2303_,
		_w2304_,
		_w2306_,
		_w4126_
	);
	LUT3 #(
		.INIT('h2a)
	) name4093 (
		_w376_,
		_w1973_,
		_w1997_,
		_w4127_
	);
	LUT3 #(
		.INIT('h70)
	) name4094 (
		_w1898_,
		_w1928_,
		_w2527_,
		_w4128_
	);
	LUT3 #(
		.INIT('h70)
	) name4095 (
		_w1501_,
		_w1949_,
		_w2407_,
		_w4129_
	);
	LUT3 #(
		.INIT('h01)
	) name4096 (
		_w4128_,
		_w4129_,
		_w4127_,
		_w4130_
	);
	LUT3 #(
		.INIT('h70)
	) name4097 (
		_w377_,
		_w4126_,
		_w4130_,
		_w4131_
	);
	LUT2 #(
		.INIT('h2)
	) name4098 (
		_w4125_,
		_w4131_,
		_w4132_
	);
	LUT4 #(
		.INIT('h135f)
	) name4099 (
		_w106_,
		_w55_,
		_w90_,
		_w176_,
		_w4133_
	);
	LUT2 #(
		.INIT('h8)
	) name4100 (
		_w472_,
		_w4133_,
		_w4134_
	);
	LUT4 #(
		.INIT('h0400)
	) name4101 (
		_w61_,
		_w370_,
		_w462_,
		_w2454_,
		_w4135_
	);
	LUT2 #(
		.INIT('h8)
	) name4102 (
		_w4134_,
		_w4135_,
		_w4136_
	);
	LUT3 #(
		.INIT('h40)
	) name4103 (
		_w167_,
		_w877_,
		_w3521_,
		_w4137_
	);
	LUT4 #(
		.INIT('h8000)
	) name4104 (
		_w1438_,
		_w1687_,
		_w1791_,
		_w2143_,
		_w4138_
	);
	LUT3 #(
		.INIT('h80)
	) name4105 (
		_w163_,
		_w844_,
		_w1092_,
		_w4139_
	);
	LUT3 #(
		.INIT('h80)
	) name4106 (
		_w4137_,
		_w4138_,
		_w4139_,
		_w4140_
	);
	LUT3 #(
		.INIT('h80)
	) name4107 (
		_w3143_,
		_w4136_,
		_w4140_,
		_w4141_
	);
	LUT4 #(
		.INIT('h8000)
	) name4108 (
		_w1222_,
		_w1275_,
		_w1362_,
		_w1470_,
		_w4142_
	);
	LUT3 #(
		.INIT('h37)
	) name4109 (
		_w122_,
		_w67_,
		_w166_,
		_w4143_
	);
	LUT4 #(
		.INIT('h135f)
	) name4110 (
		_w122_,
		_w90_,
		_w56_,
		_w430_,
		_w4144_
	);
	LUT4 #(
		.INIT('h2000)
	) name4111 (
		_w245_,
		_w437_,
		_w4143_,
		_w4144_,
		_w4145_
	);
	LUT3 #(
		.INIT('h80)
	) name4112 (
		_w2176_,
		_w3336_,
		_w3449_,
		_w4146_
	);
	LUT4 #(
		.INIT('h8000)
	) name4113 (
		_w3102_,
		_w4146_,
		_w4142_,
		_w4145_,
		_w4147_
	);
	LUT2 #(
		.INIT('h8)
	) name4114 (
		_w1757_,
		_w4147_,
		_w4148_
	);
	LUT4 #(
		.INIT('h8000)
	) name4115 (
		_w1757_,
		_w3157_,
		_w3161_,
		_w4147_,
		_w4149_
	);
	LUT2 #(
		.INIT('h8)
	) name4116 (
		_w4141_,
		_w4149_,
		_w4150_
	);
	LUT4 #(
		.INIT('h54ab)
	) name4117 (
		_w2101_,
		_w2299_,
		_w2300_,
		_w2302_,
		_w4151_
	);
	LUT3 #(
		.INIT('h70)
	) name4118 (
		_w1973_,
		_w1997_,
		_w2527_,
		_w4152_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name4119 (
		_w376_,
		_w1874_,
		_w2076_,
		_w2099_,
		_w4153_
	);
	LUT3 #(
		.INIT('h70)
	) name4120 (
		_w2023_,
		_w2055_,
		_w2407_,
		_w4154_
	);
	LUT3 #(
		.INIT('h01)
	) name4121 (
		_w4153_,
		_w4154_,
		_w4152_,
		_w4155_
	);
	LUT3 #(
		.INIT('h70)
	) name4122 (
		_w377_,
		_w4151_,
		_w4155_,
		_w4156_
	);
	LUT4 #(
		.INIT('h2033)
	) name4123 (
		_w377_,
		_w4150_,
		_w4151_,
		_w4155_,
		_w4157_
	);
	LUT4 #(
		.INIT('h153f)
	) name4124 (
		_w56_,
		_w39_,
		_w46_,
		_w201_,
		_w4158_
	);
	LUT3 #(
		.INIT('h80)
	) name4125 (
		_w997_,
		_w1332_,
		_w4158_,
		_w4159_
	);
	LUT3 #(
		.INIT('h80)
	) name4126 (
		_w1682_,
		_w1976_,
		_w2440_,
		_w4160_
	);
	LUT4 #(
		.INIT('h8000)
	) name4127 (
		_w1003_,
		_w1216_,
		_w1704_,
		_w1687_,
		_w4161_
	);
	LUT3 #(
		.INIT('h80)
	) name4128 (
		_w4159_,
		_w4160_,
		_w4161_,
		_w4162_
	);
	LUT4 #(
		.INIT('h135f)
	) name4129 (
		_w52_,
		_w67_,
		_w176_,
		_w430_,
		_w4163_
	);
	LUT4 #(
		.INIT('h8000)
	) name4130 (
		_w538_,
		_w663_,
		_w767_,
		_w4163_,
		_w4164_
	);
	LUT4 #(
		.INIT('h135f)
	) name4131 (
		_w52_,
		_w44_,
		_w184_,
		_w378_,
		_w4165_
	);
	LUT2 #(
		.INIT('h8)
	) name4132 (
		_w1359_,
		_w4165_,
		_w4166_
	);
	LUT4 #(
		.INIT('h8000)
	) name4133 (
		_w150_,
		_w1359_,
		_w2510_,
		_w4165_,
		_w4167_
	);
	LUT4 #(
		.INIT('h8000)
	) name4134 (
		_w3458_,
		_w3461_,
		_w4164_,
		_w4167_,
		_w4168_
	);
	LUT4 #(
		.INIT('h0800)
	) name4135 (
		_w292_,
		_w274_,
		_w424_,
		_w842_,
		_w4169_
	);
	LUT4 #(
		.INIT('h153f)
	) name4136 (
		_w59_,
		_w39_,
		_w44_,
		_w184_,
		_w4170_
	);
	LUT4 #(
		.INIT('h1000)
	) name4137 (
		_w286_,
		_w390_,
		_w3439_,
		_w4170_,
		_w4171_
	);
	LUT4 #(
		.INIT('h0777)
	) name4138 (
		_w106_,
		_w59_,
		_w41_,
		_w158_,
		_w4172_
	);
	LUT4 #(
		.INIT('h8000)
	) name4139 (
		_w935_,
		_w2418_,
		_w3507_,
		_w4172_,
		_w4173_
	);
	LUT4 #(
		.INIT('h8000)
	) name4140 (
		_w3038_,
		_w4173_,
		_w4169_,
		_w4171_,
		_w4174_
	);
	LUT4 #(
		.INIT('h8000)
	) name4141 (
		_w982_,
		_w4174_,
		_w4162_,
		_w4168_,
		_w4175_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4142 (
		_w1874_,
		_w2076_,
		_w2099_,
		_w2407_,
		_w4176_
	);
	LUT3 #(
		.INIT('h2a)
	) name4143 (
		_w376_,
		_w2124_,
		_w2133_,
		_w4177_
	);
	LUT3 #(
		.INIT('h70)
	) name4144 (
		_w2023_,
		_w2055_,
		_w2527_,
		_w4178_
	);
	LUT3 #(
		.INIT('h01)
	) name4145 (
		_w4176_,
		_w4177_,
		_w4178_,
		_w4179_
	);
	LUT4 #(
		.INIT('h7d00)
	) name4146 (
		_w377_,
		_w2299_,
		_w2301_,
		_w4179_,
		_w4180_
	);
	LUT2 #(
		.INIT('h1)
	) name4147 (
		_w4175_,
		_w4180_,
		_w4181_
	);
	LUT3 #(
		.INIT('h1f)
	) name4148 (
		_w38_,
		_w46_,
		_w166_,
		_w4182_
	);
	LUT4 #(
		.INIT('h1000)
	) name4149 (
		_w339_,
		_w441_,
		_w1945_,
		_w4182_,
		_w4183_
	);
	LUT4 #(
		.INIT('h153f)
	) name4150 (
		_w67_,
		_w43_,
		_w65_,
		_w184_,
		_w4184_
	);
	LUT3 #(
		.INIT('h57)
	) name4151 (
		_w52_,
		_w158_,
		_w378_,
		_w4185_
	);
	LUT2 #(
		.INIT('h8)
	) name4152 (
		_w4184_,
		_w4185_,
		_w4186_
	);
	LUT3 #(
		.INIT('h80)
	) name4153 (
		_w744_,
		_w1456_,
		_w1562_,
		_w4187_
	);
	LUT3 #(
		.INIT('h80)
	) name4154 (
		_w4183_,
		_w4186_,
		_w4187_,
		_w4188_
	);
	LUT4 #(
		.INIT('h0777)
	) name4155 (
		_w85_,
		_w78_,
		_w56_,
		_w39_,
		_w4189_
	);
	LUT4 #(
		.INIT('h8000)
	) name4156 (
		_w966_,
		_w935_,
		_w1975_,
		_w4189_,
		_w4190_
	);
	LUT4 #(
		.INIT('h153f)
	) name4157 (
		_w55_,
		_w50_,
		_w259_,
		_w378_,
		_w4191_
	);
	LUT4 #(
		.INIT('h1000)
	) name4158 (
		_w294_,
		_w439_,
		_w1211_,
		_w4191_,
		_w4192_
	);
	LUT2 #(
		.INIT('h8)
	) name4159 (
		_w4190_,
		_w4192_,
		_w4193_
	);
	LUT4 #(
		.INIT('h8000)
	) name4160 (
		_w588_,
		_w591_,
		_w2009_,
		_w2013_,
		_w4194_
	);
	LUT3 #(
		.INIT('h80)
	) name4161 (
		_w4193_,
		_w4188_,
		_w4194_,
		_w4195_
	);
	LUT2 #(
		.INIT('h2)
	) name4162 (
		_w81_,
		_w402_,
		_w4196_
	);
	LUT4 #(
		.INIT('h135f)
	) name4163 (
		_w47_,
		_w41_,
		_w43_,
		_w158_,
		_w4197_
	);
	LUT4 #(
		.INIT('h4000)
	) name4164 (
		_w285_,
		_w908_,
		_w1617_,
		_w4197_,
		_w4198_
	);
	LUT2 #(
		.INIT('h8)
	) name4165 (
		_w4196_,
		_w4198_,
		_w4199_
	);
	LUT4 #(
		.INIT('h153f)
	) name4166 (
		_w38_,
		_w65_,
		_w176_,
		_w378_,
		_w4200_
	);
	LUT4 #(
		.INIT('h8000)
	) name4167 (
		_w1480_,
		_w1629_,
		_w1784_,
		_w4200_,
		_w4201_
	);
	LUT4 #(
		.INIT('h3337)
	) name4168 (
		_w52_,
		_w72_,
		_w93_,
		_w44_,
		_w4202_
	);
	LUT2 #(
		.INIT('h8)
	) name4169 (
		_w2149_,
		_w4202_,
		_w4203_
	);
	LUT4 #(
		.INIT('h135f)
	) name4170 (
		_w56_,
		_w65_,
		_w176_,
		_w419_,
		_w4204_
	);
	LUT3 #(
		.INIT('h40)
	) name4171 (
		_w226_,
		_w538_,
		_w4204_,
		_w4205_
	);
	LUT4 #(
		.INIT('h8000)
	) name4172 (
		_w3509_,
		_w4203_,
		_w4205_,
		_w4201_,
		_w4206_
	);
	LUT4 #(
		.INIT('h8000)
	) name4173 (
		_w3537_,
		_w3548_,
		_w4199_,
		_w4206_,
		_w4207_
	);
	LUT2 #(
		.INIT('h8)
	) name4174 (
		_w4195_,
		_w4207_,
		_w4208_
	);
	LUT4 #(
		.INIT('h54ab)
	) name4175 (
		_w2158_,
		_w2295_,
		_w2296_,
		_w2298_,
		_w4209_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4176 (
		_w1874_,
		_w2076_,
		_w2099_,
		_w2527_,
		_w4210_
	);
	LUT3 #(
		.INIT('h2a)
	) name4177 (
		_w376_,
		_w2155_,
		_w2156_,
		_w4211_
	);
	LUT3 #(
		.INIT('h70)
	) name4178 (
		_w2124_,
		_w2133_,
		_w2407_,
		_w4212_
	);
	LUT3 #(
		.INIT('h01)
	) name4179 (
		_w4210_,
		_w4211_,
		_w4212_,
		_w4213_
	);
	LUT4 #(
		.INIT('h2033)
	) name4180 (
		_w377_,
		_w4208_,
		_w4209_,
		_w4213_,
		_w4214_
	);
	LUT4 #(
		.INIT('h153f)
	) name4181 (
		_w38_,
		_w67_,
		_w39_,
		_w184_,
		_w4215_
	);
	LUT4 #(
		.INIT('h135f)
	) name4182 (
		_w55_,
		_w44_,
		_w184_,
		_w259_,
		_w4216_
	);
	LUT4 #(
		.INIT('h8000)
	) name4183 (
		_w446_,
		_w1576_,
		_w4215_,
		_w4216_,
		_w4217_
	);
	LUT4 #(
		.INIT('h153f)
	) name4184 (
		_w59_,
		_w65_,
		_w419_,
		_w378_,
		_w4218_
	);
	LUT3 #(
		.INIT('h1f)
	) name4185 (
		_w110_,
		_w44_,
		_w430_,
		_w4219_
	);
	LUT3 #(
		.INIT('h80)
	) name4186 (
		_w113_,
		_w4218_,
		_w4219_,
		_w4220_
	);
	LUT3 #(
		.INIT('h80)
	) name4187 (
		_w2926_,
		_w4217_,
		_w4220_,
		_w4221_
	);
	LUT4 #(
		.INIT('h0777)
	) name4188 (
		_w78_,
		_w41_,
		_w43_,
		_w46_,
		_w4222_
	);
	LUT4 #(
		.INIT('h153f)
	) name4189 (
		_w52_,
		_w56_,
		_w158_,
		_w378_,
		_w4223_
	);
	LUT4 #(
		.INIT('h4000)
	) name4190 (
		_w369_,
		_w1165_,
		_w4222_,
		_w4223_,
		_w4224_
	);
	LUT4 #(
		.INIT('h153f)
	) name4191 (
		_w38_,
		_w90_,
		_w39_,
		_w419_,
		_w4225_
	);
	LUT4 #(
		.INIT('h8000)
	) name4192 (
		_w265_,
		_w2671_,
		_w2672_,
		_w4225_,
		_w4226_
	);
	LUT2 #(
		.INIT('h8)
	) name4193 (
		_w4224_,
		_w4226_,
		_w4227_
	);
	LUT4 #(
		.INIT('h0777)
	) name4194 (
		_w106_,
		_w52_,
		_w90_,
		_w72_,
		_w4228_
	);
	LUT2 #(
		.INIT('h4)
	) name4195 (
		_w298_,
		_w4228_,
		_w4229_
	);
	LUT4 #(
		.INIT('h153f)
	) name4196 (
		_w90_,
		_w72_,
		_w44_,
		_w176_,
		_w4230_
	);
	LUT4 #(
		.INIT('h2000)
	) name4197 (
		_w115_,
		_w298_,
		_w4230_,
		_w4228_,
		_w4231_
	);
	LUT4 #(
		.INIT('h8000)
	) name4198 (
		_w1156_,
		_w1318_,
		_w2231_,
		_w3099_,
		_w4232_
	);
	LUT4 #(
		.INIT('h8000)
	) name4199 (
		_w96_,
		_w305_,
		_w584_,
		_w790_,
		_w4233_
	);
	LUT3 #(
		.INIT('h80)
	) name4200 (
		_w4231_,
		_w4232_,
		_w4233_,
		_w4234_
	);
	LUT3 #(
		.INIT('h80)
	) name4201 (
		_w4221_,
		_w4227_,
		_w4234_,
		_w4235_
	);
	LUT2 #(
		.INIT('h8)
	) name4202 (
		_w1973_,
		_w4235_,
		_w4236_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name4203 (
		_w376_,
		_w2193_,
		_w2183_,
		_w2213_,
		_w4237_
	);
	LUT3 #(
		.INIT('h70)
	) name4204 (
		_w2155_,
		_w2156_,
		_w2407_,
		_w4238_
	);
	LUT3 #(
		.INIT('h70)
	) name4205 (
		_w2124_,
		_w2133_,
		_w2527_,
		_w4239_
	);
	LUT3 #(
		.INIT('h01)
	) name4206 (
		_w4237_,
		_w4238_,
		_w4239_,
		_w4240_
	);
	LUT4 #(
		.INIT('h7d00)
	) name4207 (
		_w377_,
		_w2295_,
		_w2297_,
		_w4240_,
		_w4241_
	);
	LUT2 #(
		.INIT('h1)
	) name4208 (
		_w4236_,
		_w4241_,
		_w4242_
	);
	LUT4 #(
		.INIT('h135f)
	) name4209 (
		_w85_,
		_w41_,
		_w158_,
		_w259_,
		_w4243_
	);
	LUT4 #(
		.INIT('h153f)
	) name4210 (
		_w85_,
		_w46_,
		_w259_,
		_w430_,
		_w4244_
	);
	LUT2 #(
		.INIT('h8)
	) name4211 (
		_w4243_,
		_w4244_,
		_w4245_
	);
	LUT3 #(
		.INIT('h80)
	) name4212 (
		_w960_,
		_w2281_,
		_w2705_,
		_w4246_
	);
	LUT2 #(
		.INIT('h8)
	) name4213 (
		_w4245_,
		_w4246_,
		_w4247_
	);
	LUT4 #(
		.INIT('h153f)
	) name4214 (
		_w55_,
		_w50_,
		_w166_,
		_w378_,
		_w4248_
	);
	LUT4 #(
		.INIT('h8000)
	) name4215 (
		_w597_,
		_w842_,
		_w1014_,
		_w4248_,
		_w4249_
	);
	LUT4 #(
		.INIT('h8000)
	) name4216 (
		_w678_,
		_w856_,
		_w857_,
		_w1113_,
		_w4250_
	);
	LUT3 #(
		.INIT('h1f)
	) name4217 (
		_w106_,
		_w39_,
		_w50_,
		_w4251_
	);
	LUT3 #(
		.INIT('h40)
	) name4218 (
		_w321_,
		_w790_,
		_w4251_,
		_w4252_
	);
	LUT4 #(
		.INIT('h8000)
	) name4219 (
		_w1221_,
		_w1664_,
		_w2494_,
		_w2640_,
		_w4253_
	);
	LUT4 #(
		.INIT('h8000)
	) name4220 (
		_w4252_,
		_w4253_,
		_w4249_,
		_w4250_,
		_w4254_
	);
	LUT3 #(
		.INIT('h80)
	) name4221 (
		_w1884_,
		_w4247_,
		_w4254_,
		_w4255_
	);
	LUT4 #(
		.INIT('h8000)
	) name4222 (
		_w2674_,
		_w2677_,
		_w3031_,
		_w3039_,
		_w4256_
	);
	LUT2 #(
		.INIT('h8)
	) name4223 (
		_w4255_,
		_w4256_,
		_w4257_
	);
	LUT4 #(
		.INIT('h0888)
	) name4224 (
		_w2228_,
		_w2262_,
		_w2273_,
		_w2293_,
		_w4258_
	);
	LUT3 #(
		.INIT('h82)
	) name4225 (
		_w377_,
		_w2214_,
		_w4258_,
		_w4259_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4226 (
		_w2193_,
		_w2183_,
		_w2213_,
		_w2527_,
		_w4260_
	);
	LUT3 #(
		.INIT('h70)
	) name4227 (
		_w2273_,
		_w2293_,
		_w2407_,
		_w4261_
	);
	LUT3 #(
		.INIT('h2a)
	) name4228 (
		_w376_,
		_w2228_,
		_w2262_,
		_w4262_
	);
	LUT3 #(
		.INIT('h01)
	) name4229 (
		_w4261_,
		_w4262_,
		_w4260_,
		_w4263_
	);
	LUT3 #(
		.INIT('h1f)
	) name4230 (
		_w110_,
		_w47_,
		_w43_,
		_w4264_
	);
	LUT3 #(
		.INIT('h1f)
	) name4231 (
		_w67_,
		_w46_,
		_w259_,
		_w4265_
	);
	LUT4 #(
		.INIT('h0777)
	) name4232 (
		_w90_,
		_w43_,
		_w46_,
		_w176_,
		_w4266_
	);
	LUT4 #(
		.INIT('h8000)
	) name4233 (
		_w2190_,
		_w4265_,
		_w4266_,
		_w4264_,
		_w4267_
	);
	LUT3 #(
		.INIT('h40)
	) name4234 (
		_w407_,
		_w1386_,
		_w2432_,
		_w4268_
	);
	LUT2 #(
		.INIT('h8)
	) name4235 (
		_w4267_,
		_w4268_,
		_w4269_
	);
	LUT4 #(
		.INIT('h153f)
	) name4236 (
		_w41_,
		_w46_,
		_w158_,
		_w419_,
		_w4270_
	);
	LUT4 #(
		.INIT('h4000)
	) name4237 (
		_w455_,
		_w960_,
		_w1924_,
		_w4270_,
		_w4271_
	);
	LUT3 #(
		.INIT('h10)
	) name4238 (
		_w186_,
		_w268_,
		_w1198_,
		_w4272_
	);
	LUT3 #(
		.INIT('h80)
	) name4239 (
		_w1637_,
		_w4272_,
		_w4271_,
		_w4273_
	);
	LUT3 #(
		.INIT('h80)
	) name4240 (
		_w2200_,
		_w4269_,
		_w4273_,
		_w4274_
	);
	LUT3 #(
		.INIT('h80)
	) name4241 (
		_w522_,
		_w512_,
		_w650_,
		_w4275_
	);
	LUT4 #(
		.INIT('h153f)
	) name4242 (
		_w122_,
		_w85_,
		_w43_,
		_w65_,
		_w4276_
	);
	LUT4 #(
		.INIT('h135f)
	) name4243 (
		_w106_,
		_w47_,
		_w50_,
		_w158_,
		_w4277_
	);
	LUT4 #(
		.INIT('h4000)
	) name4244 (
		_w57_,
		_w1631_,
		_w4276_,
		_w4277_,
		_w4278_
	);
	LUT2 #(
		.INIT('h8)
	) name4245 (
		_w4275_,
		_w4278_,
		_w4279_
	);
	LUT3 #(
		.INIT('h37)
	) name4246 (
		_w38_,
		_w39_,
		_w44_,
		_w4280_
	);
	LUT4 #(
		.INIT('h8000)
	) name4247 (
		_w148_,
		_w790_,
		_w978_,
		_w4280_,
		_w4281_
	);
	LUT4 #(
		.INIT('h153f)
	) name4248 (
		_w47_,
		_w50_,
		_w43_,
		_w176_,
		_w4282_
	);
	LUT4 #(
		.INIT('h135f)
	) name4249 (
		_w85_,
		_w44_,
		_w236_,
		_w166_,
		_w4283_
	);
	LUT4 #(
		.INIT('h135f)
	) name4250 (
		_w38_,
		_w65_,
		_w259_,
		_w176_,
		_w4284_
	);
	LUT4 #(
		.INIT('h8000)
	) name4251 (
		_w720_,
		_w4282_,
		_w4283_,
		_w4284_,
		_w4285_
	);
	LUT3 #(
		.INIT('h10)
	) name4252 (
		_w397_,
		_w462_,
		_w1360_,
		_w4286_
	);
	LUT4 #(
		.INIT('h8000)
	) name4253 (
		_w1154_,
		_w1191_,
		_w1587_,
		_w2072_,
		_w4287_
	);
	LUT4 #(
		.INIT('h8000)
	) name4254 (
		_w4286_,
		_w4287_,
		_w4281_,
		_w4285_,
		_w4288_
	);
	LUT4 #(
		.INIT('h8000)
	) name4255 (
		_w1488_,
		_w1499_,
		_w4279_,
		_w4288_,
		_w4289_
	);
	LUT2 #(
		.INIT('h8)
	) name4256 (
		_w4274_,
		_w4289_,
		_w4290_
	);
	LUT4 #(
		.INIT('h0045)
	) name4257 (
		_w4257_,
		_w4259_,
		_w4263_,
		_w4290_,
		_w4291_
	);
	LUT4 #(
		.INIT('hba00)
	) name4258 (
		_w4257_,
		_w4259_,
		_w4263_,
		_w4290_,
		_w4292_
	);
	LUT4 #(
		.INIT('h6659)
	) name4259 (
		_w2157_,
		_w2214_,
		_w2263_,
		_w2294_,
		_w4293_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4260 (
		_w2193_,
		_w2183_,
		_w2213_,
		_w2407_,
		_w4294_
	);
	LUT3 #(
		.INIT('h70)
	) name4261 (
		_w2155_,
		_w2156_,
		_w2527_,
		_w4295_
	);
	LUT3 #(
		.INIT('h2a)
	) name4262 (
		_w376_,
		_w2273_,
		_w2293_,
		_w4296_
	);
	LUT3 #(
		.INIT('h01)
	) name4263 (
		_w4294_,
		_w4295_,
		_w4296_,
		_w4297_
	);
	LUT3 #(
		.INIT('h70)
	) name4264 (
		_w377_,
		_w4293_,
		_w4297_,
		_w4298_
	);
	LUT3 #(
		.INIT('h54)
	) name4265 (
		_w4291_,
		_w4292_,
		_w4298_,
		_w4299_
	);
	LUT2 #(
		.INIT('h8)
	) name4266 (
		_w4236_,
		_w4241_,
		_w4300_
	);
	LUT2 #(
		.INIT('h6)
	) name4267 (
		_w4236_,
		_w4241_,
		_w4301_
	);
	LUT4 #(
		.INIT('h93cc)
	) name4268 (
		_w377_,
		_w4208_,
		_w4209_,
		_w4213_,
		_w4302_
	);
	LUT4 #(
		.INIT('h1700)
	) name4269 (
		_w4236_,
		_w4241_,
		_w4299_,
		_w4302_,
		_w4303_
	);
	LUT2 #(
		.INIT('h8)
	) name4270 (
		_w4175_,
		_w4180_,
		_w4304_
	);
	LUT2 #(
		.INIT('h6)
	) name4271 (
		_w4175_,
		_w4180_,
		_w4305_
	);
	LUT4 #(
		.INIT('h5501)
	) name4272 (
		_w4181_,
		_w4214_,
		_w4303_,
		_w4304_,
		_w4306_
	);
	LUT4 #(
		.INIT('h4c00)
	) name4273 (
		_w377_,
		_w4150_,
		_w4151_,
		_w4155_,
		_w4307_
	);
	LUT4 #(
		.INIT('h93cc)
	) name4274 (
		_w377_,
		_w4150_,
		_w4151_,
		_w4155_,
		_w4308_
	);
	LUT3 #(
		.INIT('h54)
	) name4275 (
		_w4157_,
		_w4306_,
		_w4307_,
		_w4309_
	);
	LUT2 #(
		.INIT('h9)
	) name4276 (
		_w3961_,
		_w3966_,
		_w4310_
	);
	LUT4 #(
		.INIT('h1700)
	) name4277 (
		_w4150_,
		_w4156_,
		_w4306_,
		_w4310_,
		_w4311_
	);
	LUT4 #(
		.INIT('h00e8)
	) name4278 (
		_w4150_,
		_w4156_,
		_w4306_,
		_w4310_,
		_w4312_
	);
	LUT4 #(
		.INIT('h54ab)
	) name4279 (
		_w4157_,
		_w4306_,
		_w4307_,
		_w4310_,
		_w4313_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4280 (
		_w1817_,
		_w1799_,
		_w1840_,
		_w2854_,
		_w4314_
	);
	LUT3 #(
		.INIT('h70)
	) name4281 (
		_w1898_,
		_w1928_,
		_w2549_,
		_w4315_
	);
	LUT3 #(
		.INIT('h70)
	) name4282 (
		_w1863_,
		_w1875_,
		_w2617_,
		_w4316_
	);
	LUT3 #(
		.INIT('h01)
	) name4283 (
		_w4315_,
		_w4316_,
		_w4314_,
		_w4317_
	);
	LUT4 #(
		.INIT('h95aa)
	) name4284 (
		\a[29] ,
		_w2550_,
		_w3972_,
		_w4317_,
		_w4318_
	);
	LUT2 #(
		.INIT('h9)
	) name4285 (
		_w4125_,
		_w4131_,
		_w4319_
	);
	LUT4 #(
		.INIT('h4d00)
	) name4286 (
		_w4309_,
		_w4310_,
		_w4318_,
		_w4319_,
		_w4320_
	);
	LUT3 #(
		.INIT('h96)
	) name4287 (
		_w3967_,
		_w3968_,
		_w4123_,
		_w4321_
	);
	LUT4 #(
		.INIT('h0155)
	) name4288 (
		_w4124_,
		_w4132_,
		_w4320_,
		_w4321_,
		_w4322_
	);
	LUT4 #(
		.INIT('hd42b)
	) name4289 (
		\a[2] ,
		_w3931_,
		_w3967_,
		_w3969_,
		_w4323_
	);
	LUT2 #(
		.INIT('h9)
	) name4290 (
		_w3977_,
		_w4323_,
		_w4324_
	);
	LUT3 #(
		.INIT('h70)
	) name4291 (
		_w1692_,
		_w1723_,
		_w2854_,
		_w4325_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4292 (
		_w1751_,
		_w1742_,
		_w1771_,
		_w2617_,
		_w4326_
	);
	LUT3 #(
		.INIT('h70)
	) name4293 (
		_w1795_,
		_w1796_,
		_w2549_,
		_w4327_
	);
	LUT3 #(
		.INIT('h01)
	) name4294 (
		_w4326_,
		_w4327_,
		_w4325_,
		_w4328_
	);
	LUT4 #(
		.INIT('h6f00)
	) name4295 (
		_w2315_,
		_w2317_,
		_w2550_,
		_w4328_,
		_w4329_
	);
	LUT2 #(
		.INIT('h6)
	) name4296 (
		\a[29] ,
		_w4329_,
		_w4330_
	);
	LUT3 #(
		.INIT('hb2)
	) name4297 (
		_w4322_,
		_w4324_,
		_w4330_,
		_w4331_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4298 (
		_w1454_,
		_w1426_,
		_w1478_,
		_w2986_,
		_w4332_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4299 (
		_w1584_,
		_w1569_,
		_w1606_,
		_w2874_,
		_w4333_
	);
	LUT3 #(
		.INIT('h70)
	) name4300 (
		_w1501_,
		_w1545_,
		_w2975_,
		_w4334_
	);
	LUT3 #(
		.INIT('h01)
	) name4301 (
		_w4333_,
		_w4334_,
		_w4332_,
		_w4335_
	);
	LUT4 #(
		.INIT('h6f00)
	) name4302 (
		_w2323_,
		_w2325_,
		_w2875_,
		_w4335_,
		_w4336_
	);
	LUT4 #(
		.INIT('h71b2)
	) name4303 (
		\a[26] ,
		_w4118_,
		_w4331_,
		_w4336_,
		_w4337_
	);
	LUT3 #(
		.INIT('h09)
	) name4304 (
		_w4065_,
		_w4117_,
		_w4337_,
		_w4338_
	);
	LUT3 #(
		.INIT('h60)
	) name4305 (
		_w4065_,
		_w4117_,
		_w4337_,
		_w4339_
	);
	LUT3 #(
		.INIT('h70)
	) name4306 (
		_w1202_,
		_w1233_,
		_w3262_,
		_w4340_
	);
	LUT3 #(
		.INIT('h2a)
	) name4307 (
		_w3214_,
		_w1325_,
		_w1367_,
		_w4341_
	);
	LUT3 #(
		.INIT('h70)
	) name4308 (
		_w1253_,
		_w1294_,
		_w3249_,
		_w4342_
	);
	LUT3 #(
		.INIT('h01)
	) name4309 (
		_w4341_,
		_w4342_,
		_w4340_,
		_w4343_
	);
	LUT4 #(
		.INIT('h6f00)
	) name4310 (
		_w2331_,
		_w2333_,
		_w37_,
		_w4343_,
		_w4344_
	);
	LUT4 #(
		.INIT('h3132)
	) name4311 (
		\a[23] ,
		_w4338_,
		_w4339_,
		_w4344_,
		_w4345_
	);
	LUT3 #(
		.INIT('hb2)
	) name4312 (
		_w4115_,
		_w4116_,
		_w4345_,
		_w4346_
	);
	LUT4 #(
		.INIT('h9669)
	) name4313 (
		\a[23] ,
		_w4067_,
		_w4069_,
		_w4074_,
		_w4347_
	);
	LUT2 #(
		.INIT('h1)
	) name4314 (
		_w4346_,
		_w4347_,
		_w4348_
	);
	LUT2 #(
		.INIT('h8)
	) name4315 (
		_w4346_,
		_w4347_,
		_w4349_
	);
	LUT3 #(
		.INIT('h70)
	) name4316 (
		_w1009_,
		_w1050_,
		_w3311_,
		_w4350_
	);
	LUT3 #(
		.INIT('h70)
	) name4317 (
		_w871_,
		_w927_,
		_w3654_,
		_w4351_
	);
	LUT3 #(
		.INIT('h70)
	) name4318 (
		_w763_,
		_w983_,
		_w3645_,
		_w4352_
	);
	LUT3 #(
		.INIT('h01)
	) name4319 (
		_w4351_,
		_w4352_,
		_w4350_,
		_w4353_
	);
	LUT4 #(
		.INIT('h95aa)
	) name4320 (
		\a[20] ,
		_w2839_,
		_w3312_,
		_w4353_,
		_w4354_
	);
	LUT3 #(
		.INIT('h54)
	) name4321 (
		_w4348_,
		_w4349_,
		_w4354_,
		_w4355_
	);
	LUT2 #(
		.INIT('h2)
	) name4322 (
		_w4110_,
		_w4355_,
		_w4356_
	);
	LUT2 #(
		.INIT('h4)
	) name4323 (
		_w4110_,
		_w4355_,
		_w4357_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4324 (
		_w587_,
		_w608_,
		_w624_,
		_w3886_,
		_w4358_
	);
	LUT3 #(
		.INIT('h70)
	) name4325 (
		_w725_,
		_w764_,
		_w3709_,
		_w4359_
	);
	LUT3 #(
		.INIT('h70)
	) name4326 (
		_w666_,
		_w694_,
		_w3877_,
		_w4360_
	);
	LUT3 #(
		.INIT('h01)
	) name4327 (
		_w4359_,
		_w4360_,
		_w4358_,
		_w4361_
	);
	LUT4 #(
		.INIT('h95aa)
	) name4328 (
		\a[17] ,
		_w2598_,
		_w3710_,
		_w4361_,
		_w4362_
	);
	LUT3 #(
		.INIT('h54)
	) name4329 (
		_w4356_,
		_w4357_,
		_w4362_,
		_w4363_
	);
	LUT3 #(
		.INIT('h54)
	) name4330 (
		_w4106_,
		_w4107_,
		_w4363_,
		_w4364_
	);
	LUT4 #(
		.INIT('hf400)
	) name4331 (
		_w374_,
		_w2361_,
		_w2404_,
		_w4034_,
		_w4365_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4332 (
		_w121_,
		_w418_,
		_w422_,
		_w4033_,
		_w4366_
	);
	LUT3 #(
		.INIT('h18)
	) name4333 (
		\a[11] ,
		\a[12] ,
		\a[13] ,
		_w4367_
	);
	LUT3 #(
		.INIT('h70)
	) name4334 (
		_w352_,
		_w373_,
		_w4367_,
		_w4368_
	);
	LUT2 #(
		.INIT('h1)
	) name4335 (
		_w4366_,
		_w4368_,
		_w4369_
	);
	LUT3 #(
		.INIT('h9a)
	) name4336 (
		\a[14] ,
		_w4365_,
		_w4369_,
		_w4370_
	);
	LUT4 #(
		.INIT('h1211)
	) name4337 (
		\a[14] ,
		_w4364_,
		_w4365_,
		_w4369_,
		_w4371_
	);
	LUT4 #(
		.INIT('h8488)
	) name4338 (
		\a[14] ,
		_w4364_,
		_w4365_,
		_w4369_,
		_w4372_
	);
	LUT4 #(
		.INIT('h6966)
	) name4339 (
		\a[14] ,
		_w4364_,
		_w4365_,
		_w4369_,
		_w4373_
	);
	LUT2 #(
		.INIT('h9)
	) name4340 (
		_w4084_,
		_w4085_,
		_w4374_
	);
	LUT2 #(
		.INIT('h6)
	) name4341 (
		_w4092_,
		_w4374_,
		_w4375_
	);
	LUT3 #(
		.INIT('h54)
	) name4342 (
		_w4371_,
		_w4372_,
		_w4375_,
		_w4376_
	);
	LUT4 #(
		.INIT('h9669)
	) name4343 (
		\a[14] ,
		_w4035_,
		_w4093_,
		_w4095_,
		_w4377_
	);
	LUT4 #(
		.INIT('h1700)
	) name4344 (
		_w4364_,
		_w4370_,
		_w4375_,
		_w4377_,
		_w4378_
	);
	LUT4 #(
		.INIT('h54ab)
	) name4345 (
		_w4371_,
		_w4372_,
		_w4375_,
		_w4377_,
		_w4379_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4346 (
		_w486_,
		_w487_,
		_w509_,
		_w4033_,
		_w4380_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4347 (
		_w121_,
		_w418_,
		_w422_,
		_w4367_,
		_w4381_
	);
	LUT4 #(
		.INIT('h6006)
	) name4348 (
		\a[11] ,
		\a[12] ,
		\a[13] ,
		\a[14] ,
		_w4382_
	);
	LUT3 #(
		.INIT('h70)
	) name4349 (
		_w352_,
		_w373_,
		_w4382_,
		_w4383_
	);
	LUT3 #(
		.INIT('h01)
	) name4350 (
		_w4380_,
		_w4381_,
		_w4383_,
		_w4384_
	);
	LUT4 #(
		.INIT('h95aa)
	) name4351 (
		\a[14] ,
		_w2535_,
		_w4034_,
		_w4384_,
		_w4385_
	);
	LUT2 #(
		.INIT('h9)
	) name4352 (
		_w4110_,
		_w4355_,
		_w4386_
	);
	LUT3 #(
		.INIT('h96)
	) name4353 (
		_w4115_,
		_w4116_,
		_w4345_,
		_w4387_
	);
	LUT3 #(
		.INIT('h70)
	) name4354 (
		_w1071_,
		_w1102_,
		_w3311_,
		_w4388_
	);
	LUT3 #(
		.INIT('h70)
	) name4355 (
		_w763_,
		_w983_,
		_w3654_,
		_w4389_
	);
	LUT3 #(
		.INIT('h70)
	) name4356 (
		_w1009_,
		_w1050_,
		_w3645_,
		_w4390_
	);
	LUT3 #(
		.INIT('h01)
	) name4357 (
		_w4389_,
		_w4390_,
		_w4388_,
		_w4391_
	);
	LUT4 #(
		.INIT('h6f00)
	) name4358 (
		_w2339_,
		_w2341_,
		_w3312_,
		_w4391_,
		_w4392_
	);
	LUT3 #(
		.INIT('h84)
	) name4359 (
		\a[20] ,
		_w4387_,
		_w4392_,
		_w4393_
	);
	LUT3 #(
		.INIT('h12)
	) name4360 (
		\a[20] ,
		_w4387_,
		_w4392_,
		_w4394_
	);
	LUT3 #(
		.INIT('h69)
	) name4361 (
		\a[20] ,
		_w4387_,
		_w4392_,
		_w4395_
	);
	LUT3 #(
		.INIT('h96)
	) name4362 (
		_w4065_,
		_w4117_,
		_w4337_,
		_w4396_
	);
	LUT3 #(
		.INIT('h69)
	) name4363 (
		\a[23] ,
		_w4344_,
		_w4396_,
		_w4397_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4364 (
		_w1584_,
		_w1569_,
		_w1606_,
		_w2975_,
		_w4398_
	);
	LUT3 #(
		.INIT('h70)
	) name4365 (
		_w1501_,
		_w1545_,
		_w2986_,
		_w4399_
	);
	LUT3 #(
		.INIT('h70)
	) name4366 (
		_w1620_,
		_w1661_,
		_w2874_,
		_w4400_
	);
	LUT3 #(
		.INIT('h01)
	) name4367 (
		_w4398_,
		_w4399_,
		_w4400_,
		_w4401_
	);
	LUT4 #(
		.INIT('h95aa)
	) name4368 (
		\a[26] ,
		_w2875_,
		_w3495_,
		_w4401_,
		_w4402_
	);
	LUT3 #(
		.INIT('h69)
	) name4369 (
		_w4322_,
		_w4324_,
		_w4330_,
		_w4403_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4370 (
		_w1751_,
		_w1742_,
		_w1771_,
		_w2854_,
		_w4404_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4371 (
		_w1817_,
		_w1799_,
		_w1840_,
		_w2549_,
		_w4405_
	);
	LUT3 #(
		.INIT('h70)
	) name4372 (
		_w1795_,
		_w1796_,
		_w2617_,
		_w4406_
	);
	LUT3 #(
		.INIT('h01)
	) name4373 (
		_w4405_,
		_w4406_,
		_w4404_,
		_w4407_
	);
	LUT4 #(
		.INIT('h95aa)
	) name4374 (
		\a[29] ,
		_w2550_,
		_w3909_,
		_w4407_,
		_w4408_
	);
	LUT4 #(
		.INIT('h001e)
	) name4375 (
		_w4132_,
		_w4320_,
		_w4321_,
		_w4408_,
		_w4409_
	);
	LUT4 #(
		.INIT('he100)
	) name4376 (
		_w4132_,
		_w4320_,
		_w4321_,
		_w4408_,
		_w4410_
	);
	LUT3 #(
		.INIT('h70)
	) name4377 (
		_w1692_,
		_w1723_,
		_w2874_,
		_w4411_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4378 (
		_w1584_,
		_w1569_,
		_w1606_,
		_w2986_,
		_w4412_
	);
	LUT3 #(
		.INIT('h70)
	) name4379 (
		_w1620_,
		_w1661_,
		_w2975_,
		_w4413_
	);
	LUT3 #(
		.INIT('h01)
	) name4380 (
		_w4412_,
		_w4413_,
		_w4411_,
		_w4414_
	);
	LUT4 #(
		.INIT('h6f00)
	) name4381 (
		_w2319_,
		_w2321_,
		_w2875_,
		_w4414_,
		_w4415_
	);
	LUT4 #(
		.INIT('h3132)
	) name4382 (
		\a[26] ,
		_w4409_,
		_w4410_,
		_w4415_,
		_w4416_
	);
	LUT3 #(
		.INIT('he8)
	) name4383 (
		_w4402_,
		_w4403_,
		_w4416_,
		_w4417_
	);
	LUT4 #(
		.INIT('h6996)
	) name4384 (
		\a[26] ,
		_w4118_,
		_w4331_,
		_w4336_,
		_w4418_
	);
	LUT2 #(
		.INIT('h4)
	) name4385 (
		_w4417_,
		_w4418_,
		_w4419_
	);
	LUT2 #(
		.INIT('h2)
	) name4386 (
		_w4417_,
		_w4418_,
		_w4420_
	);
	LUT3 #(
		.INIT('h2a)
	) name4387 (
		_w3214_,
		_w1381_,
		_w1398_,
		_w4421_
	);
	LUT3 #(
		.INIT('h70)
	) name4388 (
		_w1325_,
		_w1367_,
		_w3249_,
		_w4422_
	);
	LUT3 #(
		.INIT('h70)
	) name4389 (
		_w1253_,
		_w1294_,
		_w3262_,
		_w4423_
	);
	LUT3 #(
		.INIT('h01)
	) name4390 (
		_w4422_,
		_w4423_,
		_w4421_,
		_w4424_
	);
	LUT4 #(
		.INIT('h95aa)
	) name4391 (
		\a[23] ,
		_w3182_,
		_w37_,
		_w4424_,
		_w4425_
	);
	LUT3 #(
		.INIT('h54)
	) name4392 (
		_w4419_,
		_w4420_,
		_w4425_,
		_w4426_
	);
	LUT2 #(
		.INIT('h2)
	) name4393 (
		_w4397_,
		_w4426_,
		_w4427_
	);
	LUT2 #(
		.INIT('h4)
	) name4394 (
		_w4397_,
		_w4426_,
		_w4428_
	);
	LUT3 #(
		.INIT('h70)
	) name4395 (
		_w1136_,
		_w1187_,
		_w3311_,
		_w4429_
	);
	LUT3 #(
		.INIT('h70)
	) name4396 (
		_w1009_,
		_w1050_,
		_w3654_,
		_w4430_
	);
	LUT3 #(
		.INIT('h70)
	) name4397 (
		_w1071_,
		_w1102_,
		_w3645_,
		_w4431_
	);
	LUT3 #(
		.INIT('h01)
	) name4398 (
		_w4430_,
		_w4431_,
		_w4429_,
		_w4432_
	);
	LUT4 #(
		.INIT('h95aa)
	) name4399 (
		\a[20] ,
		_w2936_,
		_w3312_,
		_w4432_,
		_w4433_
	);
	LUT3 #(
		.INIT('h54)
	) name4400 (
		_w4427_,
		_w4428_,
		_w4433_,
		_w4434_
	);
	LUT3 #(
		.INIT('h54)
	) name4401 (
		_w4393_,
		_w4394_,
		_w4434_,
		_w4435_
	);
	LUT2 #(
		.INIT('h6)
	) name4402 (
		_w4346_,
		_w4347_,
		_w4436_
	);
	LUT2 #(
		.INIT('h9)
	) name4403 (
		_w4354_,
		_w4436_,
		_w4437_
	);
	LUT3 #(
		.INIT('h70)
	) name4404 (
		_w725_,
		_w764_,
		_w3877_,
		_w4438_
	);
	LUT3 #(
		.INIT('h70)
	) name4405 (
		_w801_,
		_w851_,
		_w3709_,
		_w4439_
	);
	LUT3 #(
		.INIT('h70)
	) name4406 (
		_w666_,
		_w694_,
		_w3886_,
		_w4440_
	);
	LUT3 #(
		.INIT('h01)
	) name4407 (
		_w4439_,
		_w4440_,
		_w4438_,
		_w4441_
	);
	LUT4 #(
		.INIT('h6f00)
	) name4408 (
		_w2347_,
		_w2349_,
		_w3710_,
		_w4441_,
		_w4442_
	);
	LUT4 #(
		.INIT('h4d8e)
	) name4409 (
		\a[17] ,
		_w4435_,
		_w4437_,
		_w4442_,
		_w4443_
	);
	LUT3 #(
		.INIT('h09)
	) name4410 (
		_w4362_,
		_w4386_,
		_w4443_,
		_w4444_
	);
	LUT3 #(
		.INIT('h60)
	) name4411 (
		_w4362_,
		_w4386_,
		_w4443_,
		_w4445_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4412 (
		_w486_,
		_w487_,
		_w509_,
		_w4367_,
		_w4446_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4413 (
		_w121_,
		_w418_,
		_w422_,
		_w4382_,
		_w4447_
	);
	LUT3 #(
		.INIT('h70)
	) name4414 (
		_w544_,
		_w558_,
		_w4033_,
		_w4448_
	);
	LUT3 #(
		.INIT('h01)
	) name4415 (
		_w4446_,
		_w4447_,
		_w4448_,
		_w4449_
	);
	LUT4 #(
		.INIT('h6f00)
	) name4416 (
		_w2355_,
		_w2357_,
		_w4034_,
		_w4449_,
		_w4450_
	);
	LUT4 #(
		.INIT('h3132)
	) name4417 (
		\a[14] ,
		_w4444_,
		_w4445_,
		_w4450_,
		_w4451_
	);
	LUT2 #(
		.INIT('h9)
	) name4418 (
		_w4108_,
		_w4363_,
		_w4452_
	);
	LUT3 #(
		.INIT('h8e)
	) name4419 (
		_w4385_,
		_w4451_,
		_w4452_,
		_w4453_
	);
	LUT2 #(
		.INIT('h9)
	) name4420 (
		_w4373_,
		_w4375_,
		_w4454_
	);
	LUT3 #(
		.INIT('h09)
	) name4421 (
		_w4373_,
		_w4375_,
		_w4453_,
		_w4455_
	);
	LUT3 #(
		.INIT('h96)
	) name4422 (
		_w4385_,
		_w4451_,
		_w4452_,
		_w4456_
	);
	LUT2 #(
		.INIT('h9)
	) name4423 (
		\a[8] ,
		\a[9] ,
		_w4457_
	);
	LUT4 #(
		.INIT('h0180)
	) name4424 (
		\a[8] ,
		\a[9] ,
		\a[10] ,
		\a[11] ,
		_w4458_
	);
	LUT4 #(
		.INIT('h0660)
	) name4425 (
		\a[8] ,
		\a[9] ,
		\a[10] ,
		\a[11] ,
		_w4459_
	);
	LUT4 #(
		.INIT('h5150)
	) name4426 (
		_w374_,
		_w2361_,
		_w4458_,
		_w4459_,
		_w4460_
	);
	LUT3 #(
		.INIT('h70)
	) name4427 (
		_w725_,
		_w764_,
		_w3886_,
		_w4461_
	);
	LUT3 #(
		.INIT('h70)
	) name4428 (
		_w801_,
		_w851_,
		_w3877_,
		_w4462_
	);
	LUT3 #(
		.INIT('h70)
	) name4429 (
		_w871_,
		_w927_,
		_w3709_,
		_w4463_
	);
	LUT3 #(
		.INIT('h01)
	) name4430 (
		_w4462_,
		_w4463_,
		_w4461_,
		_w4464_
	);
	LUT4 #(
		.INIT('h95aa)
	) name4431 (
		\a[17] ,
		_w2724_,
		_w3710_,
		_w4464_,
		_w4465_
	);
	LUT2 #(
		.INIT('h9)
	) name4432 (
		_w4395_,
		_w4434_,
		_w4466_
	);
	LUT2 #(
		.INIT('h9)
	) name4433 (
		_w4397_,
		_w4426_,
		_w4467_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name4434 (
		_w3214_,
		_w1454_,
		_w1426_,
		_w1478_,
		_w4468_
	);
	LUT3 #(
		.INIT('h70)
	) name4435 (
		_w1325_,
		_w1367_,
		_w3262_,
		_w4469_
	);
	LUT3 #(
		.INIT('h70)
	) name4436 (
		_w1381_,
		_w1398_,
		_w3249_,
		_w4470_
	);
	LUT3 #(
		.INIT('h01)
	) name4437 (
		_w4469_,
		_w4470_,
		_w4468_,
		_w4471_
	);
	LUT4 #(
		.INIT('h6f00)
	) name4438 (
		_w2327_,
		_w2329_,
		_w37_,
		_w4471_,
		_w4472_
	);
	LUT3 #(
		.INIT('h69)
	) name4439 (
		_w4402_,
		_w4403_,
		_w4416_,
		_w4473_
	);
	LUT3 #(
		.INIT('h90)
	) name4440 (
		\a[23] ,
		_w4472_,
		_w4473_,
		_w4474_
	);
	LUT3 #(
		.INIT('h06)
	) name4441 (
		\a[23] ,
		_w4472_,
		_w4473_,
		_w4475_
	);
	LUT3 #(
		.INIT('h69)
	) name4442 (
		\a[23] ,
		_w4472_,
		_w4473_,
		_w4476_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name4443 (
		_w4132_,
		_w4320_,
		_w4321_,
		_w4408_,
		_w4477_
	);
	LUT3 #(
		.INIT('h69)
	) name4444 (
		\a[26] ,
		_w4415_,
		_w4477_,
		_w4478_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4445 (
		_w1817_,
		_w1799_,
		_w1840_,
		_w2617_,
		_w4479_
	);
	LUT3 #(
		.INIT('h70)
	) name4446 (
		_w1795_,
		_w1796_,
		_w2854_,
		_w4480_
	);
	LUT3 #(
		.INIT('h70)
	) name4447 (
		_w1863_,
		_w1875_,
		_w2549_,
		_w4481_
	);
	LUT3 #(
		.INIT('h01)
	) name4448 (
		_w4480_,
		_w4481_,
		_w4479_,
		_w4482_
	);
	LUT4 #(
		.INIT('h6f00)
	) name4449 (
		_w2311_,
		_w2313_,
		_w2550_,
		_w4482_,
		_w4483_
	);
	LUT2 #(
		.INIT('h6)
	) name4450 (
		\a[29] ,
		_w4483_,
		_w4484_
	);
	LUT4 #(
		.INIT('h54ab)
	) name4451 (
		_w4311_,
		_w4312_,
		_w4318_,
		_w4319_,
		_w4485_
	);
	LUT2 #(
		.INIT('h4)
	) name4452 (
		_w4484_,
		_w4485_,
		_w4486_
	);
	LUT2 #(
		.INIT('h2)
	) name4453 (
		_w4484_,
		_w4485_,
		_w4487_
	);
	LUT3 #(
		.INIT('h70)
	) name4454 (
		_w1692_,
		_w1723_,
		_w2975_,
		_w4488_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4455 (
		_w1751_,
		_w1742_,
		_w1771_,
		_w2874_,
		_w4489_
	);
	LUT3 #(
		.INIT('h70)
	) name4456 (
		_w1620_,
		_w1661_,
		_w2986_,
		_w4490_
	);
	LUT3 #(
		.INIT('h01)
	) name4457 (
		_w4489_,
		_w4490_,
		_w4488_,
		_w4491_
	);
	LUT4 #(
		.INIT('h95aa)
	) name4458 (
		\a[26] ,
		_w2875_,
		_w3599_,
		_w4491_,
		_w4492_
	);
	LUT3 #(
		.INIT('h54)
	) name4459 (
		_w4486_,
		_w4487_,
		_w4492_,
		_w4493_
	);
	LUT2 #(
		.INIT('h2)
	) name4460 (
		_w4478_,
		_w4493_,
		_w4494_
	);
	LUT2 #(
		.INIT('h4)
	) name4461 (
		_w4478_,
		_w4493_,
		_w4495_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4462 (
		_w1454_,
		_w1426_,
		_w1478_,
		_w3249_,
		_w4496_
	);
	LUT3 #(
		.INIT('h70)
	) name4463 (
		_w1381_,
		_w1398_,
		_w3262_,
		_w4497_
	);
	LUT3 #(
		.INIT('h2a)
	) name4464 (
		_w3214_,
		_w1501_,
		_w1545_,
		_w4498_
	);
	LUT3 #(
		.INIT('h01)
	) name4465 (
		_w4497_,
		_w4498_,
		_w4496_,
		_w4499_
	);
	LUT4 #(
		.INIT('h95aa)
	) name4466 (
		\a[23] ,
		_w37_,
		_w3362_,
		_w4499_,
		_w4500_
	);
	LUT3 #(
		.INIT('h54)
	) name4467 (
		_w4494_,
		_w4495_,
		_w4500_,
		_w4501_
	);
	LUT3 #(
		.INIT('h54)
	) name4468 (
		_w4474_,
		_w4475_,
		_w4501_,
		_w4502_
	);
	LUT2 #(
		.INIT('h9)
	) name4469 (
		_w4417_,
		_w4418_,
		_w4503_
	);
	LUT2 #(
		.INIT('h6)
	) name4470 (
		_w4425_,
		_w4503_,
		_w4504_
	);
	LUT3 #(
		.INIT('h70)
	) name4471 (
		_w1136_,
		_w1187_,
		_w3645_,
		_w4505_
	);
	LUT3 #(
		.INIT('h70)
	) name4472 (
		_w1071_,
		_w1102_,
		_w3654_,
		_w4506_
	);
	LUT3 #(
		.INIT('h70)
	) name4473 (
		_w1202_,
		_w1233_,
		_w3311_,
		_w4507_
	);
	LUT3 #(
		.INIT('h01)
	) name4474 (
		_w4506_,
		_w4507_,
		_w4505_,
		_w4508_
	);
	LUT4 #(
		.INIT('h6f00)
	) name4475 (
		_w2335_,
		_w2337_,
		_w3312_,
		_w4508_,
		_w4509_
	);
	LUT4 #(
		.INIT('hd4e8)
	) name4476 (
		\a[20] ,
		_w4502_,
		_w4504_,
		_w4509_,
		_w4510_
	);
	LUT3 #(
		.INIT('h09)
	) name4477 (
		_w4433_,
		_w4467_,
		_w4510_,
		_w4511_
	);
	LUT3 #(
		.INIT('h60)
	) name4478 (
		_w4433_,
		_w4467_,
		_w4510_,
		_w4512_
	);
	LUT3 #(
		.INIT('h70)
	) name4479 (
		_w763_,
		_w983_,
		_w3709_,
		_w4513_
	);
	LUT3 #(
		.INIT('h70)
	) name4480 (
		_w871_,
		_w927_,
		_w3877_,
		_w4514_
	);
	LUT3 #(
		.INIT('h70)
	) name4481 (
		_w801_,
		_w851_,
		_w3886_,
		_w4515_
	);
	LUT3 #(
		.INIT('h01)
	) name4482 (
		_w4514_,
		_w4515_,
		_w4513_,
		_w4516_
	);
	LUT4 #(
		.INIT('h6f00)
	) name4483 (
		_w2343_,
		_w2345_,
		_w3710_,
		_w4516_,
		_w4517_
	);
	LUT4 #(
		.INIT('h3132)
	) name4484 (
		\a[17] ,
		_w4511_,
		_w4512_,
		_w4517_,
		_w4518_
	);
	LUT3 #(
		.INIT('hb2)
	) name4485 (
		_w4465_,
		_w4466_,
		_w4518_,
		_w4519_
	);
	LUT4 #(
		.INIT('h9669)
	) name4486 (
		\a[17] ,
		_w4435_,
		_w4437_,
		_w4442_,
		_w4520_
	);
	LUT2 #(
		.INIT('h1)
	) name4487 (
		_w4519_,
		_w4520_,
		_w4521_
	);
	LUT2 #(
		.INIT('h8)
	) name4488 (
		_w4519_,
		_w4520_,
		_w4522_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4489 (
		_w486_,
		_w487_,
		_w509_,
		_w4382_,
		_w4523_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4490 (
		_w587_,
		_w608_,
		_w624_,
		_w4033_,
		_w4524_
	);
	LUT3 #(
		.INIT('h70)
	) name4491 (
		_w544_,
		_w558_,
		_w4367_,
		_w4525_
	);
	LUT3 #(
		.INIT('h01)
	) name4492 (
		_w4523_,
		_w4524_,
		_w4525_,
		_w4526_
	);
	LUT4 #(
		.INIT('h95aa)
	) name4493 (
		\a[14] ,
		_w2526_,
		_w4034_,
		_w4526_,
		_w4527_
	);
	LUT3 #(
		.INIT('h54)
	) name4494 (
		_w4521_,
		_w4522_,
		_w4527_,
		_w4528_
	);
	LUT3 #(
		.INIT('h96)
	) name4495 (
		_w4362_,
		_w4386_,
		_w4443_,
		_w4529_
	);
	LUT3 #(
		.INIT('h69)
	) name4496 (
		\a[14] ,
		_w4450_,
		_w4529_,
		_w4530_
	);
	LUT4 #(
		.INIT('h90f9)
	) name4497 (
		\a[11] ,
		_w4460_,
		_w4528_,
		_w4530_,
		_w4531_
	);
	LUT2 #(
		.INIT('h2)
	) name4498 (
		_w4456_,
		_w4531_,
		_w4532_
	);
	LUT3 #(
		.INIT('h96)
	) name4499 (
		_w4465_,
		_w4466_,
		_w4518_,
		_w4533_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4500 (
		_w587_,
		_w608_,
		_w624_,
		_w4367_,
		_w4534_
	);
	LUT3 #(
		.INIT('h70)
	) name4501 (
		_w666_,
		_w694_,
		_w4033_,
		_w4535_
	);
	LUT3 #(
		.INIT('h70)
	) name4502 (
		_w544_,
		_w558_,
		_w4382_,
		_w4536_
	);
	LUT3 #(
		.INIT('h01)
	) name4503 (
		_w4535_,
		_w4536_,
		_w4534_,
		_w4537_
	);
	LUT4 #(
		.INIT('h6f00)
	) name4504 (
		_w2351_,
		_w2353_,
		_w4034_,
		_w4537_,
		_w4538_
	);
	LUT3 #(
		.INIT('h84)
	) name4505 (
		\a[14] ,
		_w4533_,
		_w4538_,
		_w4539_
	);
	LUT3 #(
		.INIT('h12)
	) name4506 (
		\a[14] ,
		_w4533_,
		_w4538_,
		_w4540_
	);
	LUT3 #(
		.INIT('h69)
	) name4507 (
		\a[14] ,
		_w4533_,
		_w4538_,
		_w4541_
	);
	LUT3 #(
		.INIT('h96)
	) name4508 (
		_w4433_,
		_w4467_,
		_w4510_,
		_w4542_
	);
	LUT3 #(
		.INIT('h69)
	) name4509 (
		\a[17] ,
		_w4517_,
		_w4542_,
		_w4543_
	);
	LUT2 #(
		.INIT('h9)
	) name4510 (
		_w4476_,
		_w4501_,
		_w4544_
	);
	LUT3 #(
		.INIT('h70)
	) name4511 (
		_w1202_,
		_w1233_,
		_w3645_,
		_w4545_
	);
	LUT3 #(
		.INIT('h70)
	) name4512 (
		_w1253_,
		_w1294_,
		_w3311_,
		_w4546_
	);
	LUT3 #(
		.INIT('h70)
	) name4513 (
		_w1136_,
		_w1187_,
		_w3654_,
		_w4547_
	);
	LUT3 #(
		.INIT('h01)
	) name4514 (
		_w4546_,
		_w4547_,
		_w4545_,
		_w4548_
	);
	LUT4 #(
		.INIT('h95aa)
	) name4515 (
		\a[20] ,
		_w3067_,
		_w3312_,
		_w4548_,
		_w4549_
	);
	LUT2 #(
		.INIT('h9)
	) name4516 (
		_w4478_,
		_w4493_,
		_w4550_
	);
	LUT3 #(
		.INIT('h70)
	) name4517 (
		_w1501_,
		_w1949_,
		_w2549_,
		_w4551_
	);
	LUT3 #(
		.INIT('h70)
	) name4518 (
		_w1898_,
		_w1928_,
		_w2617_,
		_w4552_
	);
	LUT3 #(
		.INIT('h70)
	) name4519 (
		_w1863_,
		_w1875_,
		_w2854_,
		_w4553_
	);
	LUT3 #(
		.INIT('h01)
	) name4520 (
		_w4552_,
		_w4553_,
		_w4551_,
		_w4554_
	);
	LUT4 #(
		.INIT('h6f00)
	) name4521 (
		_w2307_,
		_w2309_,
		_w2550_,
		_w4554_,
		_w4555_
	);
	LUT4 #(
		.INIT('h8241)
	) name4522 (
		\a[29] ,
		_w4306_,
		_w4308_,
		_w4555_,
		_w4556_
	);
	LUT3 #(
		.INIT('h70)
	) name4523 (
		_w1973_,
		_w1997_,
		_w2549_,
		_w4557_
	);
	LUT3 #(
		.INIT('h70)
	) name4524 (
		_w1898_,
		_w1928_,
		_w2854_,
		_w4558_
	);
	LUT3 #(
		.INIT('h70)
	) name4525 (
		_w1501_,
		_w1949_,
		_w2617_,
		_w4559_
	);
	LUT3 #(
		.INIT('h01)
	) name4526 (
		_w4558_,
		_w4559_,
		_w4557_,
		_w4560_
	);
	LUT4 #(
		.INIT('h95aa)
	) name4527 (
		\a[29] ,
		_w2550_,
		_w4126_,
		_w4560_,
		_w4561_
	);
	LUT3 #(
		.INIT('h1e)
	) name4528 (
		_w4214_,
		_w4303_,
		_w4305_,
		_w4562_
	);
	LUT2 #(
		.INIT('h4)
	) name4529 (
		_w4561_,
		_w4562_,
		_w4563_
	);
	LUT3 #(
		.INIT('h70)
	) name4530 (
		_w1973_,
		_w1997_,
		_w2617_,
		_w4564_
	);
	LUT3 #(
		.INIT('h70)
	) name4531 (
		_w1501_,
		_w1949_,
		_w2854_,
		_w4565_
	);
	LUT3 #(
		.INIT('h70)
	) name4532 (
		_w2023_,
		_w2055_,
		_w2549_,
		_w4566_
	);
	LUT3 #(
		.INIT('h01)
	) name4533 (
		_w4565_,
		_w4566_,
		_w4564_,
		_w4567_
	);
	LUT4 #(
		.INIT('h6f00)
	) name4534 (
		_w2303_,
		_w2305_,
		_w2550_,
		_w4567_,
		_w4568_
	);
	LUT2 #(
		.INIT('h6)
	) name4535 (
		\a[29] ,
		_w4568_,
		_w4569_
	);
	LUT4 #(
		.INIT('h54ab)
	) name4536 (
		_w4242_,
		_w4299_,
		_w4300_,
		_w4302_,
		_w4570_
	);
	LUT3 #(
		.INIT('h90)
	) name4537 (
		\a[29] ,
		_w4568_,
		_w4570_,
		_w4571_
	);
	LUT3 #(
		.INIT('h70)
	) name4538 (
		_w1973_,
		_w1997_,
		_w2854_,
		_w4572_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4539 (
		_w1874_,
		_w2076_,
		_w2099_,
		_w2549_,
		_w4573_
	);
	LUT3 #(
		.INIT('h70)
	) name4540 (
		_w2023_,
		_w2055_,
		_w2617_,
		_w4574_
	);
	LUT3 #(
		.INIT('h01)
	) name4541 (
		_w4573_,
		_w4574_,
		_w4572_,
		_w4575_
	);
	LUT4 #(
		.INIT('h95aa)
	) name4542 (
		\a[29] ,
		_w2550_,
		_w4151_,
		_w4575_,
		_w4576_
	);
	LUT2 #(
		.INIT('h9)
	) name4543 (
		_w4299_,
		_w4301_,
		_w4577_
	);
	LUT2 #(
		.INIT('h4)
	) name4544 (
		_w4576_,
		_w4577_,
		_w4578_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4545 (
		_w1874_,
		_w2076_,
		_w2099_,
		_w2617_,
		_w4579_
	);
	LUT3 #(
		.INIT('h70)
	) name4546 (
		_w2124_,
		_w2133_,
		_w2549_,
		_w4580_
	);
	LUT3 #(
		.INIT('h70)
	) name4547 (
		_w2023_,
		_w2055_,
		_w2854_,
		_w4581_
	);
	LUT3 #(
		.INIT('h01)
	) name4548 (
		_w4579_,
		_w4580_,
		_w4581_,
		_w4582_
	);
	LUT4 #(
		.INIT('h6f00)
	) name4549 (
		_w2299_,
		_w2301_,
		_w2550_,
		_w4582_,
		_w4583_
	);
	LUT4 #(
		.INIT('h45ba)
	) name4550 (
		_w4257_,
		_w4259_,
		_w4263_,
		_w4290_,
		_w4584_
	);
	LUT2 #(
		.INIT('h9)
	) name4551 (
		_w4298_,
		_w4584_,
		_w4585_
	);
	LUT3 #(
		.INIT('h90)
	) name4552 (
		\a[29] ,
		_w4583_,
		_w4585_,
		_w4586_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4553 (
		_w1874_,
		_w2076_,
		_w2099_,
		_w2854_,
		_w4587_
	);
	LUT3 #(
		.INIT('h70)
	) name4554 (
		_w2124_,
		_w2133_,
		_w2617_,
		_w4588_
	);
	LUT3 #(
		.INIT('h70)
	) name4555 (
		_w2155_,
		_w2156_,
		_w2549_,
		_w4589_
	);
	LUT3 #(
		.INIT('h01)
	) name4556 (
		_w4587_,
		_w4588_,
		_w4589_,
		_w4590_
	);
	LUT4 #(
		.INIT('h95aa)
	) name4557 (
		\a[29] ,
		_w2550_,
		_w4209_,
		_w4590_,
		_w4591_
	);
	LUT3 #(
		.INIT('h9a)
	) name4558 (
		_w4257_,
		_w4259_,
		_w4263_,
		_w4592_
	);
	LUT2 #(
		.INIT('h4)
	) name4559 (
		_w4591_,
		_w4592_,
		_w4593_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4560 (
		_w2193_,
		_w2183_,
		_w2213_,
		_w2549_,
		_w4594_
	);
	LUT3 #(
		.INIT('h70)
	) name4561 (
		_w2155_,
		_w2156_,
		_w2617_,
		_w4595_
	);
	LUT3 #(
		.INIT('h70)
	) name4562 (
		_w2124_,
		_w2133_,
		_w2854_,
		_w4596_
	);
	LUT3 #(
		.INIT('h01)
	) name4563 (
		_w4594_,
		_w4595_,
		_w4596_,
		_w4597_
	);
	LUT4 #(
		.INIT('h6f00)
	) name4564 (
		_w2295_,
		_w2297_,
		_w2550_,
		_w4597_,
		_w4598_
	);
	LUT4 #(
		.INIT('h8777)
	) name4565 (
		_w2228_,
		_w2262_,
		_w2273_,
		_w2293_,
		_w4599_
	);
	LUT3 #(
		.INIT('h70)
	) name4566 (
		_w2228_,
		_w2262_,
		_w2407_,
		_w4600_
	);
	LUT3 #(
		.INIT('h70)
	) name4567 (
		_w2273_,
		_w2293_,
		_w2527_,
		_w4601_
	);
	LUT4 #(
		.INIT('h000d)
	) name4568 (
		_w377_,
		_w4599_,
		_w4600_,
		_w4601_,
		_w4602_
	);
	LUT3 #(
		.INIT('h09)
	) name4569 (
		\a[29] ,
		_w4598_,
		_w4602_,
		_w4603_
	);
	LUT3 #(
		.INIT('h15)
	) name4570 (
		_w375_,
		_w2228_,
		_w2262_,
		_w4604_
	);
	LUT3 #(
		.INIT('h70)
	) name4571 (
		_w2228_,
		_w2262_,
		_w2617_,
		_w4605_
	);
	LUT3 #(
		.INIT('h70)
	) name4572 (
		_w2273_,
		_w2293_,
		_w2854_,
		_w4606_
	);
	LUT4 #(
		.INIT('h000d)
	) name4573 (
		_w2550_,
		_w4599_,
		_w4605_,
		_w4606_,
		_w4607_
	);
	LUT3 #(
		.INIT('h07)
	) name4574 (
		_w2228_,
		_w2262_,
		_w2548_,
		_w4608_
	);
	LUT4 #(
		.INIT('haa80)
	) name4575 (
		\a[29] ,
		_w2228_,
		_w2262_,
		_w2548_,
		_w4609_
	);
	LUT3 #(
		.INIT('h84)
	) name4576 (
		_w2214_,
		_w2550_,
		_w4258_,
		_w4610_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4577 (
		_w2193_,
		_w2183_,
		_w2213_,
		_w2854_,
		_w4611_
	);
	LUT3 #(
		.INIT('h70)
	) name4578 (
		_w2228_,
		_w2262_,
		_w2549_,
		_w4612_
	);
	LUT3 #(
		.INIT('h70)
	) name4579 (
		_w2273_,
		_w2293_,
		_w2617_,
		_w4613_
	);
	LUT3 #(
		.INIT('h01)
	) name4580 (
		_w4612_,
		_w4613_,
		_w4611_,
		_w4614_
	);
	LUT2 #(
		.INIT('h4)
	) name4581 (
		_w4610_,
		_w4614_,
		_w4615_
	);
	LUT4 #(
		.INIT('h0800)
	) name4582 (
		_w4607_,
		_w4609_,
		_w4610_,
		_w4614_,
		_w4616_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4583 (
		_w2193_,
		_w2183_,
		_w2213_,
		_w2617_,
		_w4617_
	);
	LUT3 #(
		.INIT('h70)
	) name4584 (
		_w2155_,
		_w2156_,
		_w2854_,
		_w4618_
	);
	LUT3 #(
		.INIT('h70)
	) name4585 (
		_w2273_,
		_w2293_,
		_w2549_,
		_w4619_
	);
	LUT3 #(
		.INIT('h01)
	) name4586 (
		_w4617_,
		_w4618_,
		_w4619_,
		_w4620_
	);
	LUT4 #(
		.INIT('h95aa)
	) name4587 (
		\a[29] ,
		_w2550_,
		_w4293_,
		_w4620_,
		_w4621_
	);
	LUT3 #(
		.INIT('h71)
	) name4588 (
		_w4604_,
		_w4616_,
		_w4621_,
		_w4622_
	);
	LUT3 #(
		.INIT('h60)
	) name4589 (
		\a[29] ,
		_w4598_,
		_w4602_,
		_w4623_
	);
	LUT3 #(
		.INIT('h96)
	) name4590 (
		\a[29] ,
		_w4598_,
		_w4602_,
		_w4624_
	);
	LUT3 #(
		.INIT('h54)
	) name4591 (
		_w4603_,
		_w4622_,
		_w4623_,
		_w4625_
	);
	LUT2 #(
		.INIT('h2)
	) name4592 (
		_w4591_,
		_w4592_,
		_w4626_
	);
	LUT2 #(
		.INIT('h9)
	) name4593 (
		_w4591_,
		_w4592_,
		_w4627_
	);
	LUT3 #(
		.INIT('h69)
	) name4594 (
		\a[29] ,
		_w4583_,
		_w4585_,
		_w4628_
	);
	LUT4 #(
		.INIT('h4d00)
	) name4595 (
		_w4591_,
		_w4592_,
		_w4625_,
		_w4628_,
		_w4629_
	);
	LUT2 #(
		.INIT('h2)
	) name4596 (
		_w4576_,
		_w4577_,
		_w4630_
	);
	LUT2 #(
		.INIT('h9)
	) name4597 (
		_w4576_,
		_w4577_,
		_w4631_
	);
	LUT4 #(
		.INIT('h5501)
	) name4598 (
		_w4578_,
		_w4586_,
		_w4629_,
		_w4630_,
		_w4632_
	);
	LUT3 #(
		.INIT('h06)
	) name4599 (
		\a[29] ,
		_w4568_,
		_w4570_,
		_w4633_
	);
	LUT3 #(
		.INIT('h69)
	) name4600 (
		\a[29] ,
		_w4568_,
		_w4570_,
		_w4634_
	);
	LUT2 #(
		.INIT('h9)
	) name4601 (
		_w4561_,
		_w4562_,
		_w4635_
	);
	LUT4 #(
		.INIT('h4d00)
	) name4602 (
		_w4569_,
		_w4570_,
		_w4632_,
		_w4635_,
		_w4636_
	);
	LUT4 #(
		.INIT('h6996)
	) name4603 (
		\a[29] ,
		_w4306_,
		_w4308_,
		_w4555_,
		_w4637_
	);
	LUT4 #(
		.INIT('h0155)
	) name4604 (
		_w4556_,
		_w4563_,
		_w4636_,
		_w4637_,
		_w4638_
	);
	LUT2 #(
		.INIT('h9)
	) name4605 (
		_w4313_,
		_w4318_,
		_w4639_
	);
	LUT3 #(
		.INIT('h70)
	) name4606 (
		_w1692_,
		_w1723_,
		_w2986_,
		_w4640_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4607 (
		_w1751_,
		_w1742_,
		_w1771_,
		_w2975_,
		_w4641_
	);
	LUT3 #(
		.INIT('h70)
	) name4608 (
		_w1795_,
		_w1796_,
		_w2874_,
		_w4642_
	);
	LUT3 #(
		.INIT('h01)
	) name4609 (
		_w4641_,
		_w4642_,
		_w4640_,
		_w4643_
	);
	LUT4 #(
		.INIT('h6f00)
	) name4610 (
		_w2315_,
		_w2317_,
		_w2875_,
		_w4643_,
		_w4644_
	);
	LUT2 #(
		.INIT('h6)
	) name4611 (
		\a[26] ,
		_w4644_,
		_w4645_
	);
	LUT3 #(
		.INIT('hb2)
	) name4612 (
		_w4638_,
		_w4639_,
		_w4645_,
		_w4646_
	);
	LUT2 #(
		.INIT('h9)
	) name4613 (
		_w4484_,
		_w4485_,
		_w4647_
	);
	LUT2 #(
		.INIT('h9)
	) name4614 (
		_w4492_,
		_w4647_,
		_w4648_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4615 (
		_w1454_,
		_w1426_,
		_w1478_,
		_w3262_,
		_w4649_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name4616 (
		_w3214_,
		_w1584_,
		_w1569_,
		_w1606_,
		_w4650_
	);
	LUT3 #(
		.INIT('h70)
	) name4617 (
		_w1501_,
		_w1545_,
		_w3249_,
		_w4651_
	);
	LUT3 #(
		.INIT('h01)
	) name4618 (
		_w4650_,
		_w4651_,
		_w4649_,
		_w4652_
	);
	LUT4 #(
		.INIT('h6f00)
	) name4619 (
		_w2323_,
		_w2325_,
		_w37_,
		_w4652_,
		_w4653_
	);
	LUT4 #(
		.INIT('h4d8e)
	) name4620 (
		\a[23] ,
		_w4646_,
		_w4648_,
		_w4653_,
		_w4654_
	);
	LUT3 #(
		.INIT('h09)
	) name4621 (
		_w4500_,
		_w4550_,
		_w4654_,
		_w4655_
	);
	LUT3 #(
		.INIT('h60)
	) name4622 (
		_w4500_,
		_w4550_,
		_w4654_,
		_w4656_
	);
	LUT3 #(
		.INIT('h70)
	) name4623 (
		_w1202_,
		_w1233_,
		_w3654_,
		_w4657_
	);
	LUT3 #(
		.INIT('h70)
	) name4624 (
		_w1325_,
		_w1367_,
		_w3311_,
		_w4658_
	);
	LUT3 #(
		.INIT('h70)
	) name4625 (
		_w1253_,
		_w1294_,
		_w3645_,
		_w4659_
	);
	LUT3 #(
		.INIT('h01)
	) name4626 (
		_w4658_,
		_w4659_,
		_w4657_,
		_w4660_
	);
	LUT4 #(
		.INIT('h6f00)
	) name4627 (
		_w2331_,
		_w2333_,
		_w3312_,
		_w4660_,
		_w4661_
	);
	LUT4 #(
		.INIT('h3132)
	) name4628 (
		\a[20] ,
		_w4655_,
		_w4656_,
		_w4661_,
		_w4662_
	);
	LUT3 #(
		.INIT('hd4)
	) name4629 (
		_w4544_,
		_w4549_,
		_w4662_,
		_w4663_
	);
	LUT4 #(
		.INIT('h9669)
	) name4630 (
		\a[20] ,
		_w4502_,
		_w4504_,
		_w4509_,
		_w4664_
	);
	LUT2 #(
		.INIT('h4)
	) name4631 (
		_w4663_,
		_w4664_,
		_w4665_
	);
	LUT2 #(
		.INIT('h2)
	) name4632 (
		_w4663_,
		_w4664_,
		_w4666_
	);
	LUT3 #(
		.INIT('h70)
	) name4633 (
		_w1009_,
		_w1050_,
		_w3709_,
		_w4667_
	);
	LUT3 #(
		.INIT('h70)
	) name4634 (
		_w871_,
		_w927_,
		_w3886_,
		_w4668_
	);
	LUT3 #(
		.INIT('h70)
	) name4635 (
		_w763_,
		_w983_,
		_w3877_,
		_w4669_
	);
	LUT3 #(
		.INIT('h01)
	) name4636 (
		_w4668_,
		_w4669_,
		_w4667_,
		_w4670_
	);
	LUT4 #(
		.INIT('h95aa)
	) name4637 (
		\a[17] ,
		_w2839_,
		_w3710_,
		_w4670_,
		_w4671_
	);
	LUT3 #(
		.INIT('h54)
	) name4638 (
		_w4665_,
		_w4666_,
		_w4671_,
		_w4672_
	);
	LUT2 #(
		.INIT('h2)
	) name4639 (
		_w4543_,
		_w4672_,
		_w4673_
	);
	LUT2 #(
		.INIT('h4)
	) name4640 (
		_w4543_,
		_w4672_,
		_w4674_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4641 (
		_w587_,
		_w608_,
		_w624_,
		_w4382_,
		_w4675_
	);
	LUT3 #(
		.INIT('h70)
	) name4642 (
		_w725_,
		_w764_,
		_w4033_,
		_w4676_
	);
	LUT3 #(
		.INIT('h70)
	) name4643 (
		_w666_,
		_w694_,
		_w4367_,
		_w4677_
	);
	LUT3 #(
		.INIT('h01)
	) name4644 (
		_w4676_,
		_w4677_,
		_w4675_,
		_w4678_
	);
	LUT4 #(
		.INIT('h95aa)
	) name4645 (
		\a[14] ,
		_w2598_,
		_w4034_,
		_w4678_,
		_w4679_
	);
	LUT3 #(
		.INIT('h54)
	) name4646 (
		_w4673_,
		_w4674_,
		_w4679_,
		_w4680_
	);
	LUT3 #(
		.INIT('h54)
	) name4647 (
		_w4539_,
		_w4540_,
		_w4680_,
		_w4681_
	);
	LUT4 #(
		.INIT('hf400)
	) name4648 (
		_w374_,
		_w2361_,
		_w2404_,
		_w4459_,
		_w4682_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4649 (
		_w121_,
		_w418_,
		_w422_,
		_w4458_,
		_w4683_
	);
	LUT3 #(
		.INIT('h18)
	) name4650 (
		\a[8] ,
		\a[9] ,
		\a[10] ,
		_w4684_
	);
	LUT3 #(
		.INIT('h70)
	) name4651 (
		_w352_,
		_w373_,
		_w4684_,
		_w4685_
	);
	LUT2 #(
		.INIT('h1)
	) name4652 (
		_w4683_,
		_w4685_,
		_w4686_
	);
	LUT3 #(
		.INIT('h9a)
	) name4653 (
		\a[11] ,
		_w4682_,
		_w4686_,
		_w4687_
	);
	LUT4 #(
		.INIT('h1211)
	) name4654 (
		\a[11] ,
		_w4681_,
		_w4682_,
		_w4686_,
		_w4688_
	);
	LUT4 #(
		.INIT('h8488)
	) name4655 (
		\a[11] ,
		_w4681_,
		_w4682_,
		_w4686_,
		_w4689_
	);
	LUT4 #(
		.INIT('h6966)
	) name4656 (
		\a[11] ,
		_w4681_,
		_w4682_,
		_w4686_,
		_w4690_
	);
	LUT2 #(
		.INIT('h6)
	) name4657 (
		_w4519_,
		_w4520_,
		_w4691_
	);
	LUT2 #(
		.INIT('h9)
	) name4658 (
		_w4527_,
		_w4691_,
		_w4692_
	);
	LUT3 #(
		.INIT('h45)
	) name4659 (
		_w4688_,
		_w4689_,
		_w4692_,
		_w4693_
	);
	LUT4 #(
		.INIT('h9669)
	) name4660 (
		\a[11] ,
		_w4460_,
		_w4528_,
		_w4530_,
		_w4694_
	);
	LUT4 #(
		.INIT('h7100)
	) name4661 (
		_w4681_,
		_w4687_,
		_w4692_,
		_w4694_,
		_w4695_
	);
	LUT4 #(
		.INIT('h45ba)
	) name4662 (
		_w4688_,
		_w4689_,
		_w4692_,
		_w4694_,
		_w4696_
	);
	LUT2 #(
		.INIT('h6)
	) name4663 (
		_w4690_,
		_w4692_,
		_w4697_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4664 (
		_w486_,
		_w487_,
		_w509_,
		_w4458_,
		_w4698_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4665 (
		_w121_,
		_w418_,
		_w422_,
		_w4684_,
		_w4699_
	);
	LUT4 #(
		.INIT('h6006)
	) name4666 (
		\a[8] ,
		\a[9] ,
		\a[10] ,
		\a[11] ,
		_w4700_
	);
	LUT3 #(
		.INIT('h70)
	) name4667 (
		_w352_,
		_w373_,
		_w4700_,
		_w4701_
	);
	LUT3 #(
		.INIT('h01)
	) name4668 (
		_w4698_,
		_w4699_,
		_w4701_,
		_w4702_
	);
	LUT4 #(
		.INIT('h95aa)
	) name4669 (
		\a[11] ,
		_w2535_,
		_w4459_,
		_w4702_,
		_w4703_
	);
	LUT2 #(
		.INIT('h9)
	) name4670 (
		_w4543_,
		_w4672_,
		_w4704_
	);
	LUT3 #(
		.INIT('h70)
	) name4671 (
		_w1071_,
		_w1102_,
		_w3709_,
		_w4705_
	);
	LUT3 #(
		.INIT('h70)
	) name4672 (
		_w763_,
		_w983_,
		_w3886_,
		_w4706_
	);
	LUT3 #(
		.INIT('h70)
	) name4673 (
		_w1009_,
		_w1050_,
		_w3877_,
		_w4707_
	);
	LUT3 #(
		.INIT('h01)
	) name4674 (
		_w4706_,
		_w4707_,
		_w4705_,
		_w4708_
	);
	LUT4 #(
		.INIT('h6f00)
	) name4675 (
		_w2339_,
		_w2341_,
		_w3710_,
		_w4708_,
		_w4709_
	);
	LUT3 #(
		.INIT('h96)
	) name4676 (
		_w4544_,
		_w4549_,
		_w4662_,
		_w4710_
	);
	LUT3 #(
		.INIT('h90)
	) name4677 (
		\a[17] ,
		_w4709_,
		_w4710_,
		_w4711_
	);
	LUT3 #(
		.INIT('h06)
	) name4678 (
		\a[17] ,
		_w4709_,
		_w4710_,
		_w4712_
	);
	LUT3 #(
		.INIT('h69)
	) name4679 (
		\a[17] ,
		_w4709_,
		_w4710_,
		_w4713_
	);
	LUT3 #(
		.INIT('h96)
	) name4680 (
		_w4500_,
		_w4550_,
		_w4654_,
		_w4714_
	);
	LUT3 #(
		.INIT('h69)
	) name4681 (
		\a[20] ,
		_w4661_,
		_w4714_,
		_w4715_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4682 (
		_w1751_,
		_w1742_,
		_w1771_,
		_w2986_,
		_w4716_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4683 (
		_w1817_,
		_w1799_,
		_w1840_,
		_w2874_,
		_w4717_
	);
	LUT3 #(
		.INIT('h70)
	) name4684 (
		_w1795_,
		_w1796_,
		_w2975_,
		_w4718_
	);
	LUT3 #(
		.INIT('h01)
	) name4685 (
		_w4717_,
		_w4718_,
		_w4716_,
		_w4719_
	);
	LUT4 #(
		.INIT('h95aa)
	) name4686 (
		\a[26] ,
		_w2875_,
		_w3909_,
		_w4719_,
		_w4720_
	);
	LUT4 #(
		.INIT('h001e)
	) name4687 (
		_w4563_,
		_w4636_,
		_w4637_,
		_w4720_,
		_w4721_
	);
	LUT4 #(
		.INIT('h54ab)
	) name4688 (
		_w4571_,
		_w4632_,
		_w4633_,
		_w4635_,
		_w4722_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4689 (
		_w1817_,
		_w1799_,
		_w1840_,
		_w2975_,
		_w4723_
	);
	LUT3 #(
		.INIT('h70)
	) name4690 (
		_w1795_,
		_w1796_,
		_w2986_,
		_w4724_
	);
	LUT3 #(
		.INIT('h70)
	) name4691 (
		_w1863_,
		_w1875_,
		_w2874_,
		_w4725_
	);
	LUT3 #(
		.INIT('h01)
	) name4692 (
		_w4724_,
		_w4725_,
		_w4723_,
		_w4726_
	);
	LUT4 #(
		.INIT('h6f00)
	) name4693 (
		_w2311_,
		_w2313_,
		_w2875_,
		_w4726_,
		_w4727_
	);
	LUT2 #(
		.INIT('h6)
	) name4694 (
		\a[26] ,
		_w4727_,
		_w4728_
	);
	LUT2 #(
		.INIT('h2)
	) name4695 (
		_w4722_,
		_w4728_,
		_w4729_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4696 (
		_w1817_,
		_w1799_,
		_w1840_,
		_w2986_,
		_w4730_
	);
	LUT3 #(
		.INIT('h70)
	) name4697 (
		_w1898_,
		_w1928_,
		_w2874_,
		_w4731_
	);
	LUT3 #(
		.INIT('h70)
	) name4698 (
		_w1863_,
		_w1875_,
		_w2975_,
		_w4732_
	);
	LUT3 #(
		.INIT('h01)
	) name4699 (
		_w4731_,
		_w4732_,
		_w4730_,
		_w4733_
	);
	LUT4 #(
		.INIT('h95aa)
	) name4700 (
		\a[26] ,
		_w2875_,
		_w3972_,
		_w4733_,
		_w4734_
	);
	LUT3 #(
		.INIT('h09)
	) name4701 (
		_w4632_,
		_w4634_,
		_w4734_,
		_w4735_
	);
	LUT3 #(
		.INIT('h1e)
	) name4702 (
		_w4586_,
		_w4629_,
		_w4631_,
		_w4736_
	);
	LUT3 #(
		.INIT('h70)
	) name4703 (
		_w1501_,
		_w1949_,
		_w2874_,
		_w4737_
	);
	LUT3 #(
		.INIT('h70)
	) name4704 (
		_w1898_,
		_w1928_,
		_w2975_,
		_w4738_
	);
	LUT3 #(
		.INIT('h70)
	) name4705 (
		_w1863_,
		_w1875_,
		_w2986_,
		_w4739_
	);
	LUT3 #(
		.INIT('h01)
	) name4706 (
		_w4738_,
		_w4739_,
		_w4737_,
		_w4740_
	);
	LUT4 #(
		.INIT('h6f00)
	) name4707 (
		_w2307_,
		_w2309_,
		_w2875_,
		_w4740_,
		_w4741_
	);
	LUT2 #(
		.INIT('h6)
	) name4708 (
		\a[26] ,
		_w4741_,
		_w4742_
	);
	LUT2 #(
		.INIT('h2)
	) name4709 (
		_w4736_,
		_w4742_,
		_w4743_
	);
	LUT4 #(
		.INIT('h54ab)
	) name4710 (
		_w4593_,
		_w4625_,
		_w4626_,
		_w4628_,
		_w4744_
	);
	LUT3 #(
		.INIT('h70)
	) name4711 (
		_w1973_,
		_w1997_,
		_w2874_,
		_w4745_
	);
	LUT3 #(
		.INIT('h70)
	) name4712 (
		_w1898_,
		_w1928_,
		_w2986_,
		_w4746_
	);
	LUT3 #(
		.INIT('h70)
	) name4713 (
		_w1501_,
		_w1949_,
		_w2975_,
		_w4747_
	);
	LUT3 #(
		.INIT('h01)
	) name4714 (
		_w4746_,
		_w4747_,
		_w4745_,
		_w4748_
	);
	LUT4 #(
		.INIT('h95aa)
	) name4715 (
		\a[26] ,
		_w2875_,
		_w4126_,
		_w4748_,
		_w4749_
	);
	LUT2 #(
		.INIT('h2)
	) name4716 (
		_w4744_,
		_w4749_,
		_w4750_
	);
	LUT2 #(
		.INIT('h9)
	) name4717 (
		_w4625_,
		_w4627_,
		_w4751_
	);
	LUT3 #(
		.INIT('h70)
	) name4718 (
		_w1973_,
		_w1997_,
		_w2975_,
		_w4752_
	);
	LUT3 #(
		.INIT('h70)
	) name4719 (
		_w1501_,
		_w1949_,
		_w2986_,
		_w4753_
	);
	LUT3 #(
		.INIT('h70)
	) name4720 (
		_w2023_,
		_w2055_,
		_w2874_,
		_w4754_
	);
	LUT3 #(
		.INIT('h01)
	) name4721 (
		_w4753_,
		_w4754_,
		_w4752_,
		_w4755_
	);
	LUT4 #(
		.INIT('h6f00)
	) name4722 (
		_w2303_,
		_w2305_,
		_w2875_,
		_w4755_,
		_w4756_
	);
	LUT2 #(
		.INIT('h6)
	) name4723 (
		\a[26] ,
		_w4756_,
		_w4757_
	);
	LUT4 #(
		.INIT('h8241)
	) name4724 (
		\a[26] ,
		_w4625_,
		_w4627_,
		_w4756_,
		_w4758_
	);
	LUT3 #(
		.INIT('h70)
	) name4725 (
		_w1973_,
		_w1997_,
		_w2986_,
		_w4759_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4726 (
		_w1874_,
		_w2076_,
		_w2099_,
		_w2874_,
		_w4760_
	);
	LUT3 #(
		.INIT('h70)
	) name4727 (
		_w2023_,
		_w2055_,
		_w2975_,
		_w4761_
	);
	LUT3 #(
		.INIT('h01)
	) name4728 (
		_w4760_,
		_w4761_,
		_w4759_,
		_w4762_
	);
	LUT4 #(
		.INIT('h95aa)
	) name4729 (
		\a[26] ,
		_w2875_,
		_w4151_,
		_w4762_,
		_w4763_
	);
	LUT2 #(
		.INIT('h9)
	) name4730 (
		_w4622_,
		_w4624_,
		_w4764_
	);
	LUT2 #(
		.INIT('h4)
	) name4731 (
		_w4763_,
		_w4764_,
		_w4765_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4732 (
		_w1874_,
		_w2076_,
		_w2099_,
		_w2975_,
		_w4766_
	);
	LUT3 #(
		.INIT('h70)
	) name4733 (
		_w2124_,
		_w2133_,
		_w2874_,
		_w4767_
	);
	LUT3 #(
		.INIT('h70)
	) name4734 (
		_w2023_,
		_w2055_,
		_w2986_,
		_w4768_
	);
	LUT3 #(
		.INIT('h01)
	) name4735 (
		_w4766_,
		_w4767_,
		_w4768_,
		_w4769_
	);
	LUT4 #(
		.INIT('h6f00)
	) name4736 (
		_w2299_,
		_w2301_,
		_w2875_,
		_w4769_,
		_w4770_
	);
	LUT3 #(
		.INIT('h69)
	) name4737 (
		_w4604_,
		_w4616_,
		_w4621_,
		_w4771_
	);
	LUT3 #(
		.INIT('h90)
	) name4738 (
		\a[26] ,
		_w4770_,
		_w4771_,
		_w4772_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4739 (
		_w1874_,
		_w2076_,
		_w2099_,
		_w2986_,
		_w4773_
	);
	LUT3 #(
		.INIT('h70)
	) name4740 (
		_w2124_,
		_w2133_,
		_w2975_,
		_w4774_
	);
	LUT3 #(
		.INIT('h70)
	) name4741 (
		_w2155_,
		_w2156_,
		_w2874_,
		_w4775_
	);
	LUT3 #(
		.INIT('h01)
	) name4742 (
		_w4773_,
		_w4774_,
		_w4775_,
		_w4776_
	);
	LUT4 #(
		.INIT('h95aa)
	) name4743 (
		\a[26] ,
		_w2875_,
		_w4209_,
		_w4776_,
		_w4777_
	);
	LUT3 #(
		.INIT('h8a)
	) name4744 (
		\a[29] ,
		_w4608_,
		_w4607_,
		_w4778_
	);
	LUT2 #(
		.INIT('h9)
	) name4745 (
		_w4615_,
		_w4778_,
		_w4779_
	);
	LUT2 #(
		.INIT('h4)
	) name4746 (
		_w4777_,
		_w4779_,
		_w4780_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4747 (
		_w2193_,
		_w2183_,
		_w2213_,
		_w2874_,
		_w4781_
	);
	LUT3 #(
		.INIT('h70)
	) name4748 (
		_w2155_,
		_w2156_,
		_w2975_,
		_w4782_
	);
	LUT3 #(
		.INIT('h70)
	) name4749 (
		_w2124_,
		_w2133_,
		_w2986_,
		_w4783_
	);
	LUT3 #(
		.INIT('h01)
	) name4750 (
		_w4781_,
		_w4782_,
		_w4783_,
		_w4784_
	);
	LUT4 #(
		.INIT('h6f00)
	) name4751 (
		_w2295_,
		_w2297_,
		_w2875_,
		_w4784_,
		_w4785_
	);
	LUT4 #(
		.INIT('h002a)
	) name4752 (
		\a[29] ,
		_w2228_,
		_w2262_,
		_w2548_,
		_w4786_
	);
	LUT2 #(
		.INIT('h9)
	) name4753 (
		_w4607_,
		_w4786_,
		_w4787_
	);
	LUT3 #(
		.INIT('h90)
	) name4754 (
		\a[26] ,
		_w4785_,
		_w4787_,
		_w4788_
	);
	LUT3 #(
		.INIT('h70)
	) name4755 (
		_w2228_,
		_w2262_,
		_w2975_,
		_w4789_
	);
	LUT3 #(
		.INIT('h70)
	) name4756 (
		_w2273_,
		_w2293_,
		_w2986_,
		_w4790_
	);
	LUT4 #(
		.INIT('h000d)
	) name4757 (
		_w2875_,
		_w4599_,
		_w4789_,
		_w4790_,
		_w4791_
	);
	LUT3 #(
		.INIT('h07)
	) name4758 (
		_w2228_,
		_w2262_,
		_w2873_,
		_w4792_
	);
	LUT4 #(
		.INIT('haa80)
	) name4759 (
		\a[26] ,
		_w2228_,
		_w2262_,
		_w2873_,
		_w4793_
	);
	LUT3 #(
		.INIT('h84)
	) name4760 (
		_w2214_,
		_w2875_,
		_w4258_,
		_w4794_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4761 (
		_w2193_,
		_w2183_,
		_w2213_,
		_w2986_,
		_w4795_
	);
	LUT3 #(
		.INIT('h70)
	) name4762 (
		_w2228_,
		_w2262_,
		_w2874_,
		_w4796_
	);
	LUT3 #(
		.INIT('h70)
	) name4763 (
		_w2273_,
		_w2293_,
		_w2975_,
		_w4797_
	);
	LUT3 #(
		.INIT('h01)
	) name4764 (
		_w4796_,
		_w4797_,
		_w4795_,
		_w4798_
	);
	LUT2 #(
		.INIT('h4)
	) name4765 (
		_w4794_,
		_w4798_,
		_w4799_
	);
	LUT4 #(
		.INIT('h0800)
	) name4766 (
		_w4791_,
		_w4793_,
		_w4794_,
		_w4798_,
		_w4800_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4767 (
		_w2193_,
		_w2183_,
		_w2213_,
		_w2975_,
		_w4801_
	);
	LUT3 #(
		.INIT('h70)
	) name4768 (
		_w2155_,
		_w2156_,
		_w2986_,
		_w4802_
	);
	LUT3 #(
		.INIT('h70)
	) name4769 (
		_w2273_,
		_w2293_,
		_w2874_,
		_w4803_
	);
	LUT3 #(
		.INIT('h01)
	) name4770 (
		_w4801_,
		_w4802_,
		_w4803_,
		_w4804_
	);
	LUT4 #(
		.INIT('h95aa)
	) name4771 (
		\a[26] ,
		_w2875_,
		_w4293_,
		_w4804_,
		_w4805_
	);
	LUT3 #(
		.INIT('h71)
	) name4772 (
		_w4608_,
		_w4800_,
		_w4805_,
		_w4806_
	);
	LUT3 #(
		.INIT('h06)
	) name4773 (
		\a[26] ,
		_w4785_,
		_w4787_,
		_w4807_
	);
	LUT3 #(
		.INIT('h69)
	) name4774 (
		\a[26] ,
		_w4785_,
		_w4787_,
		_w4808_
	);
	LUT3 #(
		.INIT('h54)
	) name4775 (
		_w4788_,
		_w4806_,
		_w4807_,
		_w4809_
	);
	LUT2 #(
		.INIT('h2)
	) name4776 (
		_w4777_,
		_w4779_,
		_w4810_
	);
	LUT2 #(
		.INIT('h9)
	) name4777 (
		_w4777_,
		_w4779_,
		_w4811_
	);
	LUT3 #(
		.INIT('h69)
	) name4778 (
		\a[26] ,
		_w4770_,
		_w4771_,
		_w4812_
	);
	LUT4 #(
		.INIT('h4d00)
	) name4779 (
		_w4777_,
		_w4779_,
		_w4809_,
		_w4812_,
		_w4813_
	);
	LUT2 #(
		.INIT('h2)
	) name4780 (
		_w4763_,
		_w4764_,
		_w4814_
	);
	LUT2 #(
		.INIT('h9)
	) name4781 (
		_w4763_,
		_w4764_,
		_w4815_
	);
	LUT4 #(
		.INIT('h5501)
	) name4782 (
		_w4765_,
		_w4772_,
		_w4813_,
		_w4814_,
		_w4816_
	);
	LUT4 #(
		.INIT('h1428)
	) name4783 (
		\a[26] ,
		_w4625_,
		_w4627_,
		_w4756_,
		_w4817_
	);
	LUT4 #(
		.INIT('h6996)
	) name4784 (
		\a[26] ,
		_w4625_,
		_w4627_,
		_w4756_,
		_w4818_
	);
	LUT2 #(
		.INIT('h9)
	) name4785 (
		_w4744_,
		_w4749_,
		_w4819_
	);
	LUT4 #(
		.INIT('h2b00)
	) name4786 (
		_w4751_,
		_w4757_,
		_w4816_,
		_w4819_,
		_w4820_
	);
	LUT2 #(
		.INIT('h4)
	) name4787 (
		_w4736_,
		_w4742_,
		_w4821_
	);
	LUT2 #(
		.INIT('h9)
	) name4788 (
		_w4736_,
		_w4742_,
		_w4822_
	);
	LUT4 #(
		.INIT('h5501)
	) name4789 (
		_w4743_,
		_w4750_,
		_w4820_,
		_w4821_,
		_w4823_
	);
	LUT3 #(
		.INIT('h60)
	) name4790 (
		_w4632_,
		_w4634_,
		_w4734_,
		_w4824_
	);
	LUT3 #(
		.INIT('h96)
	) name4791 (
		_w4632_,
		_w4634_,
		_w4734_,
		_w4825_
	);
	LUT2 #(
		.INIT('h9)
	) name4792 (
		_w4722_,
		_w4728_,
		_w4826_
	);
	LUT4 #(
		.INIT('hba00)
	) name4793 (
		_w4735_,
		_w4823_,
		_w4825_,
		_w4826_,
		_w4827_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name4794 (
		_w4563_,
		_w4636_,
		_w4637_,
		_w4720_,
		_w4828_
	);
	LUT4 #(
		.INIT('h0155)
	) name4795 (
		_w4721_,
		_w4729_,
		_w4827_,
		_w4828_,
		_w4829_
	);
	LUT3 #(
		.INIT('h96)
	) name4796 (
		_w4638_,
		_w4639_,
		_w4645_,
		_w4830_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4797 (
		_w1584_,
		_w1569_,
		_w1606_,
		_w3249_,
		_w4831_
	);
	LUT3 #(
		.INIT('h70)
	) name4798 (
		_w1501_,
		_w1545_,
		_w3262_,
		_w4832_
	);
	LUT3 #(
		.INIT('h2a)
	) name4799 (
		_w3214_,
		_w1620_,
		_w1661_,
		_w4833_
	);
	LUT3 #(
		.INIT('h01)
	) name4800 (
		_w4831_,
		_w4832_,
		_w4833_,
		_w4834_
	);
	LUT4 #(
		.INIT('h95aa)
	) name4801 (
		\a[23] ,
		_w37_,
		_w3495_,
		_w4834_,
		_w4835_
	);
	LUT4 #(
		.INIT('h9669)
	) name4802 (
		\a[23] ,
		_w4646_,
		_w4648_,
		_w4653_,
		_w4836_
	);
	LUT4 #(
		.INIT('h004d)
	) name4803 (
		_w4829_,
		_w4830_,
		_w4835_,
		_w4836_,
		_w4837_
	);
	LUT4 #(
		.INIT('hb200)
	) name4804 (
		_w4829_,
		_w4830_,
		_w4835_,
		_w4836_,
		_w4838_
	);
	LUT3 #(
		.INIT('h70)
	) name4805 (
		_w1381_,
		_w1398_,
		_w3311_,
		_w4839_
	);
	LUT3 #(
		.INIT('h70)
	) name4806 (
		_w1325_,
		_w1367_,
		_w3645_,
		_w4840_
	);
	LUT3 #(
		.INIT('h70)
	) name4807 (
		_w1253_,
		_w1294_,
		_w3654_,
		_w4841_
	);
	LUT3 #(
		.INIT('h01)
	) name4808 (
		_w4840_,
		_w4841_,
		_w4839_,
		_w4842_
	);
	LUT4 #(
		.INIT('h95aa)
	) name4809 (
		\a[20] ,
		_w3182_,
		_w3312_,
		_w4842_,
		_w4843_
	);
	LUT3 #(
		.INIT('h54)
	) name4810 (
		_w4837_,
		_w4838_,
		_w4843_,
		_w4844_
	);
	LUT2 #(
		.INIT('h2)
	) name4811 (
		_w4715_,
		_w4844_,
		_w4845_
	);
	LUT2 #(
		.INIT('h4)
	) name4812 (
		_w4715_,
		_w4844_,
		_w4846_
	);
	LUT3 #(
		.INIT('h70)
	) name4813 (
		_w1136_,
		_w1187_,
		_w3709_,
		_w4847_
	);
	LUT3 #(
		.INIT('h70)
	) name4814 (
		_w1009_,
		_w1050_,
		_w3886_,
		_w4848_
	);
	LUT3 #(
		.INIT('h70)
	) name4815 (
		_w1071_,
		_w1102_,
		_w3877_,
		_w4849_
	);
	LUT3 #(
		.INIT('h01)
	) name4816 (
		_w4848_,
		_w4849_,
		_w4847_,
		_w4850_
	);
	LUT4 #(
		.INIT('h95aa)
	) name4817 (
		\a[17] ,
		_w2936_,
		_w3710_,
		_w4850_,
		_w4851_
	);
	LUT3 #(
		.INIT('h54)
	) name4818 (
		_w4845_,
		_w4846_,
		_w4851_,
		_w4852_
	);
	LUT3 #(
		.INIT('h54)
	) name4819 (
		_w4711_,
		_w4712_,
		_w4852_,
		_w4853_
	);
	LUT2 #(
		.INIT('h9)
	) name4820 (
		_w4663_,
		_w4664_,
		_w4854_
	);
	LUT2 #(
		.INIT('h6)
	) name4821 (
		_w4671_,
		_w4854_,
		_w4855_
	);
	LUT3 #(
		.INIT('h70)
	) name4822 (
		_w725_,
		_w764_,
		_w4367_,
		_w4856_
	);
	LUT3 #(
		.INIT('h70)
	) name4823 (
		_w801_,
		_w851_,
		_w4033_,
		_w4857_
	);
	LUT3 #(
		.INIT('h70)
	) name4824 (
		_w666_,
		_w694_,
		_w4382_,
		_w4858_
	);
	LUT3 #(
		.INIT('h01)
	) name4825 (
		_w4857_,
		_w4858_,
		_w4856_,
		_w4859_
	);
	LUT4 #(
		.INIT('h6f00)
	) name4826 (
		_w2347_,
		_w2349_,
		_w4034_,
		_w4859_,
		_w4860_
	);
	LUT4 #(
		.INIT('hd4e8)
	) name4827 (
		\a[14] ,
		_w4853_,
		_w4855_,
		_w4860_,
		_w4861_
	);
	LUT3 #(
		.INIT('h09)
	) name4828 (
		_w4679_,
		_w4704_,
		_w4861_,
		_w4862_
	);
	LUT3 #(
		.INIT('h60)
	) name4829 (
		_w4679_,
		_w4704_,
		_w4861_,
		_w4863_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4830 (
		_w486_,
		_w487_,
		_w509_,
		_w4684_,
		_w4864_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4831 (
		_w121_,
		_w418_,
		_w422_,
		_w4700_,
		_w4865_
	);
	LUT3 #(
		.INIT('h70)
	) name4832 (
		_w544_,
		_w558_,
		_w4458_,
		_w4866_
	);
	LUT3 #(
		.INIT('h01)
	) name4833 (
		_w4864_,
		_w4865_,
		_w4866_,
		_w4867_
	);
	LUT4 #(
		.INIT('h6f00)
	) name4834 (
		_w2355_,
		_w2357_,
		_w4459_,
		_w4867_,
		_w4868_
	);
	LUT4 #(
		.INIT('h3132)
	) name4835 (
		\a[11] ,
		_w4862_,
		_w4863_,
		_w4868_,
		_w4869_
	);
	LUT2 #(
		.INIT('h9)
	) name4836 (
		_w4541_,
		_w4680_,
		_w4870_
	);
	LUT3 #(
		.INIT('h8e)
	) name4837 (
		_w4703_,
		_w4869_,
		_w4870_,
		_w4871_
	);
	LUT3 #(
		.INIT('h06)
	) name4838 (
		_w4690_,
		_w4692_,
		_w4871_,
		_w4872_
	);
	LUT3 #(
		.INIT('h96)
	) name4839 (
		_w4703_,
		_w4869_,
		_w4870_,
		_w4873_
	);
	LUT2 #(
		.INIT('h9)
	) name4840 (
		\a[5] ,
		\a[6] ,
		_w4874_
	);
	LUT4 #(
		.INIT('h0180)
	) name4841 (
		\a[5] ,
		\a[6] ,
		\a[7] ,
		\a[8] ,
		_w4875_
	);
	LUT4 #(
		.INIT('h0660)
	) name4842 (
		\a[5] ,
		\a[6] ,
		\a[7] ,
		\a[8] ,
		_w4876_
	);
	LUT4 #(
		.INIT('h5150)
	) name4843 (
		_w374_,
		_w2361_,
		_w4875_,
		_w4876_,
		_w4877_
	);
	LUT2 #(
		.INIT('h9)
	) name4844 (
		_w4713_,
		_w4852_,
		_w4878_
	);
	LUT3 #(
		.INIT('h70)
	) name4845 (
		_w725_,
		_w764_,
		_w4382_,
		_w4879_
	);
	LUT3 #(
		.INIT('h70)
	) name4846 (
		_w801_,
		_w851_,
		_w4367_,
		_w4880_
	);
	LUT3 #(
		.INIT('h70)
	) name4847 (
		_w871_,
		_w927_,
		_w4033_,
		_w4881_
	);
	LUT3 #(
		.INIT('h01)
	) name4848 (
		_w4880_,
		_w4881_,
		_w4879_,
		_w4882_
	);
	LUT4 #(
		.INIT('h95aa)
	) name4849 (
		\a[14] ,
		_w2724_,
		_w4034_,
		_w4882_,
		_w4883_
	);
	LUT2 #(
		.INIT('h9)
	) name4850 (
		_w4715_,
		_w4844_,
		_w4884_
	);
	LUT2 #(
		.INIT('h9)
	) name4851 (
		_w4851_,
		_w4884_,
		_w4885_
	);
	LUT3 #(
		.INIT('h2a)
	) name4852 (
		_w3214_,
		_w1692_,
		_w1723_,
		_w4886_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4853 (
		_w1584_,
		_w1569_,
		_w1606_,
		_w3262_,
		_w4887_
	);
	LUT3 #(
		.INIT('h70)
	) name4854 (
		_w1620_,
		_w1661_,
		_w3249_,
		_w4888_
	);
	LUT3 #(
		.INIT('h01)
	) name4855 (
		_w4887_,
		_w4888_,
		_w4886_,
		_w4889_
	);
	LUT4 #(
		.INIT('h6f00)
	) name4856 (
		_w2319_,
		_w2321_,
		_w37_,
		_w4889_,
		_w4890_
	);
	LUT2 #(
		.INIT('h6)
	) name4857 (
		\a[23] ,
		_w4890_,
		_w4891_
	);
	LUT4 #(
		.INIT('h001e)
	) name4858 (
		_w4729_,
		_w4827_,
		_w4828_,
		_w4891_,
		_w4892_
	);
	LUT3 #(
		.INIT('h70)
	) name4859 (
		_w1692_,
		_w1723_,
		_w3249_,
		_w4893_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name4860 (
		_w3214_,
		_w1751_,
		_w1742_,
		_w1771_,
		_w4894_
	);
	LUT3 #(
		.INIT('h70)
	) name4861 (
		_w1620_,
		_w1661_,
		_w3262_,
		_w4895_
	);
	LUT3 #(
		.INIT('h01)
	) name4862 (
		_w4894_,
		_w4895_,
		_w4893_,
		_w4896_
	);
	LUT4 #(
		.INIT('h95aa)
	) name4863 (
		\a[23] ,
		_w37_,
		_w3599_,
		_w4896_,
		_w4897_
	);
	LUT4 #(
		.INIT('h54ab)
	) name4864 (
		_w4735_,
		_w4823_,
		_w4824_,
		_w4826_,
		_w4898_
	);
	LUT2 #(
		.INIT('h4)
	) name4865 (
		_w4897_,
		_w4898_,
		_w4899_
	);
	LUT3 #(
		.INIT('h70)
	) name4866 (
		_w1692_,
		_w1723_,
		_w3262_,
		_w4900_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4867 (
		_w1751_,
		_w1742_,
		_w1771_,
		_w3249_,
		_w4901_
	);
	LUT3 #(
		.INIT('h2a)
	) name4868 (
		_w3214_,
		_w1795_,
		_w1796_,
		_w4902_
	);
	LUT3 #(
		.INIT('h01)
	) name4869 (
		_w4901_,
		_w4902_,
		_w4900_,
		_w4903_
	);
	LUT4 #(
		.INIT('h6f00)
	) name4870 (
		_w2315_,
		_w2317_,
		_w37_,
		_w4903_,
		_w4904_
	);
	LUT2 #(
		.INIT('h6)
	) name4871 (
		\a[23] ,
		_w4904_,
		_w4905_
	);
	LUT2 #(
		.INIT('h9)
	) name4872 (
		_w4823_,
		_w4825_,
		_w4906_
	);
	LUT3 #(
		.INIT('h09)
	) name4873 (
		_w4823_,
		_w4825_,
		_w4905_,
		_w4907_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4874 (
		_w1751_,
		_w1742_,
		_w1771_,
		_w3262_,
		_w4908_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name4875 (
		_w3214_,
		_w1817_,
		_w1799_,
		_w1840_,
		_w4909_
	);
	LUT3 #(
		.INIT('h70)
	) name4876 (
		_w1795_,
		_w1796_,
		_w3249_,
		_w4910_
	);
	LUT3 #(
		.INIT('h01)
	) name4877 (
		_w4909_,
		_w4910_,
		_w4908_,
		_w4911_
	);
	LUT4 #(
		.INIT('h95aa)
	) name4878 (
		\a[23] ,
		_w37_,
		_w3909_,
		_w4911_,
		_w4912_
	);
	LUT4 #(
		.INIT('h001e)
	) name4879 (
		_w4750_,
		_w4820_,
		_w4822_,
		_w4912_,
		_w4913_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4880 (
		_w1817_,
		_w1799_,
		_w1840_,
		_w3249_,
		_w4914_
	);
	LUT3 #(
		.INIT('h70)
	) name4881 (
		_w1795_,
		_w1796_,
		_w3262_,
		_w4915_
	);
	LUT3 #(
		.INIT('h2a)
	) name4882 (
		_w3214_,
		_w1863_,
		_w1875_,
		_w4916_
	);
	LUT3 #(
		.INIT('h01)
	) name4883 (
		_w4915_,
		_w4916_,
		_w4914_,
		_w4917_
	);
	LUT4 #(
		.INIT('h6f00)
	) name4884 (
		_w2311_,
		_w2313_,
		_w37_,
		_w4917_,
		_w4918_
	);
	LUT2 #(
		.INIT('h6)
	) name4885 (
		\a[23] ,
		_w4918_,
		_w4919_
	);
	LUT4 #(
		.INIT('h54ab)
	) name4886 (
		_w4758_,
		_w4816_,
		_w4817_,
		_w4819_,
		_w4920_
	);
	LUT2 #(
		.INIT('h4)
	) name4887 (
		_w4919_,
		_w4920_,
		_w4921_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4888 (
		_w1817_,
		_w1799_,
		_w1840_,
		_w3262_,
		_w4922_
	);
	LUT3 #(
		.INIT('h2a)
	) name4889 (
		_w3214_,
		_w1898_,
		_w1928_,
		_w4923_
	);
	LUT3 #(
		.INIT('h70)
	) name4890 (
		_w1863_,
		_w1875_,
		_w3249_,
		_w4924_
	);
	LUT3 #(
		.INIT('h01)
	) name4891 (
		_w4923_,
		_w4924_,
		_w4922_,
		_w4925_
	);
	LUT4 #(
		.INIT('h95aa)
	) name4892 (
		\a[23] ,
		_w37_,
		_w3972_,
		_w4925_,
		_w4926_
	);
	LUT3 #(
		.INIT('h09)
	) name4893 (
		_w4816_,
		_w4818_,
		_w4926_,
		_w4927_
	);
	LUT3 #(
		.INIT('h2a)
	) name4894 (
		_w3214_,
		_w1501_,
		_w1949_,
		_w4928_
	);
	LUT3 #(
		.INIT('h70)
	) name4895 (
		_w1898_,
		_w1928_,
		_w3249_,
		_w4929_
	);
	LUT3 #(
		.INIT('h70)
	) name4896 (
		_w1863_,
		_w1875_,
		_w3262_,
		_w4930_
	);
	LUT3 #(
		.INIT('h01)
	) name4897 (
		_w4929_,
		_w4930_,
		_w4928_,
		_w4931_
	);
	LUT4 #(
		.INIT('h6f00)
	) name4898 (
		_w2307_,
		_w2309_,
		_w37_,
		_w4931_,
		_w4932_
	);
	LUT2 #(
		.INIT('h6)
	) name4899 (
		\a[23] ,
		_w4932_,
		_w4933_
	);
	LUT3 #(
		.INIT('h1e)
	) name4900 (
		_w4772_,
		_w4813_,
		_w4815_,
		_w4934_
	);
	LUT2 #(
		.INIT('h4)
	) name4901 (
		_w4933_,
		_w4934_,
		_w4935_
	);
	LUT4 #(
		.INIT('h54ab)
	) name4902 (
		_w4780_,
		_w4809_,
		_w4810_,
		_w4812_,
		_w4936_
	);
	LUT3 #(
		.INIT('h2a)
	) name4903 (
		_w3214_,
		_w1973_,
		_w1997_,
		_w4937_
	);
	LUT3 #(
		.INIT('h70)
	) name4904 (
		_w1898_,
		_w1928_,
		_w3262_,
		_w4938_
	);
	LUT3 #(
		.INIT('h70)
	) name4905 (
		_w1501_,
		_w1949_,
		_w3249_,
		_w4939_
	);
	LUT3 #(
		.INIT('h01)
	) name4906 (
		_w4938_,
		_w4939_,
		_w4937_,
		_w4940_
	);
	LUT4 #(
		.INIT('h95aa)
	) name4907 (
		\a[23] ,
		_w37_,
		_w4126_,
		_w4940_,
		_w4941_
	);
	LUT2 #(
		.INIT('h2)
	) name4908 (
		_w4936_,
		_w4941_,
		_w4942_
	);
	LUT2 #(
		.INIT('h9)
	) name4909 (
		_w4809_,
		_w4811_,
		_w4943_
	);
	LUT3 #(
		.INIT('h70)
	) name4910 (
		_w1973_,
		_w1997_,
		_w3249_,
		_w4944_
	);
	LUT3 #(
		.INIT('h70)
	) name4911 (
		_w1501_,
		_w1949_,
		_w3262_,
		_w4945_
	);
	LUT3 #(
		.INIT('h2a)
	) name4912 (
		_w3214_,
		_w2023_,
		_w2055_,
		_w4946_
	);
	LUT3 #(
		.INIT('h01)
	) name4913 (
		_w4945_,
		_w4946_,
		_w4944_,
		_w4947_
	);
	LUT4 #(
		.INIT('h6f00)
	) name4914 (
		_w2303_,
		_w2305_,
		_w37_,
		_w4947_,
		_w4948_
	);
	LUT2 #(
		.INIT('h6)
	) name4915 (
		\a[23] ,
		_w4948_,
		_w4949_
	);
	LUT4 #(
		.INIT('h8241)
	) name4916 (
		\a[23] ,
		_w4809_,
		_w4811_,
		_w4948_,
		_w4950_
	);
	LUT3 #(
		.INIT('h70)
	) name4917 (
		_w1973_,
		_w1997_,
		_w3262_,
		_w4951_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name4918 (
		_w3214_,
		_w1874_,
		_w2076_,
		_w2099_,
		_w4952_
	);
	LUT3 #(
		.INIT('h70)
	) name4919 (
		_w2023_,
		_w2055_,
		_w3249_,
		_w4953_
	);
	LUT3 #(
		.INIT('h01)
	) name4920 (
		_w4952_,
		_w4953_,
		_w4951_,
		_w4954_
	);
	LUT4 #(
		.INIT('h95aa)
	) name4921 (
		\a[23] ,
		_w37_,
		_w4151_,
		_w4954_,
		_w4955_
	);
	LUT2 #(
		.INIT('h9)
	) name4922 (
		_w4806_,
		_w4808_,
		_w4956_
	);
	LUT2 #(
		.INIT('h4)
	) name4923 (
		_w4955_,
		_w4956_,
		_w4957_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4924 (
		_w1874_,
		_w2076_,
		_w2099_,
		_w3249_,
		_w4958_
	);
	LUT3 #(
		.INIT('h2a)
	) name4925 (
		_w3214_,
		_w2124_,
		_w2133_,
		_w4959_
	);
	LUT3 #(
		.INIT('h70)
	) name4926 (
		_w2023_,
		_w2055_,
		_w3262_,
		_w4960_
	);
	LUT3 #(
		.INIT('h01)
	) name4927 (
		_w4958_,
		_w4959_,
		_w4960_,
		_w4961_
	);
	LUT4 #(
		.INIT('h6f00)
	) name4928 (
		_w2299_,
		_w2301_,
		_w37_,
		_w4961_,
		_w4962_
	);
	LUT3 #(
		.INIT('h69)
	) name4929 (
		_w4608_,
		_w4800_,
		_w4805_,
		_w4963_
	);
	LUT3 #(
		.INIT('h90)
	) name4930 (
		\a[23] ,
		_w4962_,
		_w4963_,
		_w4964_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4931 (
		_w1874_,
		_w2076_,
		_w2099_,
		_w3262_,
		_w4965_
	);
	LUT3 #(
		.INIT('h70)
	) name4932 (
		_w2124_,
		_w2133_,
		_w3249_,
		_w4966_
	);
	LUT3 #(
		.INIT('h2a)
	) name4933 (
		_w3214_,
		_w2155_,
		_w2156_,
		_w4967_
	);
	LUT3 #(
		.INIT('h01)
	) name4934 (
		_w4965_,
		_w4966_,
		_w4967_,
		_w4968_
	);
	LUT4 #(
		.INIT('h95aa)
	) name4935 (
		\a[23] ,
		_w37_,
		_w4209_,
		_w4968_,
		_w4969_
	);
	LUT3 #(
		.INIT('h8a)
	) name4936 (
		\a[26] ,
		_w4792_,
		_w4791_,
		_w4970_
	);
	LUT2 #(
		.INIT('h9)
	) name4937 (
		_w4799_,
		_w4970_,
		_w4971_
	);
	LUT2 #(
		.INIT('h4)
	) name4938 (
		_w4969_,
		_w4971_,
		_w4972_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name4939 (
		_w3214_,
		_w2193_,
		_w2183_,
		_w2213_,
		_w4973_
	);
	LUT3 #(
		.INIT('h70)
	) name4940 (
		_w2155_,
		_w2156_,
		_w3249_,
		_w4974_
	);
	LUT3 #(
		.INIT('h70)
	) name4941 (
		_w2124_,
		_w2133_,
		_w3262_,
		_w4975_
	);
	LUT3 #(
		.INIT('h01)
	) name4942 (
		_w4973_,
		_w4974_,
		_w4975_,
		_w4976_
	);
	LUT4 #(
		.INIT('h6f00)
	) name4943 (
		_w2295_,
		_w2297_,
		_w37_,
		_w4976_,
		_w4977_
	);
	LUT4 #(
		.INIT('h002a)
	) name4944 (
		\a[26] ,
		_w2228_,
		_w2262_,
		_w2873_,
		_w4978_
	);
	LUT2 #(
		.INIT('h9)
	) name4945 (
		_w4791_,
		_w4978_,
		_w4979_
	);
	LUT3 #(
		.INIT('h90)
	) name4946 (
		\a[23] ,
		_w4977_,
		_w4979_,
		_w4980_
	);
	LUT3 #(
		.INIT('h70)
	) name4947 (
		_w2228_,
		_w2262_,
		_w3249_,
		_w4981_
	);
	LUT3 #(
		.INIT('h70)
	) name4948 (
		_w2273_,
		_w2293_,
		_w3262_,
		_w4982_
	);
	LUT4 #(
		.INIT('h000d)
	) name4949 (
		_w37_,
		_w4599_,
		_w4981_,
		_w4982_,
		_w4983_
	);
	LUT3 #(
		.INIT('h15)
	) name4950 (
		_w36_,
		_w2228_,
		_w2262_,
		_w4984_
	);
	LUT4 #(
		.INIT('ha888)
	) name4951 (
		\a[23] ,
		_w36_,
		_w2228_,
		_w2262_,
		_w4985_
	);
	LUT3 #(
		.INIT('h84)
	) name4952 (
		_w2214_,
		_w37_,
		_w4258_,
		_w4986_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4953 (
		_w2193_,
		_w2183_,
		_w2213_,
		_w3262_,
		_w4987_
	);
	LUT3 #(
		.INIT('h2a)
	) name4954 (
		_w3214_,
		_w2228_,
		_w2262_,
		_w4988_
	);
	LUT3 #(
		.INIT('h70)
	) name4955 (
		_w2273_,
		_w2293_,
		_w3249_,
		_w4989_
	);
	LUT3 #(
		.INIT('h01)
	) name4956 (
		_w4988_,
		_w4989_,
		_w4987_,
		_w4990_
	);
	LUT2 #(
		.INIT('h4)
	) name4957 (
		_w4986_,
		_w4990_,
		_w4991_
	);
	LUT4 #(
		.INIT('h0800)
	) name4958 (
		_w4983_,
		_w4985_,
		_w4986_,
		_w4990_,
		_w4992_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4959 (
		_w2193_,
		_w2183_,
		_w2213_,
		_w3249_,
		_w4993_
	);
	LUT3 #(
		.INIT('h70)
	) name4960 (
		_w2155_,
		_w2156_,
		_w3262_,
		_w4994_
	);
	LUT3 #(
		.INIT('h2a)
	) name4961 (
		_w3214_,
		_w2273_,
		_w2293_,
		_w4995_
	);
	LUT3 #(
		.INIT('h01)
	) name4962 (
		_w4993_,
		_w4994_,
		_w4995_,
		_w4996_
	);
	LUT4 #(
		.INIT('h95aa)
	) name4963 (
		\a[23] ,
		_w37_,
		_w4293_,
		_w4996_,
		_w4997_
	);
	LUT3 #(
		.INIT('h71)
	) name4964 (
		_w4792_,
		_w4992_,
		_w4997_,
		_w4998_
	);
	LUT3 #(
		.INIT('h06)
	) name4965 (
		\a[23] ,
		_w4977_,
		_w4979_,
		_w4999_
	);
	LUT3 #(
		.INIT('h69)
	) name4966 (
		\a[23] ,
		_w4977_,
		_w4979_,
		_w5000_
	);
	LUT3 #(
		.INIT('h54)
	) name4967 (
		_w4980_,
		_w4998_,
		_w4999_,
		_w5001_
	);
	LUT2 #(
		.INIT('h2)
	) name4968 (
		_w4969_,
		_w4971_,
		_w5002_
	);
	LUT2 #(
		.INIT('h9)
	) name4969 (
		_w4969_,
		_w4971_,
		_w5003_
	);
	LUT3 #(
		.INIT('h69)
	) name4970 (
		\a[23] ,
		_w4962_,
		_w4963_,
		_w5004_
	);
	LUT4 #(
		.INIT('h4d00)
	) name4971 (
		_w4969_,
		_w4971_,
		_w5001_,
		_w5004_,
		_w5005_
	);
	LUT2 #(
		.INIT('h2)
	) name4972 (
		_w4955_,
		_w4956_,
		_w5006_
	);
	LUT2 #(
		.INIT('h9)
	) name4973 (
		_w4955_,
		_w4956_,
		_w5007_
	);
	LUT4 #(
		.INIT('h5501)
	) name4974 (
		_w4957_,
		_w4964_,
		_w5005_,
		_w5006_,
		_w5008_
	);
	LUT4 #(
		.INIT('h1428)
	) name4975 (
		\a[23] ,
		_w4809_,
		_w4811_,
		_w4948_,
		_w5009_
	);
	LUT4 #(
		.INIT('h6996)
	) name4976 (
		\a[23] ,
		_w4809_,
		_w4811_,
		_w4948_,
		_w5010_
	);
	LUT2 #(
		.INIT('h9)
	) name4977 (
		_w4936_,
		_w4941_,
		_w5011_
	);
	LUT4 #(
		.INIT('h2b00)
	) name4978 (
		_w4943_,
		_w4949_,
		_w5008_,
		_w5011_,
		_w5012_
	);
	LUT2 #(
		.INIT('h2)
	) name4979 (
		_w4933_,
		_w4934_,
		_w5013_
	);
	LUT2 #(
		.INIT('h9)
	) name4980 (
		_w4933_,
		_w4934_,
		_w5014_
	);
	LUT4 #(
		.INIT('h5501)
	) name4981 (
		_w4935_,
		_w4942_,
		_w5012_,
		_w5013_,
		_w5015_
	);
	LUT3 #(
		.INIT('h60)
	) name4982 (
		_w4816_,
		_w4818_,
		_w4926_,
		_w5016_
	);
	LUT3 #(
		.INIT('h96)
	) name4983 (
		_w4816_,
		_w4818_,
		_w4926_,
		_w5017_
	);
	LUT2 #(
		.INIT('h9)
	) name4984 (
		_w4919_,
		_w4920_,
		_w5018_
	);
	LUT4 #(
		.INIT('hba00)
	) name4985 (
		_w4927_,
		_w5015_,
		_w5017_,
		_w5018_,
		_w5019_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name4986 (
		_w4750_,
		_w4820_,
		_w4822_,
		_w4912_,
		_w5020_
	);
	LUT4 #(
		.INIT('h0155)
	) name4987 (
		_w4913_,
		_w4921_,
		_w5019_,
		_w5020_,
		_w5021_
	);
	LUT3 #(
		.INIT('h60)
	) name4988 (
		_w4823_,
		_w4825_,
		_w4905_,
		_w5022_
	);
	LUT3 #(
		.INIT('h96)
	) name4989 (
		_w4823_,
		_w4825_,
		_w4905_,
		_w5023_
	);
	LUT2 #(
		.INIT('h9)
	) name4990 (
		_w4897_,
		_w4898_,
		_w5024_
	);
	LUT4 #(
		.INIT('h4d00)
	) name4991 (
		_w4905_,
		_w4906_,
		_w5021_,
		_w5024_,
		_w5025_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name4992 (
		_w4729_,
		_w4827_,
		_w4828_,
		_w4891_,
		_w5026_
	);
	LUT4 #(
		.INIT('h0155)
	) name4993 (
		_w4892_,
		_w4899_,
		_w5025_,
		_w5026_,
		_w5027_
	);
	LUT3 #(
		.INIT('h96)
	) name4994 (
		_w4829_,
		_w4830_,
		_w4835_,
		_w5028_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4995 (
		_w1454_,
		_w1426_,
		_w1478_,
		_w3311_,
		_w5029_
	);
	LUT3 #(
		.INIT('h70)
	) name4996 (
		_w1325_,
		_w1367_,
		_w3654_,
		_w5030_
	);
	LUT3 #(
		.INIT('h70)
	) name4997 (
		_w1381_,
		_w1398_,
		_w3645_,
		_w5031_
	);
	LUT3 #(
		.INIT('h01)
	) name4998 (
		_w5030_,
		_w5031_,
		_w5029_,
		_w5032_
	);
	LUT4 #(
		.INIT('h6f00)
	) name4999 (
		_w2327_,
		_w2329_,
		_w3312_,
		_w5032_,
		_w5033_
	);
	LUT2 #(
		.INIT('h6)
	) name5000 (
		\a[20] ,
		_w5033_,
		_w5034_
	);
	LUT4 #(
		.INIT('h4db2)
	) name5001 (
		_w4829_,
		_w4830_,
		_w4835_,
		_w4836_,
		_w5035_
	);
	LUT2 #(
		.INIT('h9)
	) name5002 (
		_w4843_,
		_w5035_,
		_w5036_
	);
	LUT4 #(
		.INIT('h4d00)
	) name5003 (
		_w5027_,
		_w5028_,
		_w5034_,
		_w5036_,
		_w5037_
	);
	LUT4 #(
		.INIT('h00b2)
	) name5004 (
		_w5027_,
		_w5028_,
		_w5034_,
		_w5036_,
		_w5038_
	);
	LUT3 #(
		.INIT('h70)
	) name5005 (
		_w1136_,
		_w1187_,
		_w3877_,
		_w5039_
	);
	LUT3 #(
		.INIT('h70)
	) name5006 (
		_w1071_,
		_w1102_,
		_w3886_,
		_w5040_
	);
	LUT3 #(
		.INIT('h70)
	) name5007 (
		_w1202_,
		_w1233_,
		_w3709_,
		_w5041_
	);
	LUT3 #(
		.INIT('h01)
	) name5008 (
		_w5040_,
		_w5041_,
		_w5039_,
		_w5042_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5009 (
		_w2335_,
		_w2337_,
		_w3710_,
		_w5042_,
		_w5043_
	);
	LUT2 #(
		.INIT('h6)
	) name5010 (
		\a[17] ,
		_w5043_,
		_w5044_
	);
	LUT3 #(
		.INIT('h54)
	) name5011 (
		_w5037_,
		_w5038_,
		_w5044_,
		_w5045_
	);
	LUT3 #(
		.INIT('h70)
	) name5012 (
		_w763_,
		_w983_,
		_w4033_,
		_w5046_
	);
	LUT3 #(
		.INIT('h70)
	) name5013 (
		_w871_,
		_w927_,
		_w4367_,
		_w5047_
	);
	LUT3 #(
		.INIT('h70)
	) name5014 (
		_w801_,
		_w851_,
		_w4382_,
		_w5048_
	);
	LUT3 #(
		.INIT('h01)
	) name5015 (
		_w5047_,
		_w5048_,
		_w5046_,
		_w5049_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5016 (
		_w2343_,
		_w2345_,
		_w4034_,
		_w5049_,
		_w5050_
	);
	LUT4 #(
		.INIT('h71b2)
	) name5017 (
		\a[14] ,
		_w4885_,
		_w5045_,
		_w5050_,
		_w5051_
	);
	LUT3 #(
		.INIT('hd4)
	) name5018 (
		_w4878_,
		_w4883_,
		_w5051_,
		_w5052_
	);
	LUT4 #(
		.INIT('h9669)
	) name5019 (
		\a[14] ,
		_w4853_,
		_w4855_,
		_w4860_,
		_w5053_
	);
	LUT2 #(
		.INIT('h4)
	) name5020 (
		_w5052_,
		_w5053_,
		_w5054_
	);
	LUT2 #(
		.INIT('h2)
	) name5021 (
		_w5052_,
		_w5053_,
		_w5055_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5022 (
		_w486_,
		_w487_,
		_w509_,
		_w4700_,
		_w5056_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5023 (
		_w587_,
		_w608_,
		_w624_,
		_w4458_,
		_w5057_
	);
	LUT3 #(
		.INIT('h70)
	) name5024 (
		_w544_,
		_w558_,
		_w4684_,
		_w5058_
	);
	LUT3 #(
		.INIT('h01)
	) name5025 (
		_w5056_,
		_w5057_,
		_w5058_,
		_w5059_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5026 (
		\a[11] ,
		_w2526_,
		_w4459_,
		_w5059_,
		_w5060_
	);
	LUT3 #(
		.INIT('h54)
	) name5027 (
		_w5054_,
		_w5055_,
		_w5060_,
		_w5061_
	);
	LUT3 #(
		.INIT('h96)
	) name5028 (
		_w4679_,
		_w4704_,
		_w4861_,
		_w5062_
	);
	LUT3 #(
		.INIT('h69)
	) name5029 (
		\a[11] ,
		_w4868_,
		_w5062_,
		_w5063_
	);
	LUT4 #(
		.INIT('h90f9)
	) name5030 (
		\a[8] ,
		_w4877_,
		_w5061_,
		_w5063_,
		_w5064_
	);
	LUT2 #(
		.INIT('h2)
	) name5031 (
		_w4873_,
		_w5064_,
		_w5065_
	);
	LUT2 #(
		.INIT('h4)
	) name5032 (
		_w4873_,
		_w5064_,
		_w5066_
	);
	LUT2 #(
		.INIT('h9)
	) name5033 (
		_w4873_,
		_w5064_,
		_w5067_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5034 (
		_w587_,
		_w608_,
		_w624_,
		_w4684_,
		_w5068_
	);
	LUT3 #(
		.INIT('h70)
	) name5035 (
		_w666_,
		_w694_,
		_w4458_,
		_w5069_
	);
	LUT3 #(
		.INIT('h70)
	) name5036 (
		_w544_,
		_w558_,
		_w4700_,
		_w5070_
	);
	LUT3 #(
		.INIT('h01)
	) name5037 (
		_w5069_,
		_w5070_,
		_w5068_,
		_w5071_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5038 (
		_w2351_,
		_w2353_,
		_w4459_,
		_w5071_,
		_w5072_
	);
	LUT2 #(
		.INIT('h6)
	) name5039 (
		\a[11] ,
		_w5072_,
		_w5073_
	);
	LUT4 #(
		.INIT('h6996)
	) name5040 (
		\a[14] ,
		_w4885_,
		_w5045_,
		_w5050_,
		_w5074_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5041 (
		_w1454_,
		_w1426_,
		_w1478_,
		_w3645_,
		_w5075_
	);
	LUT3 #(
		.INIT('h70)
	) name5042 (
		_w1381_,
		_w1398_,
		_w3654_,
		_w5076_
	);
	LUT3 #(
		.INIT('h70)
	) name5043 (
		_w1501_,
		_w1545_,
		_w3311_,
		_w5077_
	);
	LUT3 #(
		.INIT('h01)
	) name5044 (
		_w5076_,
		_w5077_,
		_w5075_,
		_w5078_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5045 (
		\a[20] ,
		_w3312_,
		_w3362_,
		_w5078_,
		_w5079_
	);
	LUT4 #(
		.INIT('h001e)
	) name5046 (
		_w4899_,
		_w5025_,
		_w5026_,
		_w5079_,
		_w5080_
	);
	LUT4 #(
		.INIT('h54ab)
	) name5047 (
		_w4907_,
		_w5021_,
		_w5022_,
		_w5024_,
		_w5081_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5048 (
		_w1454_,
		_w1426_,
		_w1478_,
		_w3654_,
		_w5082_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5049 (
		_w1584_,
		_w1569_,
		_w1606_,
		_w3311_,
		_w5083_
	);
	LUT3 #(
		.INIT('h70)
	) name5050 (
		_w1501_,
		_w1545_,
		_w3645_,
		_w5084_
	);
	LUT3 #(
		.INIT('h01)
	) name5051 (
		_w5083_,
		_w5084_,
		_w5082_,
		_w5085_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5052 (
		_w2323_,
		_w2325_,
		_w3312_,
		_w5085_,
		_w5086_
	);
	LUT2 #(
		.INIT('h6)
	) name5053 (
		\a[20] ,
		_w5086_,
		_w5087_
	);
	LUT2 #(
		.INIT('h2)
	) name5054 (
		_w5081_,
		_w5087_,
		_w5088_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5055 (
		_w1584_,
		_w1569_,
		_w1606_,
		_w3645_,
		_w5089_
	);
	LUT3 #(
		.INIT('h70)
	) name5056 (
		_w1501_,
		_w1545_,
		_w3654_,
		_w5090_
	);
	LUT3 #(
		.INIT('h70)
	) name5057 (
		_w1620_,
		_w1661_,
		_w3311_,
		_w5091_
	);
	LUT3 #(
		.INIT('h01)
	) name5058 (
		_w5089_,
		_w5090_,
		_w5091_,
		_w5092_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5059 (
		\a[20] ,
		_w3312_,
		_w3495_,
		_w5092_,
		_w5093_
	);
	LUT3 #(
		.INIT('h09)
	) name5060 (
		_w5021_,
		_w5023_,
		_w5093_,
		_w5094_
	);
	LUT3 #(
		.INIT('h70)
	) name5061 (
		_w1692_,
		_w1723_,
		_w3311_,
		_w5095_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5062 (
		_w1584_,
		_w1569_,
		_w1606_,
		_w3654_,
		_w5096_
	);
	LUT3 #(
		.INIT('h70)
	) name5063 (
		_w1620_,
		_w1661_,
		_w3645_,
		_w5097_
	);
	LUT3 #(
		.INIT('h01)
	) name5064 (
		_w5096_,
		_w5097_,
		_w5095_,
		_w5098_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5065 (
		_w2319_,
		_w2321_,
		_w3312_,
		_w5098_,
		_w5099_
	);
	LUT2 #(
		.INIT('h6)
	) name5066 (
		\a[20] ,
		_w5099_,
		_w5100_
	);
	LUT4 #(
		.INIT('h001e)
	) name5067 (
		_w4921_,
		_w5019_,
		_w5020_,
		_w5100_,
		_w5101_
	);
	LUT4 #(
		.INIT('h54ab)
	) name5068 (
		_w4927_,
		_w5015_,
		_w5016_,
		_w5018_,
		_w5102_
	);
	LUT3 #(
		.INIT('h70)
	) name5069 (
		_w1692_,
		_w1723_,
		_w3645_,
		_w5103_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5070 (
		_w1751_,
		_w1742_,
		_w1771_,
		_w3311_,
		_w5104_
	);
	LUT3 #(
		.INIT('h70)
	) name5071 (
		_w1620_,
		_w1661_,
		_w3654_,
		_w5105_
	);
	LUT3 #(
		.INIT('h01)
	) name5072 (
		_w5104_,
		_w5105_,
		_w5103_,
		_w5106_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5073 (
		\a[20] ,
		_w3312_,
		_w3599_,
		_w5106_,
		_w5107_
	);
	LUT2 #(
		.INIT('h2)
	) name5074 (
		_w5102_,
		_w5107_,
		_w5108_
	);
	LUT2 #(
		.INIT('h9)
	) name5075 (
		_w5015_,
		_w5017_,
		_w5109_
	);
	LUT3 #(
		.INIT('h70)
	) name5076 (
		_w1692_,
		_w1723_,
		_w3654_,
		_w5110_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5077 (
		_w1751_,
		_w1742_,
		_w1771_,
		_w3645_,
		_w5111_
	);
	LUT3 #(
		.INIT('h70)
	) name5078 (
		_w1795_,
		_w1796_,
		_w3311_,
		_w5112_
	);
	LUT3 #(
		.INIT('h01)
	) name5079 (
		_w5111_,
		_w5112_,
		_w5110_,
		_w5113_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5080 (
		_w2315_,
		_w2317_,
		_w3312_,
		_w5113_,
		_w5114_
	);
	LUT2 #(
		.INIT('h6)
	) name5081 (
		\a[20] ,
		_w5114_,
		_w5115_
	);
	LUT3 #(
		.INIT('h09)
	) name5082 (
		_w5015_,
		_w5017_,
		_w5115_,
		_w5116_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5083 (
		_w1751_,
		_w1742_,
		_w1771_,
		_w3654_,
		_w5117_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5084 (
		_w1817_,
		_w1799_,
		_w1840_,
		_w3311_,
		_w5118_
	);
	LUT3 #(
		.INIT('h70)
	) name5085 (
		_w1795_,
		_w1796_,
		_w3645_,
		_w5119_
	);
	LUT3 #(
		.INIT('h01)
	) name5086 (
		_w5118_,
		_w5119_,
		_w5117_,
		_w5120_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5087 (
		\a[20] ,
		_w3312_,
		_w3909_,
		_w5120_,
		_w5121_
	);
	LUT4 #(
		.INIT('h001e)
	) name5088 (
		_w4942_,
		_w5012_,
		_w5014_,
		_w5121_,
		_w5122_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5089 (
		_w1817_,
		_w1799_,
		_w1840_,
		_w3645_,
		_w5123_
	);
	LUT3 #(
		.INIT('h70)
	) name5090 (
		_w1795_,
		_w1796_,
		_w3654_,
		_w5124_
	);
	LUT3 #(
		.INIT('h70)
	) name5091 (
		_w1863_,
		_w1875_,
		_w3311_,
		_w5125_
	);
	LUT3 #(
		.INIT('h01)
	) name5092 (
		_w5124_,
		_w5125_,
		_w5123_,
		_w5126_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5093 (
		_w2311_,
		_w2313_,
		_w3312_,
		_w5126_,
		_w5127_
	);
	LUT2 #(
		.INIT('h6)
	) name5094 (
		\a[20] ,
		_w5127_,
		_w5128_
	);
	LUT4 #(
		.INIT('h54ab)
	) name5095 (
		_w4950_,
		_w5008_,
		_w5009_,
		_w5011_,
		_w5129_
	);
	LUT2 #(
		.INIT('h4)
	) name5096 (
		_w5128_,
		_w5129_,
		_w5130_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5097 (
		_w1817_,
		_w1799_,
		_w1840_,
		_w3654_,
		_w5131_
	);
	LUT3 #(
		.INIT('h70)
	) name5098 (
		_w1898_,
		_w1928_,
		_w3311_,
		_w5132_
	);
	LUT3 #(
		.INIT('h70)
	) name5099 (
		_w1863_,
		_w1875_,
		_w3645_,
		_w5133_
	);
	LUT3 #(
		.INIT('h01)
	) name5100 (
		_w5132_,
		_w5133_,
		_w5131_,
		_w5134_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5101 (
		\a[20] ,
		_w3312_,
		_w3972_,
		_w5134_,
		_w5135_
	);
	LUT3 #(
		.INIT('h09)
	) name5102 (
		_w5008_,
		_w5010_,
		_w5135_,
		_w5136_
	);
	LUT3 #(
		.INIT('h1e)
	) name5103 (
		_w4964_,
		_w5005_,
		_w5007_,
		_w5137_
	);
	LUT3 #(
		.INIT('h70)
	) name5104 (
		_w1501_,
		_w1949_,
		_w3311_,
		_w5138_
	);
	LUT3 #(
		.INIT('h70)
	) name5105 (
		_w1898_,
		_w1928_,
		_w3645_,
		_w5139_
	);
	LUT3 #(
		.INIT('h70)
	) name5106 (
		_w1863_,
		_w1875_,
		_w3654_,
		_w5140_
	);
	LUT3 #(
		.INIT('h01)
	) name5107 (
		_w5139_,
		_w5140_,
		_w5138_,
		_w5141_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5108 (
		_w2307_,
		_w2309_,
		_w3312_,
		_w5141_,
		_w5142_
	);
	LUT2 #(
		.INIT('h6)
	) name5109 (
		\a[20] ,
		_w5142_,
		_w5143_
	);
	LUT2 #(
		.INIT('h2)
	) name5110 (
		_w5137_,
		_w5143_,
		_w5144_
	);
	LUT4 #(
		.INIT('h54ab)
	) name5111 (
		_w4972_,
		_w5001_,
		_w5002_,
		_w5004_,
		_w5145_
	);
	LUT3 #(
		.INIT('h70)
	) name5112 (
		_w1973_,
		_w1997_,
		_w3311_,
		_w5146_
	);
	LUT3 #(
		.INIT('h70)
	) name5113 (
		_w1898_,
		_w1928_,
		_w3654_,
		_w5147_
	);
	LUT3 #(
		.INIT('h70)
	) name5114 (
		_w1501_,
		_w1949_,
		_w3645_,
		_w5148_
	);
	LUT3 #(
		.INIT('h01)
	) name5115 (
		_w5147_,
		_w5148_,
		_w5146_,
		_w5149_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5116 (
		\a[20] ,
		_w3312_,
		_w4126_,
		_w5149_,
		_w5150_
	);
	LUT2 #(
		.INIT('h2)
	) name5117 (
		_w5145_,
		_w5150_,
		_w5151_
	);
	LUT2 #(
		.INIT('h9)
	) name5118 (
		_w5001_,
		_w5003_,
		_w5152_
	);
	LUT3 #(
		.INIT('h70)
	) name5119 (
		_w1973_,
		_w1997_,
		_w3645_,
		_w5153_
	);
	LUT3 #(
		.INIT('h70)
	) name5120 (
		_w1501_,
		_w1949_,
		_w3654_,
		_w5154_
	);
	LUT3 #(
		.INIT('h70)
	) name5121 (
		_w2023_,
		_w2055_,
		_w3311_,
		_w5155_
	);
	LUT3 #(
		.INIT('h01)
	) name5122 (
		_w5154_,
		_w5155_,
		_w5153_,
		_w5156_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5123 (
		_w2303_,
		_w2305_,
		_w3312_,
		_w5156_,
		_w5157_
	);
	LUT2 #(
		.INIT('h6)
	) name5124 (
		\a[20] ,
		_w5157_,
		_w5158_
	);
	LUT4 #(
		.INIT('h8241)
	) name5125 (
		\a[20] ,
		_w5001_,
		_w5003_,
		_w5157_,
		_w5159_
	);
	LUT3 #(
		.INIT('h70)
	) name5126 (
		_w1973_,
		_w1997_,
		_w3654_,
		_w5160_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5127 (
		_w1874_,
		_w2076_,
		_w2099_,
		_w3311_,
		_w5161_
	);
	LUT3 #(
		.INIT('h70)
	) name5128 (
		_w2023_,
		_w2055_,
		_w3645_,
		_w5162_
	);
	LUT3 #(
		.INIT('h01)
	) name5129 (
		_w5161_,
		_w5162_,
		_w5160_,
		_w5163_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5130 (
		\a[20] ,
		_w3312_,
		_w4151_,
		_w5163_,
		_w5164_
	);
	LUT2 #(
		.INIT('h9)
	) name5131 (
		_w4998_,
		_w5000_,
		_w5165_
	);
	LUT2 #(
		.INIT('h4)
	) name5132 (
		_w5164_,
		_w5165_,
		_w5166_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5133 (
		_w1874_,
		_w2076_,
		_w2099_,
		_w3645_,
		_w5167_
	);
	LUT3 #(
		.INIT('h70)
	) name5134 (
		_w2124_,
		_w2133_,
		_w3311_,
		_w5168_
	);
	LUT3 #(
		.INIT('h70)
	) name5135 (
		_w2023_,
		_w2055_,
		_w3654_,
		_w5169_
	);
	LUT3 #(
		.INIT('h01)
	) name5136 (
		_w5167_,
		_w5168_,
		_w5169_,
		_w5170_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5137 (
		_w2299_,
		_w2301_,
		_w3312_,
		_w5170_,
		_w5171_
	);
	LUT3 #(
		.INIT('h69)
	) name5138 (
		_w4792_,
		_w4992_,
		_w4997_,
		_w5172_
	);
	LUT3 #(
		.INIT('h90)
	) name5139 (
		\a[20] ,
		_w5171_,
		_w5172_,
		_w5173_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5140 (
		_w1874_,
		_w2076_,
		_w2099_,
		_w3654_,
		_w5174_
	);
	LUT3 #(
		.INIT('h70)
	) name5141 (
		_w2124_,
		_w2133_,
		_w3645_,
		_w5175_
	);
	LUT3 #(
		.INIT('h70)
	) name5142 (
		_w2155_,
		_w2156_,
		_w3311_,
		_w5176_
	);
	LUT3 #(
		.INIT('h01)
	) name5143 (
		_w5174_,
		_w5175_,
		_w5176_,
		_w5177_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5144 (
		\a[20] ,
		_w3312_,
		_w4209_,
		_w5177_,
		_w5178_
	);
	LUT3 #(
		.INIT('h8a)
	) name5145 (
		\a[23] ,
		_w4984_,
		_w4983_,
		_w5179_
	);
	LUT2 #(
		.INIT('h9)
	) name5146 (
		_w4991_,
		_w5179_,
		_w5180_
	);
	LUT2 #(
		.INIT('h4)
	) name5147 (
		_w5178_,
		_w5180_,
		_w5181_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5148 (
		_w2193_,
		_w2183_,
		_w2213_,
		_w3311_,
		_w5182_
	);
	LUT3 #(
		.INIT('h70)
	) name5149 (
		_w2155_,
		_w2156_,
		_w3645_,
		_w5183_
	);
	LUT3 #(
		.INIT('h70)
	) name5150 (
		_w2124_,
		_w2133_,
		_w3654_,
		_w5184_
	);
	LUT3 #(
		.INIT('h01)
	) name5151 (
		_w5182_,
		_w5183_,
		_w5184_,
		_w5185_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5152 (
		_w2295_,
		_w2297_,
		_w3312_,
		_w5185_,
		_w5186_
	);
	LUT4 #(
		.INIT('h0222)
	) name5153 (
		\a[23] ,
		_w36_,
		_w2228_,
		_w2262_,
		_w5187_
	);
	LUT2 #(
		.INIT('h9)
	) name5154 (
		_w4983_,
		_w5187_,
		_w5188_
	);
	LUT3 #(
		.INIT('h90)
	) name5155 (
		\a[20] ,
		_w5186_,
		_w5188_,
		_w5189_
	);
	LUT3 #(
		.INIT('h70)
	) name5156 (
		_w2228_,
		_w2262_,
		_w3645_,
		_w5190_
	);
	LUT3 #(
		.INIT('h70)
	) name5157 (
		_w2273_,
		_w2293_,
		_w3654_,
		_w5191_
	);
	LUT4 #(
		.INIT('h000d)
	) name5158 (
		_w3312_,
		_w4599_,
		_w5190_,
		_w5191_,
		_w5192_
	);
	LUT3 #(
		.INIT('h07)
	) name5159 (
		_w2228_,
		_w2262_,
		_w3310_,
		_w5193_
	);
	LUT4 #(
		.INIT('haa80)
	) name5160 (
		\a[20] ,
		_w2228_,
		_w2262_,
		_w3310_,
		_w5194_
	);
	LUT3 #(
		.INIT('h84)
	) name5161 (
		_w2214_,
		_w3312_,
		_w4258_,
		_w5195_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5162 (
		_w2193_,
		_w2183_,
		_w2213_,
		_w3654_,
		_w5196_
	);
	LUT3 #(
		.INIT('h70)
	) name5163 (
		_w2228_,
		_w2262_,
		_w3311_,
		_w5197_
	);
	LUT3 #(
		.INIT('h70)
	) name5164 (
		_w2273_,
		_w2293_,
		_w3645_,
		_w5198_
	);
	LUT3 #(
		.INIT('h01)
	) name5165 (
		_w5197_,
		_w5198_,
		_w5196_,
		_w5199_
	);
	LUT2 #(
		.INIT('h4)
	) name5166 (
		_w5195_,
		_w5199_,
		_w5200_
	);
	LUT4 #(
		.INIT('h0800)
	) name5167 (
		_w5192_,
		_w5194_,
		_w5195_,
		_w5199_,
		_w5201_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5168 (
		_w2193_,
		_w2183_,
		_w2213_,
		_w3645_,
		_w5202_
	);
	LUT3 #(
		.INIT('h70)
	) name5169 (
		_w2155_,
		_w2156_,
		_w3654_,
		_w5203_
	);
	LUT3 #(
		.INIT('h70)
	) name5170 (
		_w2273_,
		_w2293_,
		_w3311_,
		_w5204_
	);
	LUT3 #(
		.INIT('h01)
	) name5171 (
		_w5202_,
		_w5203_,
		_w5204_,
		_w5205_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5172 (
		\a[20] ,
		_w3312_,
		_w4293_,
		_w5205_,
		_w5206_
	);
	LUT3 #(
		.INIT('h71)
	) name5173 (
		_w4984_,
		_w5201_,
		_w5206_,
		_w5207_
	);
	LUT3 #(
		.INIT('h06)
	) name5174 (
		\a[20] ,
		_w5186_,
		_w5188_,
		_w5208_
	);
	LUT3 #(
		.INIT('h69)
	) name5175 (
		\a[20] ,
		_w5186_,
		_w5188_,
		_w5209_
	);
	LUT3 #(
		.INIT('h54)
	) name5176 (
		_w5189_,
		_w5207_,
		_w5208_,
		_w5210_
	);
	LUT2 #(
		.INIT('h2)
	) name5177 (
		_w5178_,
		_w5180_,
		_w5211_
	);
	LUT2 #(
		.INIT('h9)
	) name5178 (
		_w5178_,
		_w5180_,
		_w5212_
	);
	LUT3 #(
		.INIT('h69)
	) name5179 (
		\a[20] ,
		_w5171_,
		_w5172_,
		_w5213_
	);
	LUT4 #(
		.INIT('h4d00)
	) name5180 (
		_w5178_,
		_w5180_,
		_w5210_,
		_w5213_,
		_w5214_
	);
	LUT2 #(
		.INIT('h2)
	) name5181 (
		_w5164_,
		_w5165_,
		_w5215_
	);
	LUT2 #(
		.INIT('h9)
	) name5182 (
		_w5164_,
		_w5165_,
		_w5216_
	);
	LUT4 #(
		.INIT('h5501)
	) name5183 (
		_w5166_,
		_w5173_,
		_w5214_,
		_w5215_,
		_w5217_
	);
	LUT4 #(
		.INIT('h1428)
	) name5184 (
		\a[20] ,
		_w5001_,
		_w5003_,
		_w5157_,
		_w5218_
	);
	LUT4 #(
		.INIT('h6996)
	) name5185 (
		\a[20] ,
		_w5001_,
		_w5003_,
		_w5157_,
		_w5219_
	);
	LUT2 #(
		.INIT('h9)
	) name5186 (
		_w5145_,
		_w5150_,
		_w5220_
	);
	LUT4 #(
		.INIT('h2b00)
	) name5187 (
		_w5152_,
		_w5158_,
		_w5217_,
		_w5220_,
		_w5221_
	);
	LUT2 #(
		.INIT('h4)
	) name5188 (
		_w5137_,
		_w5143_,
		_w5222_
	);
	LUT2 #(
		.INIT('h9)
	) name5189 (
		_w5137_,
		_w5143_,
		_w5223_
	);
	LUT4 #(
		.INIT('h5501)
	) name5190 (
		_w5144_,
		_w5151_,
		_w5221_,
		_w5222_,
		_w5224_
	);
	LUT3 #(
		.INIT('h60)
	) name5191 (
		_w5008_,
		_w5010_,
		_w5135_,
		_w5225_
	);
	LUT3 #(
		.INIT('h96)
	) name5192 (
		_w5008_,
		_w5010_,
		_w5135_,
		_w5226_
	);
	LUT2 #(
		.INIT('h9)
	) name5193 (
		_w5128_,
		_w5129_,
		_w5227_
	);
	LUT4 #(
		.INIT('hba00)
	) name5194 (
		_w5136_,
		_w5224_,
		_w5226_,
		_w5227_,
		_w5228_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name5195 (
		_w4942_,
		_w5012_,
		_w5014_,
		_w5121_,
		_w5229_
	);
	LUT4 #(
		.INIT('h0155)
	) name5196 (
		_w5122_,
		_w5130_,
		_w5228_,
		_w5229_,
		_w5230_
	);
	LUT3 #(
		.INIT('h60)
	) name5197 (
		_w5015_,
		_w5017_,
		_w5115_,
		_w5231_
	);
	LUT3 #(
		.INIT('h96)
	) name5198 (
		_w5015_,
		_w5017_,
		_w5115_,
		_w5232_
	);
	LUT2 #(
		.INIT('h9)
	) name5199 (
		_w5102_,
		_w5107_,
		_w5233_
	);
	LUT4 #(
		.INIT('h2b00)
	) name5200 (
		_w5109_,
		_w5115_,
		_w5230_,
		_w5233_,
		_w5234_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name5201 (
		_w4921_,
		_w5019_,
		_w5020_,
		_w5100_,
		_w5235_
	);
	LUT4 #(
		.INIT('h0155)
	) name5202 (
		_w5101_,
		_w5108_,
		_w5234_,
		_w5235_,
		_w5236_
	);
	LUT3 #(
		.INIT('h60)
	) name5203 (
		_w5021_,
		_w5023_,
		_w5093_,
		_w5237_
	);
	LUT3 #(
		.INIT('h96)
	) name5204 (
		_w5021_,
		_w5023_,
		_w5093_,
		_w5238_
	);
	LUT2 #(
		.INIT('h9)
	) name5205 (
		_w5081_,
		_w5087_,
		_w5239_
	);
	LUT4 #(
		.INIT('hba00)
	) name5206 (
		_w5094_,
		_w5236_,
		_w5238_,
		_w5239_,
		_w5240_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name5207 (
		_w4899_,
		_w5025_,
		_w5026_,
		_w5079_,
		_w5241_
	);
	LUT4 #(
		.INIT('h0155)
	) name5208 (
		_w5080_,
		_w5088_,
		_w5240_,
		_w5241_,
		_w5242_
	);
	LUT3 #(
		.INIT('h96)
	) name5209 (
		_w5027_,
		_w5028_,
		_w5034_,
		_w5243_
	);
	LUT3 #(
		.INIT('h70)
	) name5210 (
		_w1202_,
		_w1233_,
		_w3877_,
		_w5244_
	);
	LUT3 #(
		.INIT('h70)
	) name5211 (
		_w1253_,
		_w1294_,
		_w3709_,
		_w5245_
	);
	LUT3 #(
		.INIT('h70)
	) name5212 (
		_w1136_,
		_w1187_,
		_w3886_,
		_w5246_
	);
	LUT3 #(
		.INIT('h01)
	) name5213 (
		_w5245_,
		_w5246_,
		_w5244_,
		_w5247_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5214 (
		\a[17] ,
		_w3067_,
		_w3710_,
		_w5247_,
		_w5248_
	);
	LUT3 #(
		.INIT('hb2)
	) name5215 (
		_w5242_,
		_w5243_,
		_w5248_,
		_w5249_
	);
	LUT4 #(
		.INIT('hb24d)
	) name5216 (
		_w5027_,
		_w5028_,
		_w5034_,
		_w5036_,
		_w5250_
	);
	LUT2 #(
		.INIT('h6)
	) name5217 (
		_w5044_,
		_w5250_,
		_w5251_
	);
	LUT4 #(
		.INIT('h004d)
	) name5218 (
		_w5242_,
		_w5243_,
		_w5248_,
		_w5251_,
		_w5252_
	);
	LUT4 #(
		.INIT('hb200)
	) name5219 (
		_w5242_,
		_w5243_,
		_w5248_,
		_w5251_,
		_w5253_
	);
	LUT3 #(
		.INIT('h70)
	) name5220 (
		_w1009_,
		_w1050_,
		_w4033_,
		_w5254_
	);
	LUT3 #(
		.INIT('h70)
	) name5221 (
		_w871_,
		_w927_,
		_w4382_,
		_w5255_
	);
	LUT3 #(
		.INIT('h70)
	) name5222 (
		_w763_,
		_w983_,
		_w4367_,
		_w5256_
	);
	LUT3 #(
		.INIT('h01)
	) name5223 (
		_w5255_,
		_w5256_,
		_w5254_,
		_w5257_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5224 (
		\a[14] ,
		_w2839_,
		_w4034_,
		_w5257_,
		_w5258_
	);
	LUT4 #(
		.INIT('h022a)
	) name5225 (
		_w5074_,
		_w5249_,
		_w5251_,
		_w5258_,
		_w5259_
	);
	LUT4 #(
		.INIT('h5440)
	) name5226 (
		_w5074_,
		_w5249_,
		_w5251_,
		_w5258_,
		_w5260_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5227 (
		_w587_,
		_w608_,
		_w624_,
		_w4700_,
		_w5261_
	);
	LUT3 #(
		.INIT('h70)
	) name5228 (
		_w725_,
		_w764_,
		_w4458_,
		_w5262_
	);
	LUT3 #(
		.INIT('h70)
	) name5229 (
		_w666_,
		_w694_,
		_w4684_,
		_w5263_
	);
	LUT3 #(
		.INIT('h01)
	) name5230 (
		_w5262_,
		_w5263_,
		_w5261_,
		_w5264_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5231 (
		\a[11] ,
		_w2598_,
		_w4459_,
		_w5264_,
		_w5265_
	);
	LUT3 #(
		.INIT('h54)
	) name5232 (
		_w5259_,
		_w5260_,
		_w5265_,
		_w5266_
	);
	LUT3 #(
		.INIT('h96)
	) name5233 (
		_w4878_,
		_w4883_,
		_w5051_,
		_w5267_
	);
	LUT3 #(
		.INIT('h8e)
	) name5234 (
		_w5073_,
		_w5266_,
		_w5267_,
		_w5268_
	);
	LUT4 #(
		.INIT('hf400)
	) name5235 (
		_w374_,
		_w2361_,
		_w2404_,
		_w4876_,
		_w5269_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5236 (
		_w121_,
		_w418_,
		_w422_,
		_w4875_,
		_w5270_
	);
	LUT3 #(
		.INIT('h18)
	) name5237 (
		\a[5] ,
		\a[6] ,
		\a[7] ,
		_w5271_
	);
	LUT3 #(
		.INIT('h70)
	) name5238 (
		_w352_,
		_w373_,
		_w5271_,
		_w5272_
	);
	LUT2 #(
		.INIT('h1)
	) name5239 (
		_w5270_,
		_w5272_,
		_w5273_
	);
	LUT3 #(
		.INIT('h9a)
	) name5240 (
		\a[8] ,
		_w5269_,
		_w5273_,
		_w5274_
	);
	LUT4 #(
		.INIT('h1211)
	) name5241 (
		\a[8] ,
		_w5268_,
		_w5269_,
		_w5273_,
		_w5275_
	);
	LUT4 #(
		.INIT('h8488)
	) name5242 (
		\a[8] ,
		_w5268_,
		_w5269_,
		_w5273_,
		_w5276_
	);
	LUT4 #(
		.INIT('h6966)
	) name5243 (
		\a[8] ,
		_w5268_,
		_w5269_,
		_w5273_,
		_w5277_
	);
	LUT2 #(
		.INIT('h9)
	) name5244 (
		_w5052_,
		_w5053_,
		_w5278_
	);
	LUT2 #(
		.INIT('h6)
	) name5245 (
		_w5060_,
		_w5278_,
		_w5279_
	);
	LUT3 #(
		.INIT('h54)
	) name5246 (
		_w5275_,
		_w5276_,
		_w5279_,
		_w5280_
	);
	LUT4 #(
		.INIT('h9669)
	) name5247 (
		\a[8] ,
		_w4877_,
		_w5061_,
		_w5063_,
		_w5281_
	);
	LUT4 #(
		.INIT('h1700)
	) name5248 (
		_w5268_,
		_w5274_,
		_w5279_,
		_w5281_,
		_w5282_
	);
	LUT4 #(
		.INIT('h54ab)
	) name5249 (
		_w5275_,
		_w5276_,
		_w5279_,
		_w5281_,
		_w5283_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5250 (
		_w486_,
		_w487_,
		_w509_,
		_w4875_,
		_w5284_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5251 (
		_w121_,
		_w418_,
		_w422_,
		_w5271_,
		_w5285_
	);
	LUT4 #(
		.INIT('h6006)
	) name5252 (
		\a[5] ,
		\a[6] ,
		\a[7] ,
		\a[8] ,
		_w5286_
	);
	LUT3 #(
		.INIT('h70)
	) name5253 (
		_w352_,
		_w373_,
		_w5286_,
		_w5287_
	);
	LUT3 #(
		.INIT('h01)
	) name5254 (
		_w5284_,
		_w5285_,
		_w5287_,
		_w5288_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5255 (
		\a[8] ,
		_w2535_,
		_w4876_,
		_w5288_,
		_w5289_
	);
	LUT4 #(
		.INIT('h6665)
	) name5256 (
		_w5074_,
		_w5252_,
		_w5253_,
		_w5258_,
		_w5290_
	);
	LUT2 #(
		.INIT('h9)
	) name5257 (
		_w5265_,
		_w5290_,
		_w5291_
	);
	LUT3 #(
		.INIT('h70)
	) name5258 (
		_w1202_,
		_w1233_,
		_w3886_,
		_w5292_
	);
	LUT3 #(
		.INIT('h70)
	) name5259 (
		_w1325_,
		_w1367_,
		_w3709_,
		_w5293_
	);
	LUT3 #(
		.INIT('h70)
	) name5260 (
		_w1253_,
		_w1294_,
		_w3877_,
		_w5294_
	);
	LUT3 #(
		.INIT('h01)
	) name5261 (
		_w5293_,
		_w5294_,
		_w5292_,
		_w5295_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5262 (
		_w2331_,
		_w2333_,
		_w3710_,
		_w5295_,
		_w5296_
	);
	LUT2 #(
		.INIT('h6)
	) name5263 (
		\a[17] ,
		_w5296_,
		_w5297_
	);
	LUT4 #(
		.INIT('h001e)
	) name5264 (
		_w5088_,
		_w5240_,
		_w5241_,
		_w5297_,
		_w5298_
	);
	LUT3 #(
		.INIT('h70)
	) name5265 (
		_w1381_,
		_w1398_,
		_w3709_,
		_w5299_
	);
	LUT3 #(
		.INIT('h70)
	) name5266 (
		_w1325_,
		_w1367_,
		_w3877_,
		_w5300_
	);
	LUT3 #(
		.INIT('h70)
	) name5267 (
		_w1253_,
		_w1294_,
		_w3886_,
		_w5301_
	);
	LUT3 #(
		.INIT('h01)
	) name5268 (
		_w5300_,
		_w5301_,
		_w5299_,
		_w5302_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5269 (
		\a[17] ,
		_w3182_,
		_w3710_,
		_w5302_,
		_w5303_
	);
	LUT4 #(
		.INIT('h54ab)
	) name5270 (
		_w5094_,
		_w5236_,
		_w5237_,
		_w5239_,
		_w5304_
	);
	LUT2 #(
		.INIT('h4)
	) name5271 (
		_w5303_,
		_w5304_,
		_w5305_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5272 (
		_w1454_,
		_w1426_,
		_w1478_,
		_w3709_,
		_w5306_
	);
	LUT3 #(
		.INIT('h70)
	) name5273 (
		_w1325_,
		_w1367_,
		_w3886_,
		_w5307_
	);
	LUT3 #(
		.INIT('h70)
	) name5274 (
		_w1381_,
		_w1398_,
		_w3877_,
		_w5308_
	);
	LUT3 #(
		.INIT('h01)
	) name5275 (
		_w5307_,
		_w5308_,
		_w5306_,
		_w5309_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5276 (
		_w2327_,
		_w2329_,
		_w3710_,
		_w5309_,
		_w5310_
	);
	LUT2 #(
		.INIT('h6)
	) name5277 (
		\a[17] ,
		_w5310_,
		_w5311_
	);
	LUT2 #(
		.INIT('h9)
	) name5278 (
		_w5236_,
		_w5238_,
		_w5312_
	);
	LUT3 #(
		.INIT('h09)
	) name5279 (
		_w5236_,
		_w5238_,
		_w5311_,
		_w5313_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5280 (
		_w1454_,
		_w1426_,
		_w1478_,
		_w3877_,
		_w5314_
	);
	LUT3 #(
		.INIT('h70)
	) name5281 (
		_w1381_,
		_w1398_,
		_w3886_,
		_w5315_
	);
	LUT3 #(
		.INIT('h70)
	) name5282 (
		_w1501_,
		_w1545_,
		_w3709_,
		_w5316_
	);
	LUT3 #(
		.INIT('h01)
	) name5283 (
		_w5315_,
		_w5316_,
		_w5314_,
		_w5317_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5284 (
		\a[17] ,
		_w3362_,
		_w3710_,
		_w5317_,
		_w5318_
	);
	LUT4 #(
		.INIT('h001e)
	) name5285 (
		_w5108_,
		_w5234_,
		_w5235_,
		_w5318_,
		_w5319_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5286 (
		_w1454_,
		_w1426_,
		_w1478_,
		_w3886_,
		_w5320_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5287 (
		_w1584_,
		_w1569_,
		_w1606_,
		_w3709_,
		_w5321_
	);
	LUT3 #(
		.INIT('h70)
	) name5288 (
		_w1501_,
		_w1545_,
		_w3877_,
		_w5322_
	);
	LUT3 #(
		.INIT('h01)
	) name5289 (
		_w5321_,
		_w5322_,
		_w5320_,
		_w5323_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5290 (
		_w2323_,
		_w2325_,
		_w3710_,
		_w5323_,
		_w5324_
	);
	LUT2 #(
		.INIT('h6)
	) name5291 (
		\a[17] ,
		_w5324_,
		_w5325_
	);
	LUT4 #(
		.INIT('h54ab)
	) name5292 (
		_w5116_,
		_w5230_,
		_w5231_,
		_w5233_,
		_w5326_
	);
	LUT2 #(
		.INIT('h4)
	) name5293 (
		_w5325_,
		_w5326_,
		_w5327_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5294 (
		_w1584_,
		_w1569_,
		_w1606_,
		_w3877_,
		_w5328_
	);
	LUT3 #(
		.INIT('h70)
	) name5295 (
		_w1501_,
		_w1545_,
		_w3886_,
		_w5329_
	);
	LUT3 #(
		.INIT('h70)
	) name5296 (
		_w1620_,
		_w1661_,
		_w3709_,
		_w5330_
	);
	LUT3 #(
		.INIT('h01)
	) name5297 (
		_w5328_,
		_w5329_,
		_w5330_,
		_w5331_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5298 (
		\a[17] ,
		_w3495_,
		_w3710_,
		_w5331_,
		_w5332_
	);
	LUT3 #(
		.INIT('h09)
	) name5299 (
		_w5230_,
		_w5232_,
		_w5332_,
		_w5333_
	);
	LUT3 #(
		.INIT('h70)
	) name5300 (
		_w1692_,
		_w1723_,
		_w3709_,
		_w5334_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5301 (
		_w1584_,
		_w1569_,
		_w1606_,
		_w3886_,
		_w5335_
	);
	LUT3 #(
		.INIT('h70)
	) name5302 (
		_w1620_,
		_w1661_,
		_w3877_,
		_w5336_
	);
	LUT3 #(
		.INIT('h01)
	) name5303 (
		_w5335_,
		_w5336_,
		_w5334_,
		_w5337_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5304 (
		_w2319_,
		_w2321_,
		_w3710_,
		_w5337_,
		_w5338_
	);
	LUT2 #(
		.INIT('h6)
	) name5305 (
		\a[17] ,
		_w5338_,
		_w5339_
	);
	LUT4 #(
		.INIT('h001e)
	) name5306 (
		_w5130_,
		_w5228_,
		_w5229_,
		_w5339_,
		_w5340_
	);
	LUT4 #(
		.INIT('h54ab)
	) name5307 (
		_w5136_,
		_w5224_,
		_w5225_,
		_w5227_,
		_w5341_
	);
	LUT3 #(
		.INIT('h70)
	) name5308 (
		_w1692_,
		_w1723_,
		_w3877_,
		_w5342_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5309 (
		_w1751_,
		_w1742_,
		_w1771_,
		_w3709_,
		_w5343_
	);
	LUT3 #(
		.INIT('h70)
	) name5310 (
		_w1620_,
		_w1661_,
		_w3886_,
		_w5344_
	);
	LUT3 #(
		.INIT('h01)
	) name5311 (
		_w5343_,
		_w5344_,
		_w5342_,
		_w5345_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5312 (
		\a[17] ,
		_w3599_,
		_w3710_,
		_w5345_,
		_w5346_
	);
	LUT2 #(
		.INIT('h2)
	) name5313 (
		_w5341_,
		_w5346_,
		_w5347_
	);
	LUT2 #(
		.INIT('h9)
	) name5314 (
		_w5224_,
		_w5226_,
		_w5348_
	);
	LUT3 #(
		.INIT('h70)
	) name5315 (
		_w1692_,
		_w1723_,
		_w3886_,
		_w5349_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5316 (
		_w1751_,
		_w1742_,
		_w1771_,
		_w3877_,
		_w5350_
	);
	LUT3 #(
		.INIT('h70)
	) name5317 (
		_w1795_,
		_w1796_,
		_w3709_,
		_w5351_
	);
	LUT3 #(
		.INIT('h01)
	) name5318 (
		_w5350_,
		_w5351_,
		_w5349_,
		_w5352_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5319 (
		_w2315_,
		_w2317_,
		_w3710_,
		_w5352_,
		_w5353_
	);
	LUT2 #(
		.INIT('h6)
	) name5320 (
		\a[17] ,
		_w5353_,
		_w5354_
	);
	LUT3 #(
		.INIT('h09)
	) name5321 (
		_w5224_,
		_w5226_,
		_w5354_,
		_w5355_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5322 (
		_w1751_,
		_w1742_,
		_w1771_,
		_w3886_,
		_w5356_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5323 (
		_w1817_,
		_w1799_,
		_w1840_,
		_w3709_,
		_w5357_
	);
	LUT3 #(
		.INIT('h70)
	) name5324 (
		_w1795_,
		_w1796_,
		_w3877_,
		_w5358_
	);
	LUT3 #(
		.INIT('h01)
	) name5325 (
		_w5357_,
		_w5358_,
		_w5356_,
		_w5359_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5326 (
		\a[17] ,
		_w3710_,
		_w3909_,
		_w5359_,
		_w5360_
	);
	LUT4 #(
		.INIT('h001e)
	) name5327 (
		_w5151_,
		_w5221_,
		_w5223_,
		_w5360_,
		_w5361_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5328 (
		_w1817_,
		_w1799_,
		_w1840_,
		_w3877_,
		_w5362_
	);
	LUT3 #(
		.INIT('h70)
	) name5329 (
		_w1795_,
		_w1796_,
		_w3886_,
		_w5363_
	);
	LUT3 #(
		.INIT('h70)
	) name5330 (
		_w1863_,
		_w1875_,
		_w3709_,
		_w5364_
	);
	LUT3 #(
		.INIT('h01)
	) name5331 (
		_w5363_,
		_w5364_,
		_w5362_,
		_w5365_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5332 (
		_w2311_,
		_w2313_,
		_w3710_,
		_w5365_,
		_w5366_
	);
	LUT2 #(
		.INIT('h6)
	) name5333 (
		\a[17] ,
		_w5366_,
		_w5367_
	);
	LUT4 #(
		.INIT('h54ab)
	) name5334 (
		_w5159_,
		_w5217_,
		_w5218_,
		_w5220_,
		_w5368_
	);
	LUT2 #(
		.INIT('h4)
	) name5335 (
		_w5367_,
		_w5368_,
		_w5369_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5336 (
		_w1817_,
		_w1799_,
		_w1840_,
		_w3886_,
		_w5370_
	);
	LUT3 #(
		.INIT('h70)
	) name5337 (
		_w1898_,
		_w1928_,
		_w3709_,
		_w5371_
	);
	LUT3 #(
		.INIT('h70)
	) name5338 (
		_w1863_,
		_w1875_,
		_w3877_,
		_w5372_
	);
	LUT3 #(
		.INIT('h01)
	) name5339 (
		_w5371_,
		_w5372_,
		_w5370_,
		_w5373_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5340 (
		\a[17] ,
		_w3710_,
		_w3972_,
		_w5373_,
		_w5374_
	);
	LUT3 #(
		.INIT('h09)
	) name5341 (
		_w5217_,
		_w5219_,
		_w5374_,
		_w5375_
	);
	LUT3 #(
		.INIT('h1e)
	) name5342 (
		_w5173_,
		_w5214_,
		_w5216_,
		_w5376_
	);
	LUT3 #(
		.INIT('h70)
	) name5343 (
		_w1501_,
		_w1949_,
		_w3709_,
		_w5377_
	);
	LUT3 #(
		.INIT('h70)
	) name5344 (
		_w1898_,
		_w1928_,
		_w3877_,
		_w5378_
	);
	LUT3 #(
		.INIT('h70)
	) name5345 (
		_w1863_,
		_w1875_,
		_w3886_,
		_w5379_
	);
	LUT3 #(
		.INIT('h01)
	) name5346 (
		_w5378_,
		_w5379_,
		_w5377_,
		_w5380_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5347 (
		_w2307_,
		_w2309_,
		_w3710_,
		_w5380_,
		_w5381_
	);
	LUT2 #(
		.INIT('h6)
	) name5348 (
		\a[17] ,
		_w5381_,
		_w5382_
	);
	LUT2 #(
		.INIT('h2)
	) name5349 (
		_w5376_,
		_w5382_,
		_w5383_
	);
	LUT4 #(
		.INIT('h54ab)
	) name5350 (
		_w5181_,
		_w5210_,
		_w5211_,
		_w5213_,
		_w5384_
	);
	LUT3 #(
		.INIT('h70)
	) name5351 (
		_w1973_,
		_w1997_,
		_w3709_,
		_w5385_
	);
	LUT3 #(
		.INIT('h70)
	) name5352 (
		_w1898_,
		_w1928_,
		_w3886_,
		_w5386_
	);
	LUT3 #(
		.INIT('h70)
	) name5353 (
		_w1501_,
		_w1949_,
		_w3877_,
		_w5387_
	);
	LUT3 #(
		.INIT('h01)
	) name5354 (
		_w5386_,
		_w5387_,
		_w5385_,
		_w5388_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5355 (
		\a[17] ,
		_w3710_,
		_w4126_,
		_w5388_,
		_w5389_
	);
	LUT2 #(
		.INIT('h2)
	) name5356 (
		_w5384_,
		_w5389_,
		_w5390_
	);
	LUT2 #(
		.INIT('h9)
	) name5357 (
		_w5210_,
		_w5212_,
		_w5391_
	);
	LUT3 #(
		.INIT('h70)
	) name5358 (
		_w1973_,
		_w1997_,
		_w3877_,
		_w5392_
	);
	LUT3 #(
		.INIT('h70)
	) name5359 (
		_w1501_,
		_w1949_,
		_w3886_,
		_w5393_
	);
	LUT3 #(
		.INIT('h70)
	) name5360 (
		_w2023_,
		_w2055_,
		_w3709_,
		_w5394_
	);
	LUT3 #(
		.INIT('h01)
	) name5361 (
		_w5393_,
		_w5394_,
		_w5392_,
		_w5395_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5362 (
		_w2303_,
		_w2305_,
		_w3710_,
		_w5395_,
		_w5396_
	);
	LUT2 #(
		.INIT('h6)
	) name5363 (
		\a[17] ,
		_w5396_,
		_w5397_
	);
	LUT4 #(
		.INIT('h8241)
	) name5364 (
		\a[17] ,
		_w5210_,
		_w5212_,
		_w5396_,
		_w5398_
	);
	LUT3 #(
		.INIT('h70)
	) name5365 (
		_w1973_,
		_w1997_,
		_w3886_,
		_w5399_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5366 (
		_w1874_,
		_w2076_,
		_w2099_,
		_w3709_,
		_w5400_
	);
	LUT3 #(
		.INIT('h70)
	) name5367 (
		_w2023_,
		_w2055_,
		_w3877_,
		_w5401_
	);
	LUT3 #(
		.INIT('h01)
	) name5368 (
		_w5400_,
		_w5401_,
		_w5399_,
		_w5402_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5369 (
		\a[17] ,
		_w3710_,
		_w4151_,
		_w5402_,
		_w5403_
	);
	LUT2 #(
		.INIT('h9)
	) name5370 (
		_w5207_,
		_w5209_,
		_w5404_
	);
	LUT2 #(
		.INIT('h4)
	) name5371 (
		_w5403_,
		_w5404_,
		_w5405_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5372 (
		_w1874_,
		_w2076_,
		_w2099_,
		_w3877_,
		_w5406_
	);
	LUT3 #(
		.INIT('h70)
	) name5373 (
		_w2124_,
		_w2133_,
		_w3709_,
		_w5407_
	);
	LUT3 #(
		.INIT('h70)
	) name5374 (
		_w2023_,
		_w2055_,
		_w3886_,
		_w5408_
	);
	LUT3 #(
		.INIT('h01)
	) name5375 (
		_w5406_,
		_w5407_,
		_w5408_,
		_w5409_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5376 (
		_w2299_,
		_w2301_,
		_w3710_,
		_w5409_,
		_w5410_
	);
	LUT3 #(
		.INIT('h69)
	) name5377 (
		_w4984_,
		_w5201_,
		_w5206_,
		_w5411_
	);
	LUT3 #(
		.INIT('h90)
	) name5378 (
		\a[17] ,
		_w5410_,
		_w5411_,
		_w5412_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5379 (
		_w1874_,
		_w2076_,
		_w2099_,
		_w3886_,
		_w5413_
	);
	LUT3 #(
		.INIT('h70)
	) name5380 (
		_w2124_,
		_w2133_,
		_w3877_,
		_w5414_
	);
	LUT3 #(
		.INIT('h70)
	) name5381 (
		_w2155_,
		_w2156_,
		_w3709_,
		_w5415_
	);
	LUT3 #(
		.INIT('h01)
	) name5382 (
		_w5413_,
		_w5414_,
		_w5415_,
		_w5416_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5383 (
		\a[17] ,
		_w3710_,
		_w4209_,
		_w5416_,
		_w5417_
	);
	LUT3 #(
		.INIT('h8a)
	) name5384 (
		\a[20] ,
		_w5193_,
		_w5192_,
		_w5418_
	);
	LUT2 #(
		.INIT('h9)
	) name5385 (
		_w5200_,
		_w5418_,
		_w5419_
	);
	LUT2 #(
		.INIT('h4)
	) name5386 (
		_w5417_,
		_w5419_,
		_w5420_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5387 (
		_w2193_,
		_w2183_,
		_w2213_,
		_w3709_,
		_w5421_
	);
	LUT3 #(
		.INIT('h70)
	) name5388 (
		_w2155_,
		_w2156_,
		_w3877_,
		_w5422_
	);
	LUT3 #(
		.INIT('h70)
	) name5389 (
		_w2124_,
		_w2133_,
		_w3886_,
		_w5423_
	);
	LUT3 #(
		.INIT('h01)
	) name5390 (
		_w5421_,
		_w5422_,
		_w5423_,
		_w5424_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5391 (
		_w2295_,
		_w2297_,
		_w3710_,
		_w5424_,
		_w5425_
	);
	LUT4 #(
		.INIT('h002a)
	) name5392 (
		\a[20] ,
		_w2228_,
		_w2262_,
		_w3310_,
		_w5426_
	);
	LUT2 #(
		.INIT('h9)
	) name5393 (
		_w5192_,
		_w5426_,
		_w5427_
	);
	LUT3 #(
		.INIT('h90)
	) name5394 (
		\a[17] ,
		_w5425_,
		_w5427_,
		_w5428_
	);
	LUT3 #(
		.INIT('h70)
	) name5395 (
		_w2228_,
		_w2262_,
		_w3877_,
		_w5429_
	);
	LUT3 #(
		.INIT('h70)
	) name5396 (
		_w2273_,
		_w2293_,
		_w3886_,
		_w5430_
	);
	LUT4 #(
		.INIT('h000d)
	) name5397 (
		_w3710_,
		_w4599_,
		_w5429_,
		_w5430_,
		_w5431_
	);
	LUT3 #(
		.INIT('h07)
	) name5398 (
		_w2228_,
		_w2262_,
		_w3708_,
		_w5432_
	);
	LUT4 #(
		.INIT('haa80)
	) name5399 (
		\a[17] ,
		_w2228_,
		_w2262_,
		_w3708_,
		_w5433_
	);
	LUT3 #(
		.INIT('h84)
	) name5400 (
		_w2214_,
		_w3710_,
		_w4258_,
		_w5434_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5401 (
		_w2193_,
		_w2183_,
		_w2213_,
		_w3886_,
		_w5435_
	);
	LUT3 #(
		.INIT('h70)
	) name5402 (
		_w2228_,
		_w2262_,
		_w3709_,
		_w5436_
	);
	LUT3 #(
		.INIT('h70)
	) name5403 (
		_w2273_,
		_w2293_,
		_w3877_,
		_w5437_
	);
	LUT3 #(
		.INIT('h01)
	) name5404 (
		_w5436_,
		_w5437_,
		_w5435_,
		_w5438_
	);
	LUT2 #(
		.INIT('h4)
	) name5405 (
		_w5434_,
		_w5438_,
		_w5439_
	);
	LUT4 #(
		.INIT('h0800)
	) name5406 (
		_w5431_,
		_w5433_,
		_w5434_,
		_w5438_,
		_w5440_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5407 (
		_w2193_,
		_w2183_,
		_w2213_,
		_w3877_,
		_w5441_
	);
	LUT3 #(
		.INIT('h70)
	) name5408 (
		_w2155_,
		_w2156_,
		_w3886_,
		_w5442_
	);
	LUT3 #(
		.INIT('h70)
	) name5409 (
		_w2273_,
		_w2293_,
		_w3709_,
		_w5443_
	);
	LUT3 #(
		.INIT('h01)
	) name5410 (
		_w5441_,
		_w5442_,
		_w5443_,
		_w5444_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5411 (
		\a[17] ,
		_w3710_,
		_w4293_,
		_w5444_,
		_w5445_
	);
	LUT3 #(
		.INIT('h71)
	) name5412 (
		_w5193_,
		_w5440_,
		_w5445_,
		_w5446_
	);
	LUT3 #(
		.INIT('h06)
	) name5413 (
		\a[17] ,
		_w5425_,
		_w5427_,
		_w5447_
	);
	LUT3 #(
		.INIT('h69)
	) name5414 (
		\a[17] ,
		_w5425_,
		_w5427_,
		_w5448_
	);
	LUT3 #(
		.INIT('h54)
	) name5415 (
		_w5428_,
		_w5446_,
		_w5447_,
		_w5449_
	);
	LUT2 #(
		.INIT('h2)
	) name5416 (
		_w5417_,
		_w5419_,
		_w5450_
	);
	LUT2 #(
		.INIT('h9)
	) name5417 (
		_w5417_,
		_w5419_,
		_w5451_
	);
	LUT3 #(
		.INIT('h69)
	) name5418 (
		\a[17] ,
		_w5410_,
		_w5411_,
		_w5452_
	);
	LUT4 #(
		.INIT('h4d00)
	) name5419 (
		_w5417_,
		_w5419_,
		_w5449_,
		_w5452_,
		_w5453_
	);
	LUT2 #(
		.INIT('h2)
	) name5420 (
		_w5403_,
		_w5404_,
		_w5454_
	);
	LUT2 #(
		.INIT('h9)
	) name5421 (
		_w5403_,
		_w5404_,
		_w5455_
	);
	LUT4 #(
		.INIT('h5501)
	) name5422 (
		_w5405_,
		_w5412_,
		_w5453_,
		_w5454_,
		_w5456_
	);
	LUT4 #(
		.INIT('h1428)
	) name5423 (
		\a[17] ,
		_w5210_,
		_w5212_,
		_w5396_,
		_w5457_
	);
	LUT4 #(
		.INIT('h6996)
	) name5424 (
		\a[17] ,
		_w5210_,
		_w5212_,
		_w5396_,
		_w5458_
	);
	LUT2 #(
		.INIT('h9)
	) name5425 (
		_w5384_,
		_w5389_,
		_w5459_
	);
	LUT4 #(
		.INIT('h2b00)
	) name5426 (
		_w5391_,
		_w5397_,
		_w5456_,
		_w5459_,
		_w5460_
	);
	LUT2 #(
		.INIT('h4)
	) name5427 (
		_w5376_,
		_w5382_,
		_w5461_
	);
	LUT2 #(
		.INIT('h9)
	) name5428 (
		_w5376_,
		_w5382_,
		_w5462_
	);
	LUT4 #(
		.INIT('h5501)
	) name5429 (
		_w5383_,
		_w5390_,
		_w5460_,
		_w5461_,
		_w5463_
	);
	LUT3 #(
		.INIT('h60)
	) name5430 (
		_w5217_,
		_w5219_,
		_w5374_,
		_w5464_
	);
	LUT3 #(
		.INIT('h96)
	) name5431 (
		_w5217_,
		_w5219_,
		_w5374_,
		_w5465_
	);
	LUT2 #(
		.INIT('h9)
	) name5432 (
		_w5367_,
		_w5368_,
		_w5466_
	);
	LUT4 #(
		.INIT('hba00)
	) name5433 (
		_w5375_,
		_w5463_,
		_w5465_,
		_w5466_,
		_w5467_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name5434 (
		_w5151_,
		_w5221_,
		_w5223_,
		_w5360_,
		_w5468_
	);
	LUT4 #(
		.INIT('h0155)
	) name5435 (
		_w5361_,
		_w5369_,
		_w5467_,
		_w5468_,
		_w5469_
	);
	LUT3 #(
		.INIT('h60)
	) name5436 (
		_w5224_,
		_w5226_,
		_w5354_,
		_w5470_
	);
	LUT3 #(
		.INIT('h96)
	) name5437 (
		_w5224_,
		_w5226_,
		_w5354_,
		_w5471_
	);
	LUT2 #(
		.INIT('h9)
	) name5438 (
		_w5341_,
		_w5346_,
		_w5472_
	);
	LUT4 #(
		.INIT('h2b00)
	) name5439 (
		_w5348_,
		_w5354_,
		_w5469_,
		_w5472_,
		_w5473_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name5440 (
		_w5130_,
		_w5228_,
		_w5229_,
		_w5339_,
		_w5474_
	);
	LUT4 #(
		.INIT('h0155)
	) name5441 (
		_w5340_,
		_w5347_,
		_w5473_,
		_w5474_,
		_w5475_
	);
	LUT3 #(
		.INIT('h60)
	) name5442 (
		_w5230_,
		_w5232_,
		_w5332_,
		_w5476_
	);
	LUT3 #(
		.INIT('h96)
	) name5443 (
		_w5230_,
		_w5232_,
		_w5332_,
		_w5477_
	);
	LUT2 #(
		.INIT('h9)
	) name5444 (
		_w5325_,
		_w5326_,
		_w5478_
	);
	LUT4 #(
		.INIT('hba00)
	) name5445 (
		_w5333_,
		_w5475_,
		_w5477_,
		_w5478_,
		_w5479_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name5446 (
		_w5108_,
		_w5234_,
		_w5235_,
		_w5318_,
		_w5480_
	);
	LUT4 #(
		.INIT('h0155)
	) name5447 (
		_w5319_,
		_w5327_,
		_w5479_,
		_w5480_,
		_w5481_
	);
	LUT3 #(
		.INIT('h60)
	) name5448 (
		_w5236_,
		_w5238_,
		_w5311_,
		_w5482_
	);
	LUT3 #(
		.INIT('h96)
	) name5449 (
		_w5236_,
		_w5238_,
		_w5311_,
		_w5483_
	);
	LUT2 #(
		.INIT('h9)
	) name5450 (
		_w5303_,
		_w5304_,
		_w5484_
	);
	LUT4 #(
		.INIT('h4d00)
	) name5451 (
		_w5311_,
		_w5312_,
		_w5481_,
		_w5484_,
		_w5485_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name5452 (
		_w5088_,
		_w5240_,
		_w5241_,
		_w5297_,
		_w5486_
	);
	LUT4 #(
		.INIT('h0155)
	) name5453 (
		_w5298_,
		_w5305_,
		_w5485_,
		_w5486_,
		_w5487_
	);
	LUT3 #(
		.INIT('h96)
	) name5454 (
		_w5242_,
		_w5243_,
		_w5248_,
		_w5488_
	);
	LUT3 #(
		.INIT('h70)
	) name5455 (
		_w1071_,
		_w1102_,
		_w4033_,
		_w5489_
	);
	LUT3 #(
		.INIT('h70)
	) name5456 (
		_w763_,
		_w983_,
		_w4382_,
		_w5490_
	);
	LUT3 #(
		.INIT('h70)
	) name5457 (
		_w1009_,
		_w1050_,
		_w4367_,
		_w5491_
	);
	LUT3 #(
		.INIT('h01)
	) name5458 (
		_w5490_,
		_w5491_,
		_w5489_,
		_w5492_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5459 (
		_w2339_,
		_w2341_,
		_w4034_,
		_w5492_,
		_w5493_
	);
	LUT2 #(
		.INIT('h6)
	) name5460 (
		\a[14] ,
		_w5493_,
		_w5494_
	);
	LUT3 #(
		.INIT('hb2)
	) name5461 (
		_w5487_,
		_w5488_,
		_w5494_,
		_w5495_
	);
	LUT4 #(
		.INIT('h4db2)
	) name5462 (
		_w5242_,
		_w5243_,
		_w5248_,
		_w5251_,
		_w5496_
	);
	LUT2 #(
		.INIT('h9)
	) name5463 (
		_w5258_,
		_w5496_,
		_w5497_
	);
	LUT4 #(
		.INIT('h4d00)
	) name5464 (
		_w5487_,
		_w5488_,
		_w5494_,
		_w5497_,
		_w5498_
	);
	LUT4 #(
		.INIT('h00b2)
	) name5465 (
		_w5487_,
		_w5488_,
		_w5494_,
		_w5497_,
		_w5499_
	);
	LUT3 #(
		.INIT('h70)
	) name5466 (
		_w725_,
		_w764_,
		_w4684_,
		_w5500_
	);
	LUT3 #(
		.INIT('h70)
	) name5467 (
		_w801_,
		_w851_,
		_w4458_,
		_w5501_
	);
	LUT3 #(
		.INIT('h70)
	) name5468 (
		_w666_,
		_w694_,
		_w4700_,
		_w5502_
	);
	LUT3 #(
		.INIT('h01)
	) name5469 (
		_w5501_,
		_w5502_,
		_w5500_,
		_w5503_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5470 (
		_w2347_,
		_w2349_,
		_w4459_,
		_w5503_,
		_w5504_
	);
	LUT2 #(
		.INIT('h6)
	) name5471 (
		\a[11] ,
		_w5504_,
		_w5505_
	);
	LUT3 #(
		.INIT('h54)
	) name5472 (
		_w5498_,
		_w5499_,
		_w5505_,
		_w5506_
	);
	LUT4 #(
		.INIT('h20a2)
	) name5473 (
		_w5291_,
		_w5495_,
		_w5497_,
		_w5505_,
		_w5507_
	);
	LUT4 #(
		.INIT('h4504)
	) name5474 (
		_w5291_,
		_w5495_,
		_w5497_,
		_w5505_,
		_w5508_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5475 (
		_w486_,
		_w487_,
		_w509_,
		_w5271_,
		_w5509_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5476 (
		_w121_,
		_w418_,
		_w422_,
		_w5286_,
		_w5510_
	);
	LUT3 #(
		.INIT('h70)
	) name5477 (
		_w544_,
		_w558_,
		_w4875_,
		_w5511_
	);
	LUT3 #(
		.INIT('h01)
	) name5478 (
		_w5509_,
		_w5510_,
		_w5511_,
		_w5512_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5479 (
		_w2355_,
		_w2357_,
		_w4876_,
		_w5512_,
		_w5513_
	);
	LUT2 #(
		.INIT('h6)
	) name5480 (
		\a[8] ,
		_w5513_,
		_w5514_
	);
	LUT4 #(
		.INIT('h0445)
	) name5481 (
		_w5289_,
		_w5291_,
		_w5506_,
		_w5514_,
		_w5515_
	);
	LUT3 #(
		.INIT('h96)
	) name5482 (
		_w5073_,
		_w5266_,
		_w5267_,
		_w5516_
	);
	LUT4 #(
		.INIT('ha220)
	) name5483 (
		_w5289_,
		_w5291_,
		_w5506_,
		_w5514_,
		_w5517_
	);
	LUT4 #(
		.INIT('h999a)
	) name5484 (
		_w5289_,
		_w5507_,
		_w5508_,
		_w5514_,
		_w5518_
	);
	LUT3 #(
		.INIT('h51)
	) name5485 (
		_w5515_,
		_w5516_,
		_w5517_,
		_w5519_
	);
	LUT2 #(
		.INIT('h9)
	) name5486 (
		_w5277_,
		_w5279_,
		_w5520_
	);
	LUT2 #(
		.INIT('h4)
	) name5487 (
		_w5519_,
		_w5520_,
		_w5521_
	);
	LUT2 #(
		.INIT('h6)
	) name5488 (
		_w5516_,
		_w5518_,
		_w5522_
	);
	LUT4 #(
		.INIT('h0990)
	) name5489 (
		\a[2] ,
		\a[3] ,
		\a[4] ,
		\a[5] ,
		_w5523_
	);
	LUT4 #(
		.INIT('h0180)
	) name5490 (
		\a[2] ,
		\a[3] ,
		\a[4] ,
		\a[5] ,
		_w5524_
	);
	LUT4 #(
		.INIT('h5150)
	) name5491 (
		_w374_,
		_w2361_,
		_w5524_,
		_w35_,
		_w5525_
	);
	LUT2 #(
		.INIT('h9)
	) name5492 (
		\a[5] ,
		_w5525_,
		_w5526_
	);
	LUT3 #(
		.INIT('h70)
	) name5493 (
		_w1136_,
		_w1187_,
		_w4033_,
		_w5527_
	);
	LUT3 #(
		.INIT('h70)
	) name5494 (
		_w1009_,
		_w1050_,
		_w4382_,
		_w5528_
	);
	LUT3 #(
		.INIT('h70)
	) name5495 (
		_w1071_,
		_w1102_,
		_w4367_,
		_w5529_
	);
	LUT3 #(
		.INIT('h01)
	) name5496 (
		_w5528_,
		_w5529_,
		_w5527_,
		_w5530_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5497 (
		\a[14] ,
		_w2936_,
		_w4034_,
		_w5530_,
		_w5531_
	);
	LUT4 #(
		.INIT('h001e)
	) name5498 (
		_w5305_,
		_w5485_,
		_w5486_,
		_w5531_,
		_w5532_
	);
	LUT4 #(
		.INIT('h54ab)
	) name5499 (
		_w5313_,
		_w5481_,
		_w5482_,
		_w5484_,
		_w5533_
	);
	LUT3 #(
		.INIT('h70)
	) name5500 (
		_w1136_,
		_w1187_,
		_w4367_,
		_w5534_
	);
	LUT3 #(
		.INIT('h70)
	) name5501 (
		_w1071_,
		_w1102_,
		_w4382_,
		_w5535_
	);
	LUT3 #(
		.INIT('h70)
	) name5502 (
		_w1202_,
		_w1233_,
		_w4033_,
		_w5536_
	);
	LUT3 #(
		.INIT('h01)
	) name5503 (
		_w5535_,
		_w5536_,
		_w5534_,
		_w5537_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5504 (
		_w2335_,
		_w2337_,
		_w4034_,
		_w5537_,
		_w5538_
	);
	LUT2 #(
		.INIT('h6)
	) name5505 (
		\a[14] ,
		_w5538_,
		_w5539_
	);
	LUT2 #(
		.INIT('h2)
	) name5506 (
		_w5533_,
		_w5539_,
		_w5540_
	);
	LUT3 #(
		.INIT('h70)
	) name5507 (
		_w1202_,
		_w1233_,
		_w4367_,
		_w5541_
	);
	LUT3 #(
		.INIT('h70)
	) name5508 (
		_w1253_,
		_w1294_,
		_w4033_,
		_w5542_
	);
	LUT3 #(
		.INIT('h70)
	) name5509 (
		_w1136_,
		_w1187_,
		_w4382_,
		_w5543_
	);
	LUT3 #(
		.INIT('h01)
	) name5510 (
		_w5542_,
		_w5543_,
		_w5541_,
		_w5544_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5511 (
		\a[14] ,
		_w3067_,
		_w4034_,
		_w5544_,
		_w5545_
	);
	LUT3 #(
		.INIT('h09)
	) name5512 (
		_w5481_,
		_w5483_,
		_w5545_,
		_w5546_
	);
	LUT3 #(
		.INIT('h70)
	) name5513 (
		_w1202_,
		_w1233_,
		_w4382_,
		_w5547_
	);
	LUT3 #(
		.INIT('h70)
	) name5514 (
		_w1325_,
		_w1367_,
		_w4033_,
		_w5548_
	);
	LUT3 #(
		.INIT('h70)
	) name5515 (
		_w1253_,
		_w1294_,
		_w4367_,
		_w5549_
	);
	LUT3 #(
		.INIT('h01)
	) name5516 (
		_w5548_,
		_w5549_,
		_w5547_,
		_w5550_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5517 (
		_w2331_,
		_w2333_,
		_w4034_,
		_w5550_,
		_w5551_
	);
	LUT2 #(
		.INIT('h6)
	) name5518 (
		\a[14] ,
		_w5551_,
		_w5552_
	);
	LUT4 #(
		.INIT('h001e)
	) name5519 (
		_w5327_,
		_w5479_,
		_w5480_,
		_w5552_,
		_w5553_
	);
	LUT4 #(
		.INIT('h54ab)
	) name5520 (
		_w5333_,
		_w5475_,
		_w5476_,
		_w5478_,
		_w5554_
	);
	LUT3 #(
		.INIT('h70)
	) name5521 (
		_w1381_,
		_w1398_,
		_w4033_,
		_w5555_
	);
	LUT3 #(
		.INIT('h70)
	) name5522 (
		_w1325_,
		_w1367_,
		_w4367_,
		_w5556_
	);
	LUT3 #(
		.INIT('h70)
	) name5523 (
		_w1253_,
		_w1294_,
		_w4382_,
		_w5557_
	);
	LUT3 #(
		.INIT('h01)
	) name5524 (
		_w5556_,
		_w5557_,
		_w5555_,
		_w5558_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5525 (
		\a[14] ,
		_w3182_,
		_w4034_,
		_w5558_,
		_w5559_
	);
	LUT2 #(
		.INIT('h2)
	) name5526 (
		_w5554_,
		_w5559_,
		_w5560_
	);
	LUT2 #(
		.INIT('h9)
	) name5527 (
		_w5475_,
		_w5477_,
		_w5561_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5528 (
		_w1454_,
		_w1426_,
		_w1478_,
		_w4033_,
		_w5562_
	);
	LUT3 #(
		.INIT('h70)
	) name5529 (
		_w1325_,
		_w1367_,
		_w4382_,
		_w5563_
	);
	LUT3 #(
		.INIT('h70)
	) name5530 (
		_w1381_,
		_w1398_,
		_w4367_,
		_w5564_
	);
	LUT3 #(
		.INIT('h01)
	) name5531 (
		_w5563_,
		_w5564_,
		_w5562_,
		_w5565_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5532 (
		_w2327_,
		_w2329_,
		_w4034_,
		_w5565_,
		_w5566_
	);
	LUT2 #(
		.INIT('h6)
	) name5533 (
		\a[14] ,
		_w5566_,
		_w5567_
	);
	LUT3 #(
		.INIT('h09)
	) name5534 (
		_w5475_,
		_w5477_,
		_w5567_,
		_w5568_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5535 (
		_w1454_,
		_w1426_,
		_w1478_,
		_w4367_,
		_w5569_
	);
	LUT3 #(
		.INIT('h70)
	) name5536 (
		_w1381_,
		_w1398_,
		_w4382_,
		_w5570_
	);
	LUT3 #(
		.INIT('h70)
	) name5537 (
		_w1501_,
		_w1545_,
		_w4033_,
		_w5571_
	);
	LUT3 #(
		.INIT('h01)
	) name5538 (
		_w5570_,
		_w5571_,
		_w5569_,
		_w5572_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5539 (
		\a[14] ,
		_w3362_,
		_w4034_,
		_w5572_,
		_w5573_
	);
	LUT4 #(
		.INIT('h001e)
	) name5540 (
		_w5347_,
		_w5473_,
		_w5474_,
		_w5573_,
		_w5574_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5541 (
		_w1454_,
		_w1426_,
		_w1478_,
		_w4382_,
		_w5575_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5542 (
		_w1584_,
		_w1569_,
		_w1606_,
		_w4033_,
		_w5576_
	);
	LUT3 #(
		.INIT('h70)
	) name5543 (
		_w1501_,
		_w1545_,
		_w4367_,
		_w5577_
	);
	LUT3 #(
		.INIT('h01)
	) name5544 (
		_w5576_,
		_w5577_,
		_w5575_,
		_w5578_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5545 (
		_w2323_,
		_w2325_,
		_w4034_,
		_w5578_,
		_w5579_
	);
	LUT2 #(
		.INIT('h6)
	) name5546 (
		\a[14] ,
		_w5579_,
		_w5580_
	);
	LUT4 #(
		.INIT('h54ab)
	) name5547 (
		_w5355_,
		_w5469_,
		_w5470_,
		_w5472_,
		_w5581_
	);
	LUT2 #(
		.INIT('h4)
	) name5548 (
		_w5580_,
		_w5581_,
		_w5582_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5549 (
		_w1584_,
		_w1569_,
		_w1606_,
		_w4367_,
		_w5583_
	);
	LUT3 #(
		.INIT('h70)
	) name5550 (
		_w1501_,
		_w1545_,
		_w4382_,
		_w5584_
	);
	LUT3 #(
		.INIT('h70)
	) name5551 (
		_w1620_,
		_w1661_,
		_w4033_,
		_w5585_
	);
	LUT3 #(
		.INIT('h01)
	) name5552 (
		_w5583_,
		_w5584_,
		_w5585_,
		_w5586_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5553 (
		\a[14] ,
		_w3495_,
		_w4034_,
		_w5586_,
		_w5587_
	);
	LUT3 #(
		.INIT('h09)
	) name5554 (
		_w5469_,
		_w5471_,
		_w5587_,
		_w5588_
	);
	LUT3 #(
		.INIT('h70)
	) name5555 (
		_w1692_,
		_w1723_,
		_w4033_,
		_w5589_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5556 (
		_w1584_,
		_w1569_,
		_w1606_,
		_w4382_,
		_w5590_
	);
	LUT3 #(
		.INIT('h70)
	) name5557 (
		_w1620_,
		_w1661_,
		_w4367_,
		_w5591_
	);
	LUT3 #(
		.INIT('h01)
	) name5558 (
		_w5590_,
		_w5591_,
		_w5589_,
		_w5592_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5559 (
		_w2319_,
		_w2321_,
		_w4034_,
		_w5592_,
		_w5593_
	);
	LUT2 #(
		.INIT('h6)
	) name5560 (
		\a[14] ,
		_w5593_,
		_w5594_
	);
	LUT4 #(
		.INIT('h001e)
	) name5561 (
		_w5369_,
		_w5467_,
		_w5468_,
		_w5594_,
		_w5595_
	);
	LUT4 #(
		.INIT('h54ab)
	) name5562 (
		_w5375_,
		_w5463_,
		_w5464_,
		_w5466_,
		_w5596_
	);
	LUT3 #(
		.INIT('h70)
	) name5563 (
		_w1692_,
		_w1723_,
		_w4367_,
		_w5597_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5564 (
		_w1751_,
		_w1742_,
		_w1771_,
		_w4033_,
		_w5598_
	);
	LUT3 #(
		.INIT('h70)
	) name5565 (
		_w1620_,
		_w1661_,
		_w4382_,
		_w5599_
	);
	LUT3 #(
		.INIT('h01)
	) name5566 (
		_w5598_,
		_w5599_,
		_w5597_,
		_w5600_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5567 (
		\a[14] ,
		_w3599_,
		_w4034_,
		_w5600_,
		_w5601_
	);
	LUT2 #(
		.INIT('h2)
	) name5568 (
		_w5596_,
		_w5601_,
		_w5602_
	);
	LUT2 #(
		.INIT('h9)
	) name5569 (
		_w5463_,
		_w5465_,
		_w5603_
	);
	LUT3 #(
		.INIT('h70)
	) name5570 (
		_w1692_,
		_w1723_,
		_w4382_,
		_w5604_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5571 (
		_w1751_,
		_w1742_,
		_w1771_,
		_w4367_,
		_w5605_
	);
	LUT3 #(
		.INIT('h70)
	) name5572 (
		_w1795_,
		_w1796_,
		_w4033_,
		_w5606_
	);
	LUT3 #(
		.INIT('h01)
	) name5573 (
		_w5605_,
		_w5606_,
		_w5604_,
		_w5607_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5574 (
		_w2315_,
		_w2317_,
		_w4034_,
		_w5607_,
		_w5608_
	);
	LUT2 #(
		.INIT('h6)
	) name5575 (
		\a[14] ,
		_w5608_,
		_w5609_
	);
	LUT3 #(
		.INIT('h09)
	) name5576 (
		_w5463_,
		_w5465_,
		_w5609_,
		_w5610_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5577 (
		_w1751_,
		_w1742_,
		_w1771_,
		_w4382_,
		_w5611_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5578 (
		_w1817_,
		_w1799_,
		_w1840_,
		_w4033_,
		_w5612_
	);
	LUT3 #(
		.INIT('h70)
	) name5579 (
		_w1795_,
		_w1796_,
		_w4367_,
		_w5613_
	);
	LUT3 #(
		.INIT('h01)
	) name5580 (
		_w5612_,
		_w5613_,
		_w5611_,
		_w5614_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5581 (
		\a[14] ,
		_w3909_,
		_w4034_,
		_w5614_,
		_w5615_
	);
	LUT4 #(
		.INIT('h001e)
	) name5582 (
		_w5390_,
		_w5460_,
		_w5462_,
		_w5615_,
		_w5616_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5583 (
		_w1817_,
		_w1799_,
		_w1840_,
		_w4367_,
		_w5617_
	);
	LUT3 #(
		.INIT('h70)
	) name5584 (
		_w1795_,
		_w1796_,
		_w4382_,
		_w5618_
	);
	LUT3 #(
		.INIT('h70)
	) name5585 (
		_w1863_,
		_w1875_,
		_w4033_,
		_w5619_
	);
	LUT3 #(
		.INIT('h01)
	) name5586 (
		_w5618_,
		_w5619_,
		_w5617_,
		_w5620_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5587 (
		_w2311_,
		_w2313_,
		_w4034_,
		_w5620_,
		_w5621_
	);
	LUT2 #(
		.INIT('h6)
	) name5588 (
		\a[14] ,
		_w5621_,
		_w5622_
	);
	LUT4 #(
		.INIT('h54ab)
	) name5589 (
		_w5398_,
		_w5456_,
		_w5457_,
		_w5459_,
		_w5623_
	);
	LUT2 #(
		.INIT('h4)
	) name5590 (
		_w5622_,
		_w5623_,
		_w5624_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5591 (
		_w1817_,
		_w1799_,
		_w1840_,
		_w4382_,
		_w5625_
	);
	LUT3 #(
		.INIT('h70)
	) name5592 (
		_w1898_,
		_w1928_,
		_w4033_,
		_w5626_
	);
	LUT3 #(
		.INIT('h70)
	) name5593 (
		_w1863_,
		_w1875_,
		_w4367_,
		_w5627_
	);
	LUT3 #(
		.INIT('h01)
	) name5594 (
		_w5626_,
		_w5627_,
		_w5625_,
		_w5628_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5595 (
		\a[14] ,
		_w3972_,
		_w4034_,
		_w5628_,
		_w5629_
	);
	LUT3 #(
		.INIT('h09)
	) name5596 (
		_w5456_,
		_w5458_,
		_w5629_,
		_w5630_
	);
	LUT3 #(
		.INIT('h1e)
	) name5597 (
		_w5412_,
		_w5453_,
		_w5455_,
		_w5631_
	);
	LUT3 #(
		.INIT('h70)
	) name5598 (
		_w1501_,
		_w1949_,
		_w4033_,
		_w5632_
	);
	LUT3 #(
		.INIT('h70)
	) name5599 (
		_w1898_,
		_w1928_,
		_w4367_,
		_w5633_
	);
	LUT3 #(
		.INIT('h70)
	) name5600 (
		_w1863_,
		_w1875_,
		_w4382_,
		_w5634_
	);
	LUT3 #(
		.INIT('h01)
	) name5601 (
		_w5633_,
		_w5634_,
		_w5632_,
		_w5635_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5602 (
		_w2307_,
		_w2309_,
		_w4034_,
		_w5635_,
		_w5636_
	);
	LUT2 #(
		.INIT('h6)
	) name5603 (
		\a[14] ,
		_w5636_,
		_w5637_
	);
	LUT2 #(
		.INIT('h2)
	) name5604 (
		_w5631_,
		_w5637_,
		_w5638_
	);
	LUT4 #(
		.INIT('h54ab)
	) name5605 (
		_w5420_,
		_w5449_,
		_w5450_,
		_w5452_,
		_w5639_
	);
	LUT3 #(
		.INIT('h70)
	) name5606 (
		_w1973_,
		_w1997_,
		_w4033_,
		_w5640_
	);
	LUT3 #(
		.INIT('h70)
	) name5607 (
		_w1898_,
		_w1928_,
		_w4382_,
		_w5641_
	);
	LUT3 #(
		.INIT('h70)
	) name5608 (
		_w1501_,
		_w1949_,
		_w4367_,
		_w5642_
	);
	LUT3 #(
		.INIT('h01)
	) name5609 (
		_w5641_,
		_w5642_,
		_w5640_,
		_w5643_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5610 (
		\a[14] ,
		_w4034_,
		_w4126_,
		_w5643_,
		_w5644_
	);
	LUT2 #(
		.INIT('h2)
	) name5611 (
		_w5639_,
		_w5644_,
		_w5645_
	);
	LUT2 #(
		.INIT('h9)
	) name5612 (
		_w5449_,
		_w5451_,
		_w5646_
	);
	LUT3 #(
		.INIT('h70)
	) name5613 (
		_w1973_,
		_w1997_,
		_w4367_,
		_w5647_
	);
	LUT3 #(
		.INIT('h70)
	) name5614 (
		_w1501_,
		_w1949_,
		_w4382_,
		_w5648_
	);
	LUT3 #(
		.INIT('h70)
	) name5615 (
		_w2023_,
		_w2055_,
		_w4033_,
		_w5649_
	);
	LUT3 #(
		.INIT('h01)
	) name5616 (
		_w5648_,
		_w5649_,
		_w5647_,
		_w5650_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5617 (
		_w2303_,
		_w2305_,
		_w4034_,
		_w5650_,
		_w5651_
	);
	LUT2 #(
		.INIT('h6)
	) name5618 (
		\a[14] ,
		_w5651_,
		_w5652_
	);
	LUT4 #(
		.INIT('h8241)
	) name5619 (
		\a[14] ,
		_w5449_,
		_w5451_,
		_w5651_,
		_w5653_
	);
	LUT3 #(
		.INIT('h70)
	) name5620 (
		_w1973_,
		_w1997_,
		_w4382_,
		_w5654_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5621 (
		_w1874_,
		_w2076_,
		_w2099_,
		_w4033_,
		_w5655_
	);
	LUT3 #(
		.INIT('h70)
	) name5622 (
		_w2023_,
		_w2055_,
		_w4367_,
		_w5656_
	);
	LUT3 #(
		.INIT('h01)
	) name5623 (
		_w5655_,
		_w5656_,
		_w5654_,
		_w5657_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5624 (
		\a[14] ,
		_w4034_,
		_w4151_,
		_w5657_,
		_w5658_
	);
	LUT2 #(
		.INIT('h9)
	) name5625 (
		_w5446_,
		_w5448_,
		_w5659_
	);
	LUT2 #(
		.INIT('h4)
	) name5626 (
		_w5658_,
		_w5659_,
		_w5660_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5627 (
		_w1874_,
		_w2076_,
		_w2099_,
		_w4367_,
		_w5661_
	);
	LUT3 #(
		.INIT('h70)
	) name5628 (
		_w2124_,
		_w2133_,
		_w4033_,
		_w5662_
	);
	LUT3 #(
		.INIT('h70)
	) name5629 (
		_w2023_,
		_w2055_,
		_w4382_,
		_w5663_
	);
	LUT3 #(
		.INIT('h01)
	) name5630 (
		_w5661_,
		_w5662_,
		_w5663_,
		_w5664_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5631 (
		_w2299_,
		_w2301_,
		_w4034_,
		_w5664_,
		_w5665_
	);
	LUT3 #(
		.INIT('h69)
	) name5632 (
		_w5193_,
		_w5440_,
		_w5445_,
		_w5666_
	);
	LUT3 #(
		.INIT('h90)
	) name5633 (
		\a[14] ,
		_w5665_,
		_w5666_,
		_w5667_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5634 (
		_w1874_,
		_w2076_,
		_w2099_,
		_w4382_,
		_w5668_
	);
	LUT3 #(
		.INIT('h70)
	) name5635 (
		_w2124_,
		_w2133_,
		_w4367_,
		_w5669_
	);
	LUT3 #(
		.INIT('h70)
	) name5636 (
		_w2155_,
		_w2156_,
		_w4033_,
		_w5670_
	);
	LUT3 #(
		.INIT('h01)
	) name5637 (
		_w5668_,
		_w5669_,
		_w5670_,
		_w5671_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5638 (
		\a[14] ,
		_w4034_,
		_w4209_,
		_w5671_,
		_w5672_
	);
	LUT3 #(
		.INIT('h8a)
	) name5639 (
		\a[17] ,
		_w5432_,
		_w5431_,
		_w5673_
	);
	LUT2 #(
		.INIT('h9)
	) name5640 (
		_w5439_,
		_w5673_,
		_w5674_
	);
	LUT2 #(
		.INIT('h4)
	) name5641 (
		_w5672_,
		_w5674_,
		_w5675_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5642 (
		_w2193_,
		_w2183_,
		_w2213_,
		_w4033_,
		_w5676_
	);
	LUT3 #(
		.INIT('h70)
	) name5643 (
		_w2155_,
		_w2156_,
		_w4367_,
		_w5677_
	);
	LUT3 #(
		.INIT('h70)
	) name5644 (
		_w2124_,
		_w2133_,
		_w4382_,
		_w5678_
	);
	LUT3 #(
		.INIT('h01)
	) name5645 (
		_w5676_,
		_w5677_,
		_w5678_,
		_w5679_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5646 (
		_w2295_,
		_w2297_,
		_w4034_,
		_w5679_,
		_w5680_
	);
	LUT4 #(
		.INIT('h002a)
	) name5647 (
		\a[17] ,
		_w2228_,
		_w2262_,
		_w3708_,
		_w5681_
	);
	LUT2 #(
		.INIT('h9)
	) name5648 (
		_w5431_,
		_w5681_,
		_w5682_
	);
	LUT3 #(
		.INIT('h90)
	) name5649 (
		\a[14] ,
		_w5680_,
		_w5682_,
		_w5683_
	);
	LUT3 #(
		.INIT('h70)
	) name5650 (
		_w2228_,
		_w2262_,
		_w4367_,
		_w5684_
	);
	LUT3 #(
		.INIT('h70)
	) name5651 (
		_w2273_,
		_w2293_,
		_w4382_,
		_w5685_
	);
	LUT4 #(
		.INIT('h000d)
	) name5652 (
		_w4034_,
		_w4599_,
		_w5684_,
		_w5685_,
		_w5686_
	);
	LUT3 #(
		.INIT('h07)
	) name5653 (
		_w2228_,
		_w2262_,
		_w4032_,
		_w5687_
	);
	LUT4 #(
		.INIT('haa80)
	) name5654 (
		\a[14] ,
		_w2228_,
		_w2262_,
		_w4032_,
		_w5688_
	);
	LUT3 #(
		.INIT('h84)
	) name5655 (
		_w2214_,
		_w4034_,
		_w4258_,
		_w5689_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5656 (
		_w2193_,
		_w2183_,
		_w2213_,
		_w4382_,
		_w5690_
	);
	LUT3 #(
		.INIT('h70)
	) name5657 (
		_w2228_,
		_w2262_,
		_w4033_,
		_w5691_
	);
	LUT3 #(
		.INIT('h70)
	) name5658 (
		_w2273_,
		_w2293_,
		_w4367_,
		_w5692_
	);
	LUT3 #(
		.INIT('h01)
	) name5659 (
		_w5691_,
		_w5692_,
		_w5690_,
		_w5693_
	);
	LUT2 #(
		.INIT('h4)
	) name5660 (
		_w5689_,
		_w5693_,
		_w5694_
	);
	LUT4 #(
		.INIT('h0800)
	) name5661 (
		_w5686_,
		_w5688_,
		_w5689_,
		_w5693_,
		_w5695_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5662 (
		_w2193_,
		_w2183_,
		_w2213_,
		_w4367_,
		_w5696_
	);
	LUT3 #(
		.INIT('h70)
	) name5663 (
		_w2155_,
		_w2156_,
		_w4382_,
		_w5697_
	);
	LUT3 #(
		.INIT('h70)
	) name5664 (
		_w2273_,
		_w2293_,
		_w4033_,
		_w5698_
	);
	LUT3 #(
		.INIT('h01)
	) name5665 (
		_w5696_,
		_w5697_,
		_w5698_,
		_w5699_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5666 (
		\a[14] ,
		_w4034_,
		_w4293_,
		_w5699_,
		_w5700_
	);
	LUT3 #(
		.INIT('h71)
	) name5667 (
		_w5432_,
		_w5695_,
		_w5700_,
		_w5701_
	);
	LUT3 #(
		.INIT('h06)
	) name5668 (
		\a[14] ,
		_w5680_,
		_w5682_,
		_w5702_
	);
	LUT3 #(
		.INIT('h69)
	) name5669 (
		\a[14] ,
		_w5680_,
		_w5682_,
		_w5703_
	);
	LUT3 #(
		.INIT('h54)
	) name5670 (
		_w5683_,
		_w5701_,
		_w5702_,
		_w5704_
	);
	LUT2 #(
		.INIT('h2)
	) name5671 (
		_w5672_,
		_w5674_,
		_w5705_
	);
	LUT2 #(
		.INIT('h9)
	) name5672 (
		_w5672_,
		_w5674_,
		_w5706_
	);
	LUT3 #(
		.INIT('h69)
	) name5673 (
		\a[14] ,
		_w5665_,
		_w5666_,
		_w5707_
	);
	LUT4 #(
		.INIT('h4d00)
	) name5674 (
		_w5672_,
		_w5674_,
		_w5704_,
		_w5707_,
		_w5708_
	);
	LUT2 #(
		.INIT('h2)
	) name5675 (
		_w5658_,
		_w5659_,
		_w5709_
	);
	LUT2 #(
		.INIT('h9)
	) name5676 (
		_w5658_,
		_w5659_,
		_w5710_
	);
	LUT4 #(
		.INIT('h5501)
	) name5677 (
		_w5660_,
		_w5667_,
		_w5708_,
		_w5709_,
		_w5711_
	);
	LUT4 #(
		.INIT('h1428)
	) name5678 (
		\a[14] ,
		_w5449_,
		_w5451_,
		_w5651_,
		_w5712_
	);
	LUT4 #(
		.INIT('h6996)
	) name5679 (
		\a[14] ,
		_w5449_,
		_w5451_,
		_w5651_,
		_w5713_
	);
	LUT2 #(
		.INIT('h9)
	) name5680 (
		_w5639_,
		_w5644_,
		_w5714_
	);
	LUT4 #(
		.INIT('h2b00)
	) name5681 (
		_w5646_,
		_w5652_,
		_w5711_,
		_w5714_,
		_w5715_
	);
	LUT2 #(
		.INIT('h4)
	) name5682 (
		_w5631_,
		_w5637_,
		_w5716_
	);
	LUT2 #(
		.INIT('h9)
	) name5683 (
		_w5631_,
		_w5637_,
		_w5717_
	);
	LUT4 #(
		.INIT('h5501)
	) name5684 (
		_w5638_,
		_w5645_,
		_w5715_,
		_w5716_,
		_w5718_
	);
	LUT3 #(
		.INIT('h60)
	) name5685 (
		_w5456_,
		_w5458_,
		_w5629_,
		_w5719_
	);
	LUT3 #(
		.INIT('h96)
	) name5686 (
		_w5456_,
		_w5458_,
		_w5629_,
		_w5720_
	);
	LUT2 #(
		.INIT('h9)
	) name5687 (
		_w5622_,
		_w5623_,
		_w5721_
	);
	LUT4 #(
		.INIT('hba00)
	) name5688 (
		_w5630_,
		_w5718_,
		_w5720_,
		_w5721_,
		_w5722_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name5689 (
		_w5390_,
		_w5460_,
		_w5462_,
		_w5615_,
		_w5723_
	);
	LUT4 #(
		.INIT('h0155)
	) name5690 (
		_w5616_,
		_w5624_,
		_w5722_,
		_w5723_,
		_w5724_
	);
	LUT3 #(
		.INIT('h60)
	) name5691 (
		_w5463_,
		_w5465_,
		_w5609_,
		_w5725_
	);
	LUT3 #(
		.INIT('h96)
	) name5692 (
		_w5463_,
		_w5465_,
		_w5609_,
		_w5726_
	);
	LUT2 #(
		.INIT('h9)
	) name5693 (
		_w5596_,
		_w5601_,
		_w5727_
	);
	LUT4 #(
		.INIT('h2b00)
	) name5694 (
		_w5603_,
		_w5609_,
		_w5724_,
		_w5727_,
		_w5728_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name5695 (
		_w5369_,
		_w5467_,
		_w5468_,
		_w5594_,
		_w5729_
	);
	LUT4 #(
		.INIT('h0155)
	) name5696 (
		_w5595_,
		_w5602_,
		_w5728_,
		_w5729_,
		_w5730_
	);
	LUT3 #(
		.INIT('h60)
	) name5697 (
		_w5469_,
		_w5471_,
		_w5587_,
		_w5731_
	);
	LUT3 #(
		.INIT('h96)
	) name5698 (
		_w5469_,
		_w5471_,
		_w5587_,
		_w5732_
	);
	LUT2 #(
		.INIT('h9)
	) name5699 (
		_w5580_,
		_w5581_,
		_w5733_
	);
	LUT4 #(
		.INIT('hba00)
	) name5700 (
		_w5588_,
		_w5730_,
		_w5732_,
		_w5733_,
		_w5734_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name5701 (
		_w5347_,
		_w5473_,
		_w5474_,
		_w5573_,
		_w5735_
	);
	LUT4 #(
		.INIT('h0155)
	) name5702 (
		_w5574_,
		_w5582_,
		_w5734_,
		_w5735_,
		_w5736_
	);
	LUT3 #(
		.INIT('h60)
	) name5703 (
		_w5475_,
		_w5477_,
		_w5567_,
		_w5737_
	);
	LUT3 #(
		.INIT('h96)
	) name5704 (
		_w5475_,
		_w5477_,
		_w5567_,
		_w5738_
	);
	LUT2 #(
		.INIT('h9)
	) name5705 (
		_w5554_,
		_w5559_,
		_w5739_
	);
	LUT4 #(
		.INIT('h2b00)
	) name5706 (
		_w5561_,
		_w5567_,
		_w5736_,
		_w5739_,
		_w5740_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name5707 (
		_w5327_,
		_w5479_,
		_w5480_,
		_w5552_,
		_w5741_
	);
	LUT4 #(
		.INIT('h0155)
	) name5708 (
		_w5553_,
		_w5560_,
		_w5740_,
		_w5741_,
		_w5742_
	);
	LUT3 #(
		.INIT('h60)
	) name5709 (
		_w5481_,
		_w5483_,
		_w5545_,
		_w5743_
	);
	LUT3 #(
		.INIT('h96)
	) name5710 (
		_w5481_,
		_w5483_,
		_w5545_,
		_w5744_
	);
	LUT2 #(
		.INIT('h9)
	) name5711 (
		_w5533_,
		_w5539_,
		_w5745_
	);
	LUT4 #(
		.INIT('hba00)
	) name5712 (
		_w5546_,
		_w5742_,
		_w5744_,
		_w5745_,
		_w5746_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name5713 (
		_w5305_,
		_w5485_,
		_w5486_,
		_w5531_,
		_w5747_
	);
	LUT4 #(
		.INIT('h0155)
	) name5714 (
		_w5532_,
		_w5540_,
		_w5746_,
		_w5747_,
		_w5748_
	);
	LUT3 #(
		.INIT('h96)
	) name5715 (
		_w5487_,
		_w5488_,
		_w5494_,
		_w5749_
	);
	LUT3 #(
		.INIT('h70)
	) name5716 (
		_w725_,
		_w764_,
		_w4700_,
		_w5750_
	);
	LUT3 #(
		.INIT('h70)
	) name5717 (
		_w801_,
		_w851_,
		_w4684_,
		_w5751_
	);
	LUT3 #(
		.INIT('h70)
	) name5718 (
		_w871_,
		_w927_,
		_w4458_,
		_w5752_
	);
	LUT3 #(
		.INIT('h01)
	) name5719 (
		_w5751_,
		_w5752_,
		_w5750_,
		_w5753_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5720 (
		\a[11] ,
		_w2724_,
		_w4459_,
		_w5753_,
		_w5754_
	);
	LUT3 #(
		.INIT('hb2)
	) name5721 (
		_w5748_,
		_w5749_,
		_w5754_,
		_w5755_
	);
	LUT4 #(
		.INIT('hb24d)
	) name5722 (
		_w5487_,
		_w5488_,
		_w5494_,
		_w5497_,
		_w5756_
	);
	LUT2 #(
		.INIT('h6)
	) name5723 (
		_w5505_,
		_w5756_,
		_w5757_
	);
	LUT4 #(
		.INIT('h004d)
	) name5724 (
		_w5748_,
		_w5749_,
		_w5754_,
		_w5757_,
		_w5758_
	);
	LUT4 #(
		.INIT('hb200)
	) name5725 (
		_w5748_,
		_w5749_,
		_w5754_,
		_w5757_,
		_w5759_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5726 (
		_w486_,
		_w487_,
		_w509_,
		_w5286_,
		_w5760_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5727 (
		_w587_,
		_w608_,
		_w624_,
		_w4875_,
		_w5761_
	);
	LUT3 #(
		.INIT('h70)
	) name5728 (
		_w544_,
		_w558_,
		_w5271_,
		_w5762_
	);
	LUT3 #(
		.INIT('h01)
	) name5729 (
		_w5760_,
		_w5761_,
		_w5762_,
		_w5763_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5730 (
		\a[8] ,
		_w2526_,
		_w4876_,
		_w5763_,
		_w5764_
	);
	LUT3 #(
		.INIT('h54)
	) name5731 (
		_w5758_,
		_w5759_,
		_w5764_,
		_w5765_
	);
	LUT4 #(
		.INIT('h0115)
	) name5732 (
		_w5526_,
		_w5755_,
		_w5757_,
		_w5764_,
		_w5766_
	);
	LUT4 #(
		.INIT('ha880)
	) name5733 (
		_w5526_,
		_w5755_,
		_w5757_,
		_w5764_,
		_w5767_
	);
	LUT4 #(
		.INIT('h6665)
	) name5734 (
		_w5291_,
		_w5498_,
		_w5499_,
		_w5505_,
		_w5768_
	);
	LUT2 #(
		.INIT('h9)
	) name5735 (
		_w5514_,
		_w5768_,
		_w5769_
	);
	LUT4 #(
		.INIT('h2a02)
	) name5736 (
		_w5522_,
		_w5526_,
		_w5765_,
		_w5769_,
		_w5770_
	);
	LUT3 #(
		.INIT('h70)
	) name5737 (
		_w763_,
		_w983_,
		_w4458_,
		_w5771_
	);
	LUT3 #(
		.INIT('h70)
	) name5738 (
		_w871_,
		_w927_,
		_w4684_,
		_w5772_
	);
	LUT3 #(
		.INIT('h70)
	) name5739 (
		_w801_,
		_w851_,
		_w4700_,
		_w5773_
	);
	LUT3 #(
		.INIT('h01)
	) name5740 (
		_w5772_,
		_w5773_,
		_w5771_,
		_w5774_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5741 (
		_w2343_,
		_w2345_,
		_w4459_,
		_w5774_,
		_w5775_
	);
	LUT2 #(
		.INIT('h6)
	) name5742 (
		\a[11] ,
		_w5775_,
		_w5776_
	);
	LUT4 #(
		.INIT('h001e)
	) name5743 (
		_w5540_,
		_w5746_,
		_w5747_,
		_w5776_,
		_w5777_
	);
	LUT3 #(
		.INIT('h70)
	) name5744 (
		_w1009_,
		_w1050_,
		_w4458_,
		_w5778_
	);
	LUT3 #(
		.INIT('h70)
	) name5745 (
		_w871_,
		_w927_,
		_w4700_,
		_w5779_
	);
	LUT3 #(
		.INIT('h70)
	) name5746 (
		_w763_,
		_w983_,
		_w4684_,
		_w5780_
	);
	LUT3 #(
		.INIT('h01)
	) name5747 (
		_w5779_,
		_w5780_,
		_w5778_,
		_w5781_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5748 (
		\a[11] ,
		_w2839_,
		_w4459_,
		_w5781_,
		_w5782_
	);
	LUT4 #(
		.INIT('h54ab)
	) name5749 (
		_w5546_,
		_w5742_,
		_w5743_,
		_w5745_,
		_w5783_
	);
	LUT2 #(
		.INIT('h4)
	) name5750 (
		_w5782_,
		_w5783_,
		_w5784_
	);
	LUT3 #(
		.INIT('h70)
	) name5751 (
		_w1071_,
		_w1102_,
		_w4458_,
		_w5785_
	);
	LUT3 #(
		.INIT('h70)
	) name5752 (
		_w763_,
		_w983_,
		_w4700_,
		_w5786_
	);
	LUT3 #(
		.INIT('h70)
	) name5753 (
		_w1009_,
		_w1050_,
		_w4684_,
		_w5787_
	);
	LUT3 #(
		.INIT('h01)
	) name5754 (
		_w5786_,
		_w5787_,
		_w5785_,
		_w5788_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5755 (
		_w2339_,
		_w2341_,
		_w4459_,
		_w5788_,
		_w5789_
	);
	LUT2 #(
		.INIT('h6)
	) name5756 (
		\a[11] ,
		_w5789_,
		_w5790_
	);
	LUT2 #(
		.INIT('h9)
	) name5757 (
		_w5742_,
		_w5744_,
		_w5791_
	);
	LUT3 #(
		.INIT('h09)
	) name5758 (
		_w5742_,
		_w5744_,
		_w5790_,
		_w5792_
	);
	LUT3 #(
		.INIT('h70)
	) name5759 (
		_w1136_,
		_w1187_,
		_w4458_,
		_w5793_
	);
	LUT3 #(
		.INIT('h70)
	) name5760 (
		_w1009_,
		_w1050_,
		_w4700_,
		_w5794_
	);
	LUT3 #(
		.INIT('h70)
	) name5761 (
		_w1071_,
		_w1102_,
		_w4684_,
		_w5795_
	);
	LUT3 #(
		.INIT('h01)
	) name5762 (
		_w5794_,
		_w5795_,
		_w5793_,
		_w5796_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5763 (
		\a[11] ,
		_w2936_,
		_w4459_,
		_w5796_,
		_w5797_
	);
	LUT4 #(
		.INIT('h001e)
	) name5764 (
		_w5560_,
		_w5740_,
		_w5741_,
		_w5797_,
		_w5798_
	);
	LUT3 #(
		.INIT('h70)
	) name5765 (
		_w1136_,
		_w1187_,
		_w4684_,
		_w5799_
	);
	LUT3 #(
		.INIT('h70)
	) name5766 (
		_w1071_,
		_w1102_,
		_w4700_,
		_w5800_
	);
	LUT3 #(
		.INIT('h70)
	) name5767 (
		_w1202_,
		_w1233_,
		_w4458_,
		_w5801_
	);
	LUT3 #(
		.INIT('h01)
	) name5768 (
		_w5800_,
		_w5801_,
		_w5799_,
		_w5802_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5769 (
		_w2335_,
		_w2337_,
		_w4459_,
		_w5802_,
		_w5803_
	);
	LUT2 #(
		.INIT('h6)
	) name5770 (
		\a[11] ,
		_w5803_,
		_w5804_
	);
	LUT4 #(
		.INIT('h54ab)
	) name5771 (
		_w5568_,
		_w5736_,
		_w5737_,
		_w5739_,
		_w5805_
	);
	LUT2 #(
		.INIT('h4)
	) name5772 (
		_w5804_,
		_w5805_,
		_w5806_
	);
	LUT3 #(
		.INIT('h70)
	) name5773 (
		_w1202_,
		_w1233_,
		_w4684_,
		_w5807_
	);
	LUT3 #(
		.INIT('h70)
	) name5774 (
		_w1253_,
		_w1294_,
		_w4458_,
		_w5808_
	);
	LUT3 #(
		.INIT('h70)
	) name5775 (
		_w1136_,
		_w1187_,
		_w4700_,
		_w5809_
	);
	LUT3 #(
		.INIT('h01)
	) name5776 (
		_w5808_,
		_w5809_,
		_w5807_,
		_w5810_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5777 (
		\a[11] ,
		_w3067_,
		_w4459_,
		_w5810_,
		_w5811_
	);
	LUT3 #(
		.INIT('h09)
	) name5778 (
		_w5736_,
		_w5738_,
		_w5811_,
		_w5812_
	);
	LUT3 #(
		.INIT('h70)
	) name5779 (
		_w1202_,
		_w1233_,
		_w4700_,
		_w5813_
	);
	LUT3 #(
		.INIT('h70)
	) name5780 (
		_w1325_,
		_w1367_,
		_w4458_,
		_w5814_
	);
	LUT3 #(
		.INIT('h70)
	) name5781 (
		_w1253_,
		_w1294_,
		_w4684_,
		_w5815_
	);
	LUT3 #(
		.INIT('h01)
	) name5782 (
		_w5814_,
		_w5815_,
		_w5813_,
		_w5816_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5783 (
		_w2331_,
		_w2333_,
		_w4459_,
		_w5816_,
		_w5817_
	);
	LUT2 #(
		.INIT('h6)
	) name5784 (
		\a[11] ,
		_w5817_,
		_w5818_
	);
	LUT4 #(
		.INIT('h001e)
	) name5785 (
		_w5582_,
		_w5734_,
		_w5735_,
		_w5818_,
		_w5819_
	);
	LUT4 #(
		.INIT('h54ab)
	) name5786 (
		_w5588_,
		_w5730_,
		_w5731_,
		_w5733_,
		_w5820_
	);
	LUT3 #(
		.INIT('h70)
	) name5787 (
		_w1381_,
		_w1398_,
		_w4458_,
		_w5821_
	);
	LUT3 #(
		.INIT('h70)
	) name5788 (
		_w1325_,
		_w1367_,
		_w4684_,
		_w5822_
	);
	LUT3 #(
		.INIT('h70)
	) name5789 (
		_w1253_,
		_w1294_,
		_w4700_,
		_w5823_
	);
	LUT3 #(
		.INIT('h01)
	) name5790 (
		_w5822_,
		_w5823_,
		_w5821_,
		_w5824_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5791 (
		\a[11] ,
		_w3182_,
		_w4459_,
		_w5824_,
		_w5825_
	);
	LUT2 #(
		.INIT('h2)
	) name5792 (
		_w5820_,
		_w5825_,
		_w5826_
	);
	LUT2 #(
		.INIT('h9)
	) name5793 (
		_w5730_,
		_w5732_,
		_w5827_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5794 (
		_w1454_,
		_w1426_,
		_w1478_,
		_w4458_,
		_w5828_
	);
	LUT3 #(
		.INIT('h70)
	) name5795 (
		_w1325_,
		_w1367_,
		_w4700_,
		_w5829_
	);
	LUT3 #(
		.INIT('h70)
	) name5796 (
		_w1381_,
		_w1398_,
		_w4684_,
		_w5830_
	);
	LUT3 #(
		.INIT('h01)
	) name5797 (
		_w5829_,
		_w5830_,
		_w5828_,
		_w5831_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5798 (
		_w2327_,
		_w2329_,
		_w4459_,
		_w5831_,
		_w5832_
	);
	LUT2 #(
		.INIT('h6)
	) name5799 (
		\a[11] ,
		_w5832_,
		_w5833_
	);
	LUT3 #(
		.INIT('h09)
	) name5800 (
		_w5730_,
		_w5732_,
		_w5833_,
		_w5834_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5801 (
		_w1454_,
		_w1426_,
		_w1478_,
		_w4684_,
		_w5835_
	);
	LUT3 #(
		.INIT('h70)
	) name5802 (
		_w1381_,
		_w1398_,
		_w4700_,
		_w5836_
	);
	LUT3 #(
		.INIT('h70)
	) name5803 (
		_w1501_,
		_w1545_,
		_w4458_,
		_w5837_
	);
	LUT3 #(
		.INIT('h01)
	) name5804 (
		_w5836_,
		_w5837_,
		_w5835_,
		_w5838_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5805 (
		\a[11] ,
		_w3362_,
		_w4459_,
		_w5838_,
		_w5839_
	);
	LUT4 #(
		.INIT('h001e)
	) name5806 (
		_w5602_,
		_w5728_,
		_w5729_,
		_w5839_,
		_w5840_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5807 (
		_w1454_,
		_w1426_,
		_w1478_,
		_w4700_,
		_w5841_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5808 (
		_w1584_,
		_w1569_,
		_w1606_,
		_w4458_,
		_w5842_
	);
	LUT3 #(
		.INIT('h70)
	) name5809 (
		_w1501_,
		_w1545_,
		_w4684_,
		_w5843_
	);
	LUT3 #(
		.INIT('h01)
	) name5810 (
		_w5842_,
		_w5843_,
		_w5841_,
		_w5844_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5811 (
		_w2323_,
		_w2325_,
		_w4459_,
		_w5844_,
		_w5845_
	);
	LUT2 #(
		.INIT('h6)
	) name5812 (
		\a[11] ,
		_w5845_,
		_w5846_
	);
	LUT4 #(
		.INIT('h54ab)
	) name5813 (
		_w5610_,
		_w5724_,
		_w5725_,
		_w5727_,
		_w5847_
	);
	LUT2 #(
		.INIT('h4)
	) name5814 (
		_w5846_,
		_w5847_,
		_w5848_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5815 (
		_w1584_,
		_w1569_,
		_w1606_,
		_w4684_,
		_w5849_
	);
	LUT3 #(
		.INIT('h70)
	) name5816 (
		_w1501_,
		_w1545_,
		_w4700_,
		_w5850_
	);
	LUT3 #(
		.INIT('h70)
	) name5817 (
		_w1620_,
		_w1661_,
		_w4458_,
		_w5851_
	);
	LUT3 #(
		.INIT('h01)
	) name5818 (
		_w5849_,
		_w5850_,
		_w5851_,
		_w5852_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5819 (
		\a[11] ,
		_w3495_,
		_w4459_,
		_w5852_,
		_w5853_
	);
	LUT3 #(
		.INIT('h09)
	) name5820 (
		_w5724_,
		_w5726_,
		_w5853_,
		_w5854_
	);
	LUT3 #(
		.INIT('h70)
	) name5821 (
		_w1692_,
		_w1723_,
		_w4458_,
		_w5855_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5822 (
		_w1584_,
		_w1569_,
		_w1606_,
		_w4700_,
		_w5856_
	);
	LUT3 #(
		.INIT('h70)
	) name5823 (
		_w1620_,
		_w1661_,
		_w4684_,
		_w5857_
	);
	LUT3 #(
		.INIT('h01)
	) name5824 (
		_w5856_,
		_w5857_,
		_w5855_,
		_w5858_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5825 (
		_w2319_,
		_w2321_,
		_w4459_,
		_w5858_,
		_w5859_
	);
	LUT2 #(
		.INIT('h6)
	) name5826 (
		\a[11] ,
		_w5859_,
		_w5860_
	);
	LUT4 #(
		.INIT('h001e)
	) name5827 (
		_w5624_,
		_w5722_,
		_w5723_,
		_w5860_,
		_w5861_
	);
	LUT4 #(
		.INIT('h54ab)
	) name5828 (
		_w5630_,
		_w5718_,
		_w5719_,
		_w5721_,
		_w5862_
	);
	LUT3 #(
		.INIT('h70)
	) name5829 (
		_w1692_,
		_w1723_,
		_w4684_,
		_w5863_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5830 (
		_w1751_,
		_w1742_,
		_w1771_,
		_w4458_,
		_w5864_
	);
	LUT3 #(
		.INIT('h70)
	) name5831 (
		_w1620_,
		_w1661_,
		_w4700_,
		_w5865_
	);
	LUT3 #(
		.INIT('h01)
	) name5832 (
		_w5864_,
		_w5865_,
		_w5863_,
		_w5866_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5833 (
		\a[11] ,
		_w3599_,
		_w4459_,
		_w5866_,
		_w5867_
	);
	LUT2 #(
		.INIT('h2)
	) name5834 (
		_w5862_,
		_w5867_,
		_w5868_
	);
	LUT2 #(
		.INIT('h9)
	) name5835 (
		_w5718_,
		_w5720_,
		_w5869_
	);
	LUT3 #(
		.INIT('h70)
	) name5836 (
		_w1692_,
		_w1723_,
		_w4700_,
		_w5870_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5837 (
		_w1751_,
		_w1742_,
		_w1771_,
		_w4684_,
		_w5871_
	);
	LUT3 #(
		.INIT('h70)
	) name5838 (
		_w1795_,
		_w1796_,
		_w4458_,
		_w5872_
	);
	LUT3 #(
		.INIT('h01)
	) name5839 (
		_w5871_,
		_w5872_,
		_w5870_,
		_w5873_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5840 (
		_w2315_,
		_w2317_,
		_w4459_,
		_w5873_,
		_w5874_
	);
	LUT2 #(
		.INIT('h6)
	) name5841 (
		\a[11] ,
		_w5874_,
		_w5875_
	);
	LUT3 #(
		.INIT('h09)
	) name5842 (
		_w5718_,
		_w5720_,
		_w5875_,
		_w5876_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5843 (
		_w1751_,
		_w1742_,
		_w1771_,
		_w4700_,
		_w5877_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5844 (
		_w1817_,
		_w1799_,
		_w1840_,
		_w4458_,
		_w5878_
	);
	LUT3 #(
		.INIT('h70)
	) name5845 (
		_w1795_,
		_w1796_,
		_w4684_,
		_w5879_
	);
	LUT3 #(
		.INIT('h01)
	) name5846 (
		_w5878_,
		_w5879_,
		_w5877_,
		_w5880_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5847 (
		\a[11] ,
		_w3909_,
		_w4459_,
		_w5880_,
		_w5881_
	);
	LUT4 #(
		.INIT('h001e)
	) name5848 (
		_w5645_,
		_w5715_,
		_w5717_,
		_w5881_,
		_w5882_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5849 (
		_w1817_,
		_w1799_,
		_w1840_,
		_w4684_,
		_w5883_
	);
	LUT3 #(
		.INIT('h70)
	) name5850 (
		_w1795_,
		_w1796_,
		_w4700_,
		_w5884_
	);
	LUT3 #(
		.INIT('h70)
	) name5851 (
		_w1863_,
		_w1875_,
		_w4458_,
		_w5885_
	);
	LUT3 #(
		.INIT('h01)
	) name5852 (
		_w5884_,
		_w5885_,
		_w5883_,
		_w5886_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5853 (
		_w2311_,
		_w2313_,
		_w4459_,
		_w5886_,
		_w5887_
	);
	LUT2 #(
		.INIT('h6)
	) name5854 (
		\a[11] ,
		_w5887_,
		_w5888_
	);
	LUT4 #(
		.INIT('h54ab)
	) name5855 (
		_w5653_,
		_w5711_,
		_w5712_,
		_w5714_,
		_w5889_
	);
	LUT2 #(
		.INIT('h4)
	) name5856 (
		_w5888_,
		_w5889_,
		_w5890_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5857 (
		_w1817_,
		_w1799_,
		_w1840_,
		_w4700_,
		_w5891_
	);
	LUT3 #(
		.INIT('h70)
	) name5858 (
		_w1898_,
		_w1928_,
		_w4458_,
		_w5892_
	);
	LUT3 #(
		.INIT('h70)
	) name5859 (
		_w1863_,
		_w1875_,
		_w4684_,
		_w5893_
	);
	LUT3 #(
		.INIT('h01)
	) name5860 (
		_w5892_,
		_w5893_,
		_w5891_,
		_w5894_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5861 (
		\a[11] ,
		_w3972_,
		_w4459_,
		_w5894_,
		_w5895_
	);
	LUT3 #(
		.INIT('h09)
	) name5862 (
		_w5711_,
		_w5713_,
		_w5895_,
		_w5896_
	);
	LUT3 #(
		.INIT('h1e)
	) name5863 (
		_w5667_,
		_w5708_,
		_w5710_,
		_w5897_
	);
	LUT3 #(
		.INIT('h70)
	) name5864 (
		_w1501_,
		_w1949_,
		_w4458_,
		_w5898_
	);
	LUT3 #(
		.INIT('h70)
	) name5865 (
		_w1898_,
		_w1928_,
		_w4684_,
		_w5899_
	);
	LUT3 #(
		.INIT('h70)
	) name5866 (
		_w1863_,
		_w1875_,
		_w4700_,
		_w5900_
	);
	LUT3 #(
		.INIT('h01)
	) name5867 (
		_w5899_,
		_w5900_,
		_w5898_,
		_w5901_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5868 (
		_w2307_,
		_w2309_,
		_w4459_,
		_w5901_,
		_w5902_
	);
	LUT2 #(
		.INIT('h6)
	) name5869 (
		\a[11] ,
		_w5902_,
		_w5903_
	);
	LUT2 #(
		.INIT('h2)
	) name5870 (
		_w5897_,
		_w5903_,
		_w5904_
	);
	LUT4 #(
		.INIT('h54ab)
	) name5871 (
		_w5675_,
		_w5704_,
		_w5705_,
		_w5707_,
		_w5905_
	);
	LUT3 #(
		.INIT('h70)
	) name5872 (
		_w1973_,
		_w1997_,
		_w4458_,
		_w5906_
	);
	LUT3 #(
		.INIT('h70)
	) name5873 (
		_w1898_,
		_w1928_,
		_w4700_,
		_w5907_
	);
	LUT3 #(
		.INIT('h70)
	) name5874 (
		_w1501_,
		_w1949_,
		_w4684_,
		_w5908_
	);
	LUT3 #(
		.INIT('h01)
	) name5875 (
		_w5907_,
		_w5908_,
		_w5906_,
		_w5909_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5876 (
		\a[11] ,
		_w4126_,
		_w4459_,
		_w5909_,
		_w5910_
	);
	LUT2 #(
		.INIT('h2)
	) name5877 (
		_w5905_,
		_w5910_,
		_w5911_
	);
	LUT2 #(
		.INIT('h9)
	) name5878 (
		_w5704_,
		_w5706_,
		_w5912_
	);
	LUT3 #(
		.INIT('h70)
	) name5879 (
		_w1973_,
		_w1997_,
		_w4684_,
		_w5913_
	);
	LUT3 #(
		.INIT('h70)
	) name5880 (
		_w1501_,
		_w1949_,
		_w4700_,
		_w5914_
	);
	LUT3 #(
		.INIT('h70)
	) name5881 (
		_w2023_,
		_w2055_,
		_w4458_,
		_w5915_
	);
	LUT3 #(
		.INIT('h01)
	) name5882 (
		_w5914_,
		_w5915_,
		_w5913_,
		_w5916_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5883 (
		_w2303_,
		_w2305_,
		_w4459_,
		_w5916_,
		_w5917_
	);
	LUT2 #(
		.INIT('h6)
	) name5884 (
		\a[11] ,
		_w5917_,
		_w5918_
	);
	LUT4 #(
		.INIT('h8241)
	) name5885 (
		\a[11] ,
		_w5704_,
		_w5706_,
		_w5917_,
		_w5919_
	);
	LUT3 #(
		.INIT('h70)
	) name5886 (
		_w1973_,
		_w1997_,
		_w4700_,
		_w5920_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5887 (
		_w1874_,
		_w2076_,
		_w2099_,
		_w4458_,
		_w5921_
	);
	LUT3 #(
		.INIT('h70)
	) name5888 (
		_w2023_,
		_w2055_,
		_w4684_,
		_w5922_
	);
	LUT3 #(
		.INIT('h01)
	) name5889 (
		_w5921_,
		_w5922_,
		_w5920_,
		_w5923_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5890 (
		\a[11] ,
		_w4151_,
		_w4459_,
		_w5923_,
		_w5924_
	);
	LUT2 #(
		.INIT('h9)
	) name5891 (
		_w5701_,
		_w5703_,
		_w5925_
	);
	LUT2 #(
		.INIT('h4)
	) name5892 (
		_w5924_,
		_w5925_,
		_w5926_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5893 (
		_w1874_,
		_w2076_,
		_w2099_,
		_w4684_,
		_w5927_
	);
	LUT3 #(
		.INIT('h70)
	) name5894 (
		_w2124_,
		_w2133_,
		_w4458_,
		_w5928_
	);
	LUT3 #(
		.INIT('h70)
	) name5895 (
		_w2023_,
		_w2055_,
		_w4700_,
		_w5929_
	);
	LUT3 #(
		.INIT('h01)
	) name5896 (
		_w5927_,
		_w5928_,
		_w5929_,
		_w5930_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5897 (
		_w2299_,
		_w2301_,
		_w4459_,
		_w5930_,
		_w5931_
	);
	LUT3 #(
		.INIT('h69)
	) name5898 (
		_w5432_,
		_w5695_,
		_w5700_,
		_w5932_
	);
	LUT3 #(
		.INIT('h90)
	) name5899 (
		\a[11] ,
		_w5931_,
		_w5932_,
		_w5933_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5900 (
		_w1874_,
		_w2076_,
		_w2099_,
		_w4700_,
		_w5934_
	);
	LUT3 #(
		.INIT('h70)
	) name5901 (
		_w2124_,
		_w2133_,
		_w4684_,
		_w5935_
	);
	LUT3 #(
		.INIT('h70)
	) name5902 (
		_w2155_,
		_w2156_,
		_w4458_,
		_w5936_
	);
	LUT3 #(
		.INIT('h01)
	) name5903 (
		_w5934_,
		_w5935_,
		_w5936_,
		_w5937_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5904 (
		\a[11] ,
		_w4209_,
		_w4459_,
		_w5937_,
		_w5938_
	);
	LUT3 #(
		.INIT('h8a)
	) name5905 (
		\a[14] ,
		_w5687_,
		_w5686_,
		_w5939_
	);
	LUT2 #(
		.INIT('h9)
	) name5906 (
		_w5694_,
		_w5939_,
		_w5940_
	);
	LUT2 #(
		.INIT('h4)
	) name5907 (
		_w5938_,
		_w5940_,
		_w5941_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5908 (
		_w2193_,
		_w2183_,
		_w2213_,
		_w4458_,
		_w5942_
	);
	LUT3 #(
		.INIT('h70)
	) name5909 (
		_w2155_,
		_w2156_,
		_w4684_,
		_w5943_
	);
	LUT3 #(
		.INIT('h70)
	) name5910 (
		_w2124_,
		_w2133_,
		_w4700_,
		_w5944_
	);
	LUT3 #(
		.INIT('h01)
	) name5911 (
		_w5942_,
		_w5943_,
		_w5944_,
		_w5945_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5912 (
		_w2295_,
		_w2297_,
		_w4459_,
		_w5945_,
		_w5946_
	);
	LUT4 #(
		.INIT('h002a)
	) name5913 (
		\a[14] ,
		_w2228_,
		_w2262_,
		_w4032_,
		_w5947_
	);
	LUT2 #(
		.INIT('h9)
	) name5914 (
		_w5686_,
		_w5947_,
		_w5948_
	);
	LUT3 #(
		.INIT('h90)
	) name5915 (
		\a[11] ,
		_w5946_,
		_w5948_,
		_w5949_
	);
	LUT3 #(
		.INIT('h70)
	) name5916 (
		_w2228_,
		_w2262_,
		_w4684_,
		_w5950_
	);
	LUT3 #(
		.INIT('h70)
	) name5917 (
		_w2273_,
		_w2293_,
		_w4700_,
		_w5951_
	);
	LUT4 #(
		.INIT('h000d)
	) name5918 (
		_w4459_,
		_w4599_,
		_w5950_,
		_w5951_,
		_w5952_
	);
	LUT3 #(
		.INIT('h07)
	) name5919 (
		_w2228_,
		_w2262_,
		_w4457_,
		_w5953_
	);
	LUT4 #(
		.INIT('haa80)
	) name5920 (
		\a[11] ,
		_w2228_,
		_w2262_,
		_w4457_,
		_w5954_
	);
	LUT3 #(
		.INIT('h90)
	) name5921 (
		_w2214_,
		_w4258_,
		_w4459_,
		_w5955_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5922 (
		_w2193_,
		_w2183_,
		_w2213_,
		_w4700_,
		_w5956_
	);
	LUT3 #(
		.INIT('h70)
	) name5923 (
		_w2228_,
		_w2262_,
		_w4458_,
		_w5957_
	);
	LUT3 #(
		.INIT('h70)
	) name5924 (
		_w2273_,
		_w2293_,
		_w4684_,
		_w5958_
	);
	LUT3 #(
		.INIT('h01)
	) name5925 (
		_w5957_,
		_w5958_,
		_w5956_,
		_w5959_
	);
	LUT2 #(
		.INIT('h4)
	) name5926 (
		_w5955_,
		_w5959_,
		_w5960_
	);
	LUT4 #(
		.INIT('h0800)
	) name5927 (
		_w5952_,
		_w5954_,
		_w5955_,
		_w5959_,
		_w5961_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5928 (
		_w2193_,
		_w2183_,
		_w2213_,
		_w4684_,
		_w5962_
	);
	LUT3 #(
		.INIT('h70)
	) name5929 (
		_w2155_,
		_w2156_,
		_w4700_,
		_w5963_
	);
	LUT3 #(
		.INIT('h70)
	) name5930 (
		_w2273_,
		_w2293_,
		_w4458_,
		_w5964_
	);
	LUT3 #(
		.INIT('h01)
	) name5931 (
		_w5962_,
		_w5963_,
		_w5964_,
		_w5965_
	);
	LUT4 #(
		.INIT('h95aa)
	) name5932 (
		\a[11] ,
		_w4293_,
		_w4459_,
		_w5965_,
		_w5966_
	);
	LUT3 #(
		.INIT('h71)
	) name5933 (
		_w5687_,
		_w5961_,
		_w5966_,
		_w5967_
	);
	LUT3 #(
		.INIT('h06)
	) name5934 (
		\a[11] ,
		_w5946_,
		_w5948_,
		_w5968_
	);
	LUT3 #(
		.INIT('h69)
	) name5935 (
		\a[11] ,
		_w5946_,
		_w5948_,
		_w5969_
	);
	LUT3 #(
		.INIT('h54)
	) name5936 (
		_w5949_,
		_w5967_,
		_w5968_,
		_w5970_
	);
	LUT2 #(
		.INIT('h2)
	) name5937 (
		_w5938_,
		_w5940_,
		_w5971_
	);
	LUT2 #(
		.INIT('h9)
	) name5938 (
		_w5938_,
		_w5940_,
		_w5972_
	);
	LUT3 #(
		.INIT('h69)
	) name5939 (
		\a[11] ,
		_w5931_,
		_w5932_,
		_w5973_
	);
	LUT4 #(
		.INIT('h4d00)
	) name5940 (
		_w5938_,
		_w5940_,
		_w5970_,
		_w5973_,
		_w5974_
	);
	LUT2 #(
		.INIT('h2)
	) name5941 (
		_w5924_,
		_w5925_,
		_w5975_
	);
	LUT2 #(
		.INIT('h9)
	) name5942 (
		_w5924_,
		_w5925_,
		_w5976_
	);
	LUT4 #(
		.INIT('h5501)
	) name5943 (
		_w5926_,
		_w5933_,
		_w5974_,
		_w5975_,
		_w5977_
	);
	LUT4 #(
		.INIT('h1428)
	) name5944 (
		\a[11] ,
		_w5704_,
		_w5706_,
		_w5917_,
		_w5978_
	);
	LUT4 #(
		.INIT('h6996)
	) name5945 (
		\a[11] ,
		_w5704_,
		_w5706_,
		_w5917_,
		_w5979_
	);
	LUT2 #(
		.INIT('h9)
	) name5946 (
		_w5905_,
		_w5910_,
		_w5980_
	);
	LUT4 #(
		.INIT('h2b00)
	) name5947 (
		_w5912_,
		_w5918_,
		_w5977_,
		_w5980_,
		_w5981_
	);
	LUT2 #(
		.INIT('h4)
	) name5948 (
		_w5897_,
		_w5903_,
		_w5982_
	);
	LUT2 #(
		.INIT('h9)
	) name5949 (
		_w5897_,
		_w5903_,
		_w5983_
	);
	LUT4 #(
		.INIT('h5501)
	) name5950 (
		_w5904_,
		_w5911_,
		_w5981_,
		_w5982_,
		_w5984_
	);
	LUT3 #(
		.INIT('h60)
	) name5951 (
		_w5711_,
		_w5713_,
		_w5895_,
		_w5985_
	);
	LUT3 #(
		.INIT('h96)
	) name5952 (
		_w5711_,
		_w5713_,
		_w5895_,
		_w5986_
	);
	LUT2 #(
		.INIT('h9)
	) name5953 (
		_w5888_,
		_w5889_,
		_w5987_
	);
	LUT4 #(
		.INIT('hba00)
	) name5954 (
		_w5896_,
		_w5984_,
		_w5986_,
		_w5987_,
		_w5988_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name5955 (
		_w5645_,
		_w5715_,
		_w5717_,
		_w5881_,
		_w5989_
	);
	LUT4 #(
		.INIT('h0155)
	) name5956 (
		_w5882_,
		_w5890_,
		_w5988_,
		_w5989_,
		_w5990_
	);
	LUT3 #(
		.INIT('h60)
	) name5957 (
		_w5718_,
		_w5720_,
		_w5875_,
		_w5991_
	);
	LUT3 #(
		.INIT('h96)
	) name5958 (
		_w5718_,
		_w5720_,
		_w5875_,
		_w5992_
	);
	LUT2 #(
		.INIT('h9)
	) name5959 (
		_w5862_,
		_w5867_,
		_w5993_
	);
	LUT4 #(
		.INIT('h2b00)
	) name5960 (
		_w5869_,
		_w5875_,
		_w5990_,
		_w5993_,
		_w5994_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name5961 (
		_w5624_,
		_w5722_,
		_w5723_,
		_w5860_,
		_w5995_
	);
	LUT4 #(
		.INIT('h0155)
	) name5962 (
		_w5861_,
		_w5868_,
		_w5994_,
		_w5995_,
		_w5996_
	);
	LUT3 #(
		.INIT('h60)
	) name5963 (
		_w5724_,
		_w5726_,
		_w5853_,
		_w5997_
	);
	LUT3 #(
		.INIT('h96)
	) name5964 (
		_w5724_,
		_w5726_,
		_w5853_,
		_w5998_
	);
	LUT2 #(
		.INIT('h9)
	) name5965 (
		_w5846_,
		_w5847_,
		_w5999_
	);
	LUT4 #(
		.INIT('hba00)
	) name5966 (
		_w5854_,
		_w5996_,
		_w5998_,
		_w5999_,
		_w6000_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name5967 (
		_w5602_,
		_w5728_,
		_w5729_,
		_w5839_,
		_w6001_
	);
	LUT4 #(
		.INIT('h0155)
	) name5968 (
		_w5840_,
		_w5848_,
		_w6000_,
		_w6001_,
		_w6002_
	);
	LUT3 #(
		.INIT('h60)
	) name5969 (
		_w5730_,
		_w5732_,
		_w5833_,
		_w6003_
	);
	LUT3 #(
		.INIT('h96)
	) name5970 (
		_w5730_,
		_w5732_,
		_w5833_,
		_w6004_
	);
	LUT2 #(
		.INIT('h9)
	) name5971 (
		_w5820_,
		_w5825_,
		_w6005_
	);
	LUT4 #(
		.INIT('h2b00)
	) name5972 (
		_w5827_,
		_w5833_,
		_w6002_,
		_w6005_,
		_w6006_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name5973 (
		_w5582_,
		_w5734_,
		_w5735_,
		_w5818_,
		_w6007_
	);
	LUT4 #(
		.INIT('h0155)
	) name5974 (
		_w5819_,
		_w5826_,
		_w6006_,
		_w6007_,
		_w6008_
	);
	LUT3 #(
		.INIT('h60)
	) name5975 (
		_w5736_,
		_w5738_,
		_w5811_,
		_w6009_
	);
	LUT3 #(
		.INIT('h96)
	) name5976 (
		_w5736_,
		_w5738_,
		_w5811_,
		_w6010_
	);
	LUT2 #(
		.INIT('h9)
	) name5977 (
		_w5804_,
		_w5805_,
		_w6011_
	);
	LUT4 #(
		.INIT('hba00)
	) name5978 (
		_w5812_,
		_w6008_,
		_w6010_,
		_w6011_,
		_w6012_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name5979 (
		_w5560_,
		_w5740_,
		_w5741_,
		_w5797_,
		_w6013_
	);
	LUT4 #(
		.INIT('h0155)
	) name5980 (
		_w5798_,
		_w5806_,
		_w6012_,
		_w6013_,
		_w6014_
	);
	LUT3 #(
		.INIT('h60)
	) name5981 (
		_w5742_,
		_w5744_,
		_w5790_,
		_w6015_
	);
	LUT3 #(
		.INIT('h96)
	) name5982 (
		_w5742_,
		_w5744_,
		_w5790_,
		_w6016_
	);
	LUT2 #(
		.INIT('h9)
	) name5983 (
		_w5782_,
		_w5783_,
		_w6017_
	);
	LUT4 #(
		.INIT('h4d00)
	) name5984 (
		_w5790_,
		_w5791_,
		_w6014_,
		_w6017_,
		_w6018_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name5985 (
		_w5540_,
		_w5746_,
		_w5747_,
		_w5776_,
		_w6019_
	);
	LUT4 #(
		.INIT('h0155)
	) name5986 (
		_w5777_,
		_w5784_,
		_w6018_,
		_w6019_,
		_w6020_
	);
	LUT3 #(
		.INIT('h96)
	) name5987 (
		_w5748_,
		_w5749_,
		_w5754_,
		_w6021_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5988 (
		_w587_,
		_w608_,
		_w624_,
		_w5271_,
		_w6022_
	);
	LUT3 #(
		.INIT('h70)
	) name5989 (
		_w666_,
		_w694_,
		_w4875_,
		_w6023_
	);
	LUT3 #(
		.INIT('h70)
	) name5990 (
		_w544_,
		_w558_,
		_w5286_,
		_w6024_
	);
	LUT3 #(
		.INIT('h01)
	) name5991 (
		_w6023_,
		_w6024_,
		_w6022_,
		_w6025_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5992 (
		_w2351_,
		_w2353_,
		_w4876_,
		_w6025_,
		_w6026_
	);
	LUT2 #(
		.INIT('h6)
	) name5993 (
		\a[8] ,
		_w6026_,
		_w6027_
	);
	LUT3 #(
		.INIT('hb2)
	) name5994 (
		_w6020_,
		_w6021_,
		_w6027_,
		_w6028_
	);
	LUT4 #(
		.INIT('hf400)
	) name5995 (
		_w374_,
		_w2361_,
		_w2404_,
		_w35_,
		_w6029_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5996 (
		_w121_,
		_w418_,
		_w422_,
		_w5524_,
		_w6030_
	);
	LUT3 #(
		.INIT('h18)
	) name5997 (
		\a[2] ,
		\a[3] ,
		\a[4] ,
		_w6031_
	);
	LUT3 #(
		.INIT('h70)
	) name5998 (
		_w352_,
		_w373_,
		_w6031_,
		_w6032_
	);
	LUT2 #(
		.INIT('h1)
	) name5999 (
		_w6030_,
		_w6032_,
		_w6033_
	);
	LUT3 #(
		.INIT('h9a)
	) name6000 (
		\a[5] ,
		_w6029_,
		_w6033_,
		_w6034_
	);
	LUT4 #(
		.INIT('h004d)
	) name6001 (
		_w6020_,
		_w6021_,
		_w6027_,
		_w6034_,
		_w6035_
	);
	LUT4 #(
		.INIT('hb200)
	) name6002 (
		_w6020_,
		_w6021_,
		_w6027_,
		_w6034_,
		_w6036_
	);
	LUT4 #(
		.INIT('h4db2)
	) name6003 (
		_w6020_,
		_w6021_,
		_w6027_,
		_w6034_,
		_w6037_
	);
	LUT4 #(
		.INIT('h4db2)
	) name6004 (
		_w5748_,
		_w5749_,
		_w5754_,
		_w5757_,
		_w6038_
	);
	LUT2 #(
		.INIT('h9)
	) name6005 (
		_w5764_,
		_w6038_,
		_w6039_
	);
	LUT3 #(
		.INIT('h45)
	) name6006 (
		_w6035_,
		_w6036_,
		_w6039_,
		_w6040_
	);
	LUT4 #(
		.INIT('h999a)
	) name6007 (
		_w5526_,
		_w5758_,
		_w5759_,
		_w5764_,
		_w6041_
	);
	LUT2 #(
		.INIT('h6)
	) name6008 (
		_w5769_,
		_w6041_,
		_w6042_
	);
	LUT4 #(
		.INIT('h7100)
	) name6009 (
		_w6028_,
		_w6034_,
		_w6039_,
		_w6042_,
		_w6043_
	);
	LUT4 #(
		.INIT('h45ba)
	) name6010 (
		_w6035_,
		_w6036_,
		_w6039_,
		_w6042_,
		_w6044_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6011 (
		_w587_,
		_w608_,
		_w624_,
		_w5286_,
		_w6045_
	);
	LUT3 #(
		.INIT('h70)
	) name6012 (
		_w725_,
		_w764_,
		_w4875_,
		_w6046_
	);
	LUT3 #(
		.INIT('h70)
	) name6013 (
		_w666_,
		_w694_,
		_w5271_,
		_w6047_
	);
	LUT3 #(
		.INIT('h01)
	) name6014 (
		_w6046_,
		_w6047_,
		_w6045_,
		_w6048_
	);
	LUT4 #(
		.INIT('h95aa)
	) name6015 (
		\a[8] ,
		_w2598_,
		_w4876_,
		_w6048_,
		_w6049_
	);
	LUT4 #(
		.INIT('h001e)
	) name6016 (
		_w5784_,
		_w6018_,
		_w6019_,
		_w6049_,
		_w6050_
	);
	LUT4 #(
		.INIT('h54ab)
	) name6017 (
		_w5792_,
		_w6014_,
		_w6015_,
		_w6017_,
		_w6051_
	);
	LUT3 #(
		.INIT('h70)
	) name6018 (
		_w725_,
		_w764_,
		_w5271_,
		_w6052_
	);
	LUT3 #(
		.INIT('h70)
	) name6019 (
		_w801_,
		_w851_,
		_w4875_,
		_w6053_
	);
	LUT3 #(
		.INIT('h70)
	) name6020 (
		_w666_,
		_w694_,
		_w5286_,
		_w6054_
	);
	LUT3 #(
		.INIT('h01)
	) name6021 (
		_w6053_,
		_w6054_,
		_w6052_,
		_w6055_
	);
	LUT4 #(
		.INIT('h6f00)
	) name6022 (
		_w2347_,
		_w2349_,
		_w4876_,
		_w6055_,
		_w6056_
	);
	LUT2 #(
		.INIT('h6)
	) name6023 (
		\a[8] ,
		_w6056_,
		_w6057_
	);
	LUT2 #(
		.INIT('h2)
	) name6024 (
		_w6051_,
		_w6057_,
		_w6058_
	);
	LUT3 #(
		.INIT('h70)
	) name6025 (
		_w725_,
		_w764_,
		_w5286_,
		_w6059_
	);
	LUT3 #(
		.INIT('h70)
	) name6026 (
		_w801_,
		_w851_,
		_w5271_,
		_w6060_
	);
	LUT3 #(
		.INIT('h70)
	) name6027 (
		_w871_,
		_w927_,
		_w4875_,
		_w6061_
	);
	LUT3 #(
		.INIT('h01)
	) name6028 (
		_w6060_,
		_w6061_,
		_w6059_,
		_w6062_
	);
	LUT4 #(
		.INIT('h95aa)
	) name6029 (
		\a[8] ,
		_w2724_,
		_w4876_,
		_w6062_,
		_w6063_
	);
	LUT3 #(
		.INIT('h09)
	) name6030 (
		_w6014_,
		_w6016_,
		_w6063_,
		_w6064_
	);
	LUT3 #(
		.INIT('h70)
	) name6031 (
		_w763_,
		_w983_,
		_w4875_,
		_w6065_
	);
	LUT3 #(
		.INIT('h70)
	) name6032 (
		_w871_,
		_w927_,
		_w5271_,
		_w6066_
	);
	LUT3 #(
		.INIT('h70)
	) name6033 (
		_w801_,
		_w851_,
		_w5286_,
		_w6067_
	);
	LUT3 #(
		.INIT('h01)
	) name6034 (
		_w6066_,
		_w6067_,
		_w6065_,
		_w6068_
	);
	LUT4 #(
		.INIT('h6f00)
	) name6035 (
		_w2343_,
		_w2345_,
		_w4876_,
		_w6068_,
		_w6069_
	);
	LUT2 #(
		.INIT('h6)
	) name6036 (
		\a[8] ,
		_w6069_,
		_w6070_
	);
	LUT4 #(
		.INIT('h001e)
	) name6037 (
		_w5806_,
		_w6012_,
		_w6013_,
		_w6070_,
		_w6071_
	);
	LUT4 #(
		.INIT('h54ab)
	) name6038 (
		_w5812_,
		_w6008_,
		_w6009_,
		_w6011_,
		_w6072_
	);
	LUT3 #(
		.INIT('h70)
	) name6039 (
		_w1009_,
		_w1050_,
		_w4875_,
		_w6073_
	);
	LUT3 #(
		.INIT('h70)
	) name6040 (
		_w871_,
		_w927_,
		_w5286_,
		_w6074_
	);
	LUT3 #(
		.INIT('h70)
	) name6041 (
		_w763_,
		_w983_,
		_w5271_,
		_w6075_
	);
	LUT3 #(
		.INIT('h01)
	) name6042 (
		_w6074_,
		_w6075_,
		_w6073_,
		_w6076_
	);
	LUT4 #(
		.INIT('h95aa)
	) name6043 (
		\a[8] ,
		_w2839_,
		_w4876_,
		_w6076_,
		_w6077_
	);
	LUT2 #(
		.INIT('h2)
	) name6044 (
		_w6072_,
		_w6077_,
		_w6078_
	);
	LUT2 #(
		.INIT('h9)
	) name6045 (
		_w6008_,
		_w6010_,
		_w6079_
	);
	LUT3 #(
		.INIT('h70)
	) name6046 (
		_w1071_,
		_w1102_,
		_w4875_,
		_w6080_
	);
	LUT3 #(
		.INIT('h70)
	) name6047 (
		_w763_,
		_w983_,
		_w5286_,
		_w6081_
	);
	LUT3 #(
		.INIT('h70)
	) name6048 (
		_w1009_,
		_w1050_,
		_w5271_,
		_w6082_
	);
	LUT3 #(
		.INIT('h01)
	) name6049 (
		_w6081_,
		_w6082_,
		_w6080_,
		_w6083_
	);
	LUT4 #(
		.INIT('h6f00)
	) name6050 (
		_w2339_,
		_w2341_,
		_w4876_,
		_w6083_,
		_w6084_
	);
	LUT2 #(
		.INIT('h6)
	) name6051 (
		\a[8] ,
		_w6084_,
		_w6085_
	);
	LUT3 #(
		.INIT('h09)
	) name6052 (
		_w6008_,
		_w6010_,
		_w6085_,
		_w6086_
	);
	LUT3 #(
		.INIT('h70)
	) name6053 (
		_w1136_,
		_w1187_,
		_w4875_,
		_w6087_
	);
	LUT3 #(
		.INIT('h70)
	) name6054 (
		_w1009_,
		_w1050_,
		_w5286_,
		_w6088_
	);
	LUT3 #(
		.INIT('h70)
	) name6055 (
		_w1071_,
		_w1102_,
		_w5271_,
		_w6089_
	);
	LUT3 #(
		.INIT('h01)
	) name6056 (
		_w6088_,
		_w6089_,
		_w6087_,
		_w6090_
	);
	LUT4 #(
		.INIT('h95aa)
	) name6057 (
		\a[8] ,
		_w2936_,
		_w4876_,
		_w6090_,
		_w6091_
	);
	LUT4 #(
		.INIT('h001e)
	) name6058 (
		_w5826_,
		_w6006_,
		_w6007_,
		_w6091_,
		_w6092_
	);
	LUT3 #(
		.INIT('h70)
	) name6059 (
		_w1136_,
		_w1187_,
		_w5271_,
		_w6093_
	);
	LUT3 #(
		.INIT('h70)
	) name6060 (
		_w1071_,
		_w1102_,
		_w5286_,
		_w6094_
	);
	LUT3 #(
		.INIT('h70)
	) name6061 (
		_w1202_,
		_w1233_,
		_w4875_,
		_w6095_
	);
	LUT3 #(
		.INIT('h01)
	) name6062 (
		_w6094_,
		_w6095_,
		_w6093_,
		_w6096_
	);
	LUT4 #(
		.INIT('h6f00)
	) name6063 (
		_w2335_,
		_w2337_,
		_w4876_,
		_w6096_,
		_w6097_
	);
	LUT2 #(
		.INIT('h6)
	) name6064 (
		\a[8] ,
		_w6097_,
		_w6098_
	);
	LUT4 #(
		.INIT('h54ab)
	) name6065 (
		_w5834_,
		_w6002_,
		_w6003_,
		_w6005_,
		_w6099_
	);
	LUT2 #(
		.INIT('h4)
	) name6066 (
		_w6098_,
		_w6099_,
		_w6100_
	);
	LUT3 #(
		.INIT('h70)
	) name6067 (
		_w1202_,
		_w1233_,
		_w5271_,
		_w6101_
	);
	LUT3 #(
		.INIT('h70)
	) name6068 (
		_w1253_,
		_w1294_,
		_w4875_,
		_w6102_
	);
	LUT3 #(
		.INIT('h70)
	) name6069 (
		_w1136_,
		_w1187_,
		_w5286_,
		_w6103_
	);
	LUT3 #(
		.INIT('h01)
	) name6070 (
		_w6102_,
		_w6103_,
		_w6101_,
		_w6104_
	);
	LUT4 #(
		.INIT('h95aa)
	) name6071 (
		\a[8] ,
		_w3067_,
		_w4876_,
		_w6104_,
		_w6105_
	);
	LUT3 #(
		.INIT('h09)
	) name6072 (
		_w6002_,
		_w6004_,
		_w6105_,
		_w6106_
	);
	LUT3 #(
		.INIT('h70)
	) name6073 (
		_w1202_,
		_w1233_,
		_w5286_,
		_w6107_
	);
	LUT3 #(
		.INIT('h70)
	) name6074 (
		_w1325_,
		_w1367_,
		_w4875_,
		_w6108_
	);
	LUT3 #(
		.INIT('h70)
	) name6075 (
		_w1253_,
		_w1294_,
		_w5271_,
		_w6109_
	);
	LUT3 #(
		.INIT('h01)
	) name6076 (
		_w6108_,
		_w6109_,
		_w6107_,
		_w6110_
	);
	LUT4 #(
		.INIT('h6f00)
	) name6077 (
		_w2331_,
		_w2333_,
		_w4876_,
		_w6110_,
		_w6111_
	);
	LUT2 #(
		.INIT('h6)
	) name6078 (
		\a[8] ,
		_w6111_,
		_w6112_
	);
	LUT4 #(
		.INIT('h001e)
	) name6079 (
		_w5848_,
		_w6000_,
		_w6001_,
		_w6112_,
		_w6113_
	);
	LUT4 #(
		.INIT('h54ab)
	) name6080 (
		_w5854_,
		_w5996_,
		_w5997_,
		_w5999_,
		_w6114_
	);
	LUT3 #(
		.INIT('h70)
	) name6081 (
		_w1381_,
		_w1398_,
		_w4875_,
		_w6115_
	);
	LUT3 #(
		.INIT('h70)
	) name6082 (
		_w1325_,
		_w1367_,
		_w5271_,
		_w6116_
	);
	LUT3 #(
		.INIT('h70)
	) name6083 (
		_w1253_,
		_w1294_,
		_w5286_,
		_w6117_
	);
	LUT3 #(
		.INIT('h01)
	) name6084 (
		_w6116_,
		_w6117_,
		_w6115_,
		_w6118_
	);
	LUT4 #(
		.INIT('h95aa)
	) name6085 (
		\a[8] ,
		_w3182_,
		_w4876_,
		_w6118_,
		_w6119_
	);
	LUT2 #(
		.INIT('h2)
	) name6086 (
		_w6114_,
		_w6119_,
		_w6120_
	);
	LUT2 #(
		.INIT('h9)
	) name6087 (
		_w5996_,
		_w5998_,
		_w6121_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6088 (
		_w1454_,
		_w1426_,
		_w1478_,
		_w4875_,
		_w6122_
	);
	LUT3 #(
		.INIT('h70)
	) name6089 (
		_w1325_,
		_w1367_,
		_w5286_,
		_w6123_
	);
	LUT3 #(
		.INIT('h70)
	) name6090 (
		_w1381_,
		_w1398_,
		_w5271_,
		_w6124_
	);
	LUT3 #(
		.INIT('h01)
	) name6091 (
		_w6123_,
		_w6124_,
		_w6122_,
		_w6125_
	);
	LUT4 #(
		.INIT('h6f00)
	) name6092 (
		_w2327_,
		_w2329_,
		_w4876_,
		_w6125_,
		_w6126_
	);
	LUT2 #(
		.INIT('h6)
	) name6093 (
		\a[8] ,
		_w6126_,
		_w6127_
	);
	LUT3 #(
		.INIT('h09)
	) name6094 (
		_w5996_,
		_w5998_,
		_w6127_,
		_w6128_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6095 (
		_w1454_,
		_w1426_,
		_w1478_,
		_w5271_,
		_w6129_
	);
	LUT3 #(
		.INIT('h70)
	) name6096 (
		_w1381_,
		_w1398_,
		_w5286_,
		_w6130_
	);
	LUT3 #(
		.INIT('h70)
	) name6097 (
		_w1501_,
		_w1545_,
		_w4875_,
		_w6131_
	);
	LUT3 #(
		.INIT('h01)
	) name6098 (
		_w6130_,
		_w6131_,
		_w6129_,
		_w6132_
	);
	LUT4 #(
		.INIT('h95aa)
	) name6099 (
		\a[8] ,
		_w3362_,
		_w4876_,
		_w6132_,
		_w6133_
	);
	LUT4 #(
		.INIT('h001e)
	) name6100 (
		_w5868_,
		_w5994_,
		_w5995_,
		_w6133_,
		_w6134_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6101 (
		_w1454_,
		_w1426_,
		_w1478_,
		_w5286_,
		_w6135_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6102 (
		_w1584_,
		_w1569_,
		_w1606_,
		_w4875_,
		_w6136_
	);
	LUT3 #(
		.INIT('h70)
	) name6103 (
		_w1501_,
		_w1545_,
		_w5271_,
		_w6137_
	);
	LUT3 #(
		.INIT('h01)
	) name6104 (
		_w6136_,
		_w6137_,
		_w6135_,
		_w6138_
	);
	LUT4 #(
		.INIT('h6f00)
	) name6105 (
		_w2323_,
		_w2325_,
		_w4876_,
		_w6138_,
		_w6139_
	);
	LUT2 #(
		.INIT('h6)
	) name6106 (
		\a[8] ,
		_w6139_,
		_w6140_
	);
	LUT4 #(
		.INIT('h54ab)
	) name6107 (
		_w5876_,
		_w5990_,
		_w5991_,
		_w5993_,
		_w6141_
	);
	LUT2 #(
		.INIT('h4)
	) name6108 (
		_w6140_,
		_w6141_,
		_w6142_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6109 (
		_w1584_,
		_w1569_,
		_w1606_,
		_w5271_,
		_w6143_
	);
	LUT3 #(
		.INIT('h70)
	) name6110 (
		_w1501_,
		_w1545_,
		_w5286_,
		_w6144_
	);
	LUT3 #(
		.INIT('h70)
	) name6111 (
		_w1620_,
		_w1661_,
		_w4875_,
		_w6145_
	);
	LUT3 #(
		.INIT('h01)
	) name6112 (
		_w6143_,
		_w6144_,
		_w6145_,
		_w6146_
	);
	LUT4 #(
		.INIT('h95aa)
	) name6113 (
		\a[8] ,
		_w3495_,
		_w4876_,
		_w6146_,
		_w6147_
	);
	LUT3 #(
		.INIT('h09)
	) name6114 (
		_w5990_,
		_w5992_,
		_w6147_,
		_w6148_
	);
	LUT3 #(
		.INIT('h70)
	) name6115 (
		_w1692_,
		_w1723_,
		_w4875_,
		_w6149_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6116 (
		_w1584_,
		_w1569_,
		_w1606_,
		_w5286_,
		_w6150_
	);
	LUT3 #(
		.INIT('h70)
	) name6117 (
		_w1620_,
		_w1661_,
		_w5271_,
		_w6151_
	);
	LUT3 #(
		.INIT('h01)
	) name6118 (
		_w6150_,
		_w6151_,
		_w6149_,
		_w6152_
	);
	LUT4 #(
		.INIT('h6f00)
	) name6119 (
		_w2319_,
		_w2321_,
		_w4876_,
		_w6152_,
		_w6153_
	);
	LUT2 #(
		.INIT('h6)
	) name6120 (
		\a[8] ,
		_w6153_,
		_w6154_
	);
	LUT4 #(
		.INIT('h001e)
	) name6121 (
		_w5890_,
		_w5988_,
		_w5989_,
		_w6154_,
		_w6155_
	);
	LUT4 #(
		.INIT('h54ab)
	) name6122 (
		_w5896_,
		_w5984_,
		_w5985_,
		_w5987_,
		_w6156_
	);
	LUT3 #(
		.INIT('h70)
	) name6123 (
		_w1692_,
		_w1723_,
		_w5271_,
		_w6157_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6124 (
		_w1751_,
		_w1742_,
		_w1771_,
		_w4875_,
		_w6158_
	);
	LUT3 #(
		.INIT('h70)
	) name6125 (
		_w1620_,
		_w1661_,
		_w5286_,
		_w6159_
	);
	LUT3 #(
		.INIT('h01)
	) name6126 (
		_w6158_,
		_w6159_,
		_w6157_,
		_w6160_
	);
	LUT4 #(
		.INIT('h95aa)
	) name6127 (
		\a[8] ,
		_w3599_,
		_w4876_,
		_w6160_,
		_w6161_
	);
	LUT2 #(
		.INIT('h2)
	) name6128 (
		_w6156_,
		_w6161_,
		_w6162_
	);
	LUT2 #(
		.INIT('h9)
	) name6129 (
		_w5984_,
		_w5986_,
		_w6163_
	);
	LUT3 #(
		.INIT('h70)
	) name6130 (
		_w1692_,
		_w1723_,
		_w5286_,
		_w6164_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6131 (
		_w1751_,
		_w1742_,
		_w1771_,
		_w5271_,
		_w6165_
	);
	LUT3 #(
		.INIT('h70)
	) name6132 (
		_w1795_,
		_w1796_,
		_w4875_,
		_w6166_
	);
	LUT3 #(
		.INIT('h01)
	) name6133 (
		_w6165_,
		_w6166_,
		_w6164_,
		_w6167_
	);
	LUT4 #(
		.INIT('h6f00)
	) name6134 (
		_w2315_,
		_w2317_,
		_w4876_,
		_w6167_,
		_w6168_
	);
	LUT2 #(
		.INIT('h6)
	) name6135 (
		\a[8] ,
		_w6168_,
		_w6169_
	);
	LUT3 #(
		.INIT('h09)
	) name6136 (
		_w5984_,
		_w5986_,
		_w6169_,
		_w6170_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6137 (
		_w1751_,
		_w1742_,
		_w1771_,
		_w5286_,
		_w6171_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6138 (
		_w1817_,
		_w1799_,
		_w1840_,
		_w4875_,
		_w6172_
	);
	LUT3 #(
		.INIT('h70)
	) name6139 (
		_w1795_,
		_w1796_,
		_w5271_,
		_w6173_
	);
	LUT3 #(
		.INIT('h01)
	) name6140 (
		_w6172_,
		_w6173_,
		_w6171_,
		_w6174_
	);
	LUT4 #(
		.INIT('h95aa)
	) name6141 (
		\a[8] ,
		_w3909_,
		_w4876_,
		_w6174_,
		_w6175_
	);
	LUT4 #(
		.INIT('h001e)
	) name6142 (
		_w5911_,
		_w5981_,
		_w5983_,
		_w6175_,
		_w6176_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6143 (
		_w1817_,
		_w1799_,
		_w1840_,
		_w5271_,
		_w6177_
	);
	LUT3 #(
		.INIT('h70)
	) name6144 (
		_w1795_,
		_w1796_,
		_w5286_,
		_w6178_
	);
	LUT3 #(
		.INIT('h70)
	) name6145 (
		_w1863_,
		_w1875_,
		_w4875_,
		_w6179_
	);
	LUT3 #(
		.INIT('h01)
	) name6146 (
		_w6178_,
		_w6179_,
		_w6177_,
		_w6180_
	);
	LUT4 #(
		.INIT('h6f00)
	) name6147 (
		_w2311_,
		_w2313_,
		_w4876_,
		_w6180_,
		_w6181_
	);
	LUT2 #(
		.INIT('h6)
	) name6148 (
		\a[8] ,
		_w6181_,
		_w6182_
	);
	LUT4 #(
		.INIT('h54ab)
	) name6149 (
		_w5919_,
		_w5977_,
		_w5978_,
		_w5980_,
		_w6183_
	);
	LUT2 #(
		.INIT('h4)
	) name6150 (
		_w6182_,
		_w6183_,
		_w6184_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6151 (
		_w1817_,
		_w1799_,
		_w1840_,
		_w5286_,
		_w6185_
	);
	LUT3 #(
		.INIT('h70)
	) name6152 (
		_w1898_,
		_w1928_,
		_w4875_,
		_w6186_
	);
	LUT3 #(
		.INIT('h70)
	) name6153 (
		_w1863_,
		_w1875_,
		_w5271_,
		_w6187_
	);
	LUT3 #(
		.INIT('h01)
	) name6154 (
		_w6186_,
		_w6187_,
		_w6185_,
		_w6188_
	);
	LUT4 #(
		.INIT('h95aa)
	) name6155 (
		\a[8] ,
		_w3972_,
		_w4876_,
		_w6188_,
		_w6189_
	);
	LUT3 #(
		.INIT('h09)
	) name6156 (
		_w5977_,
		_w5979_,
		_w6189_,
		_w6190_
	);
	LUT3 #(
		.INIT('h1e)
	) name6157 (
		_w5933_,
		_w5974_,
		_w5976_,
		_w6191_
	);
	LUT3 #(
		.INIT('h70)
	) name6158 (
		_w1501_,
		_w1949_,
		_w4875_,
		_w6192_
	);
	LUT3 #(
		.INIT('h70)
	) name6159 (
		_w1898_,
		_w1928_,
		_w5271_,
		_w6193_
	);
	LUT3 #(
		.INIT('h70)
	) name6160 (
		_w1863_,
		_w1875_,
		_w5286_,
		_w6194_
	);
	LUT3 #(
		.INIT('h01)
	) name6161 (
		_w6193_,
		_w6194_,
		_w6192_,
		_w6195_
	);
	LUT4 #(
		.INIT('h6f00)
	) name6162 (
		_w2307_,
		_w2309_,
		_w4876_,
		_w6195_,
		_w6196_
	);
	LUT2 #(
		.INIT('h6)
	) name6163 (
		\a[8] ,
		_w6196_,
		_w6197_
	);
	LUT2 #(
		.INIT('h2)
	) name6164 (
		_w6191_,
		_w6197_,
		_w6198_
	);
	LUT4 #(
		.INIT('h54ab)
	) name6165 (
		_w5941_,
		_w5970_,
		_w5971_,
		_w5973_,
		_w6199_
	);
	LUT3 #(
		.INIT('h70)
	) name6166 (
		_w1973_,
		_w1997_,
		_w4875_,
		_w6200_
	);
	LUT3 #(
		.INIT('h70)
	) name6167 (
		_w1898_,
		_w1928_,
		_w5286_,
		_w6201_
	);
	LUT3 #(
		.INIT('h70)
	) name6168 (
		_w1501_,
		_w1949_,
		_w5271_,
		_w6202_
	);
	LUT3 #(
		.INIT('h01)
	) name6169 (
		_w6201_,
		_w6202_,
		_w6200_,
		_w6203_
	);
	LUT4 #(
		.INIT('h95aa)
	) name6170 (
		\a[8] ,
		_w4126_,
		_w4876_,
		_w6203_,
		_w6204_
	);
	LUT2 #(
		.INIT('h2)
	) name6171 (
		_w6199_,
		_w6204_,
		_w6205_
	);
	LUT2 #(
		.INIT('h9)
	) name6172 (
		_w5970_,
		_w5972_,
		_w6206_
	);
	LUT3 #(
		.INIT('h70)
	) name6173 (
		_w1973_,
		_w1997_,
		_w5271_,
		_w6207_
	);
	LUT3 #(
		.INIT('h70)
	) name6174 (
		_w1501_,
		_w1949_,
		_w5286_,
		_w6208_
	);
	LUT3 #(
		.INIT('h70)
	) name6175 (
		_w2023_,
		_w2055_,
		_w4875_,
		_w6209_
	);
	LUT3 #(
		.INIT('h01)
	) name6176 (
		_w6208_,
		_w6209_,
		_w6207_,
		_w6210_
	);
	LUT4 #(
		.INIT('h6f00)
	) name6177 (
		_w2303_,
		_w2305_,
		_w4876_,
		_w6210_,
		_w6211_
	);
	LUT2 #(
		.INIT('h6)
	) name6178 (
		\a[8] ,
		_w6211_,
		_w6212_
	);
	LUT4 #(
		.INIT('h8241)
	) name6179 (
		\a[8] ,
		_w5970_,
		_w5972_,
		_w6211_,
		_w6213_
	);
	LUT3 #(
		.INIT('h70)
	) name6180 (
		_w1973_,
		_w1997_,
		_w5286_,
		_w6214_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6181 (
		_w1874_,
		_w2076_,
		_w2099_,
		_w4875_,
		_w6215_
	);
	LUT3 #(
		.INIT('h70)
	) name6182 (
		_w2023_,
		_w2055_,
		_w5271_,
		_w6216_
	);
	LUT3 #(
		.INIT('h01)
	) name6183 (
		_w6215_,
		_w6216_,
		_w6214_,
		_w6217_
	);
	LUT4 #(
		.INIT('h95aa)
	) name6184 (
		\a[8] ,
		_w4151_,
		_w4876_,
		_w6217_,
		_w6218_
	);
	LUT2 #(
		.INIT('h9)
	) name6185 (
		_w5967_,
		_w5969_,
		_w6219_
	);
	LUT2 #(
		.INIT('h4)
	) name6186 (
		_w6218_,
		_w6219_,
		_w6220_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6187 (
		_w1874_,
		_w2076_,
		_w2099_,
		_w5271_,
		_w6221_
	);
	LUT3 #(
		.INIT('h70)
	) name6188 (
		_w2124_,
		_w2133_,
		_w4875_,
		_w6222_
	);
	LUT3 #(
		.INIT('h70)
	) name6189 (
		_w2023_,
		_w2055_,
		_w5286_,
		_w6223_
	);
	LUT3 #(
		.INIT('h01)
	) name6190 (
		_w6221_,
		_w6222_,
		_w6223_,
		_w6224_
	);
	LUT4 #(
		.INIT('h6f00)
	) name6191 (
		_w2299_,
		_w2301_,
		_w4876_,
		_w6224_,
		_w6225_
	);
	LUT3 #(
		.INIT('h69)
	) name6192 (
		_w5687_,
		_w5961_,
		_w5966_,
		_w6226_
	);
	LUT3 #(
		.INIT('h90)
	) name6193 (
		\a[8] ,
		_w6225_,
		_w6226_,
		_w6227_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6194 (
		_w1874_,
		_w2076_,
		_w2099_,
		_w5286_,
		_w6228_
	);
	LUT3 #(
		.INIT('h70)
	) name6195 (
		_w2124_,
		_w2133_,
		_w5271_,
		_w6229_
	);
	LUT3 #(
		.INIT('h70)
	) name6196 (
		_w2155_,
		_w2156_,
		_w4875_,
		_w6230_
	);
	LUT3 #(
		.INIT('h01)
	) name6197 (
		_w6228_,
		_w6229_,
		_w6230_,
		_w6231_
	);
	LUT4 #(
		.INIT('h95aa)
	) name6198 (
		\a[8] ,
		_w4209_,
		_w4876_,
		_w6231_,
		_w6232_
	);
	LUT3 #(
		.INIT('h8a)
	) name6199 (
		\a[11] ,
		_w5953_,
		_w5952_,
		_w6233_
	);
	LUT2 #(
		.INIT('h9)
	) name6200 (
		_w5960_,
		_w6233_,
		_w6234_
	);
	LUT2 #(
		.INIT('h4)
	) name6201 (
		_w6232_,
		_w6234_,
		_w6235_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6202 (
		_w2193_,
		_w2183_,
		_w2213_,
		_w4875_,
		_w6236_
	);
	LUT3 #(
		.INIT('h70)
	) name6203 (
		_w2155_,
		_w2156_,
		_w5271_,
		_w6237_
	);
	LUT3 #(
		.INIT('h70)
	) name6204 (
		_w2124_,
		_w2133_,
		_w5286_,
		_w6238_
	);
	LUT3 #(
		.INIT('h01)
	) name6205 (
		_w6236_,
		_w6237_,
		_w6238_,
		_w6239_
	);
	LUT4 #(
		.INIT('h6f00)
	) name6206 (
		_w2295_,
		_w2297_,
		_w4876_,
		_w6239_,
		_w6240_
	);
	LUT4 #(
		.INIT('h002a)
	) name6207 (
		\a[11] ,
		_w2228_,
		_w2262_,
		_w4457_,
		_w6241_
	);
	LUT2 #(
		.INIT('h9)
	) name6208 (
		_w5952_,
		_w6241_,
		_w6242_
	);
	LUT3 #(
		.INIT('h90)
	) name6209 (
		\a[8] ,
		_w6240_,
		_w6242_,
		_w6243_
	);
	LUT3 #(
		.INIT('h70)
	) name6210 (
		_w2228_,
		_w2262_,
		_w5271_,
		_w6244_
	);
	LUT3 #(
		.INIT('h70)
	) name6211 (
		_w2273_,
		_w2293_,
		_w5286_,
		_w6245_
	);
	LUT4 #(
		.INIT('h000b)
	) name6212 (
		_w4599_,
		_w4876_,
		_w6244_,
		_w6245_,
		_w6246_
	);
	LUT3 #(
		.INIT('h07)
	) name6213 (
		_w2228_,
		_w2262_,
		_w4874_,
		_w6247_
	);
	LUT4 #(
		.INIT('haa80)
	) name6214 (
		\a[8] ,
		_w2228_,
		_w2262_,
		_w4874_,
		_w6248_
	);
	LUT3 #(
		.INIT('h90)
	) name6215 (
		_w2214_,
		_w4258_,
		_w4876_,
		_w6249_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6216 (
		_w2193_,
		_w2183_,
		_w2213_,
		_w5286_,
		_w6250_
	);
	LUT3 #(
		.INIT('h70)
	) name6217 (
		_w2228_,
		_w2262_,
		_w4875_,
		_w6251_
	);
	LUT3 #(
		.INIT('h70)
	) name6218 (
		_w2273_,
		_w2293_,
		_w5271_,
		_w6252_
	);
	LUT3 #(
		.INIT('h01)
	) name6219 (
		_w6251_,
		_w6252_,
		_w6250_,
		_w6253_
	);
	LUT2 #(
		.INIT('h4)
	) name6220 (
		_w6249_,
		_w6253_,
		_w6254_
	);
	LUT4 #(
		.INIT('h0800)
	) name6221 (
		_w6246_,
		_w6248_,
		_w6249_,
		_w6253_,
		_w6255_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6222 (
		_w2193_,
		_w2183_,
		_w2213_,
		_w5271_,
		_w6256_
	);
	LUT3 #(
		.INIT('h70)
	) name6223 (
		_w2155_,
		_w2156_,
		_w5286_,
		_w6257_
	);
	LUT3 #(
		.INIT('h70)
	) name6224 (
		_w2273_,
		_w2293_,
		_w4875_,
		_w6258_
	);
	LUT3 #(
		.INIT('h01)
	) name6225 (
		_w6256_,
		_w6257_,
		_w6258_,
		_w6259_
	);
	LUT4 #(
		.INIT('h95aa)
	) name6226 (
		\a[8] ,
		_w4293_,
		_w4876_,
		_w6259_,
		_w6260_
	);
	LUT3 #(
		.INIT('h71)
	) name6227 (
		_w5953_,
		_w6255_,
		_w6260_,
		_w6261_
	);
	LUT3 #(
		.INIT('h06)
	) name6228 (
		\a[8] ,
		_w6240_,
		_w6242_,
		_w6262_
	);
	LUT3 #(
		.INIT('h69)
	) name6229 (
		\a[8] ,
		_w6240_,
		_w6242_,
		_w6263_
	);
	LUT3 #(
		.INIT('h54)
	) name6230 (
		_w6243_,
		_w6261_,
		_w6262_,
		_w6264_
	);
	LUT2 #(
		.INIT('h2)
	) name6231 (
		_w6232_,
		_w6234_,
		_w6265_
	);
	LUT2 #(
		.INIT('h9)
	) name6232 (
		_w6232_,
		_w6234_,
		_w6266_
	);
	LUT3 #(
		.INIT('h69)
	) name6233 (
		\a[8] ,
		_w6225_,
		_w6226_,
		_w6267_
	);
	LUT4 #(
		.INIT('h4d00)
	) name6234 (
		_w6232_,
		_w6234_,
		_w6264_,
		_w6267_,
		_w6268_
	);
	LUT2 #(
		.INIT('h2)
	) name6235 (
		_w6218_,
		_w6219_,
		_w6269_
	);
	LUT2 #(
		.INIT('h9)
	) name6236 (
		_w6218_,
		_w6219_,
		_w6270_
	);
	LUT4 #(
		.INIT('h5501)
	) name6237 (
		_w6220_,
		_w6227_,
		_w6268_,
		_w6269_,
		_w6271_
	);
	LUT4 #(
		.INIT('h1428)
	) name6238 (
		\a[8] ,
		_w5970_,
		_w5972_,
		_w6211_,
		_w6272_
	);
	LUT4 #(
		.INIT('h6996)
	) name6239 (
		\a[8] ,
		_w5970_,
		_w5972_,
		_w6211_,
		_w6273_
	);
	LUT2 #(
		.INIT('h9)
	) name6240 (
		_w6199_,
		_w6204_,
		_w6274_
	);
	LUT4 #(
		.INIT('h2b00)
	) name6241 (
		_w6206_,
		_w6212_,
		_w6271_,
		_w6274_,
		_w6275_
	);
	LUT2 #(
		.INIT('h4)
	) name6242 (
		_w6191_,
		_w6197_,
		_w6276_
	);
	LUT2 #(
		.INIT('h9)
	) name6243 (
		_w6191_,
		_w6197_,
		_w6277_
	);
	LUT4 #(
		.INIT('h5501)
	) name6244 (
		_w6198_,
		_w6205_,
		_w6275_,
		_w6276_,
		_w6278_
	);
	LUT3 #(
		.INIT('h60)
	) name6245 (
		_w5977_,
		_w5979_,
		_w6189_,
		_w6279_
	);
	LUT3 #(
		.INIT('h96)
	) name6246 (
		_w5977_,
		_w5979_,
		_w6189_,
		_w6280_
	);
	LUT2 #(
		.INIT('h9)
	) name6247 (
		_w6182_,
		_w6183_,
		_w6281_
	);
	LUT4 #(
		.INIT('hba00)
	) name6248 (
		_w6190_,
		_w6278_,
		_w6280_,
		_w6281_,
		_w6282_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name6249 (
		_w5911_,
		_w5981_,
		_w5983_,
		_w6175_,
		_w6283_
	);
	LUT4 #(
		.INIT('h0155)
	) name6250 (
		_w6176_,
		_w6184_,
		_w6282_,
		_w6283_,
		_w6284_
	);
	LUT3 #(
		.INIT('h60)
	) name6251 (
		_w5984_,
		_w5986_,
		_w6169_,
		_w6285_
	);
	LUT3 #(
		.INIT('h96)
	) name6252 (
		_w5984_,
		_w5986_,
		_w6169_,
		_w6286_
	);
	LUT2 #(
		.INIT('h9)
	) name6253 (
		_w6156_,
		_w6161_,
		_w6287_
	);
	LUT4 #(
		.INIT('h2b00)
	) name6254 (
		_w6163_,
		_w6169_,
		_w6284_,
		_w6287_,
		_w6288_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name6255 (
		_w5890_,
		_w5988_,
		_w5989_,
		_w6154_,
		_w6289_
	);
	LUT4 #(
		.INIT('h0155)
	) name6256 (
		_w6155_,
		_w6162_,
		_w6288_,
		_w6289_,
		_w6290_
	);
	LUT3 #(
		.INIT('h60)
	) name6257 (
		_w5990_,
		_w5992_,
		_w6147_,
		_w6291_
	);
	LUT3 #(
		.INIT('h96)
	) name6258 (
		_w5990_,
		_w5992_,
		_w6147_,
		_w6292_
	);
	LUT2 #(
		.INIT('h9)
	) name6259 (
		_w6140_,
		_w6141_,
		_w6293_
	);
	LUT4 #(
		.INIT('hba00)
	) name6260 (
		_w6148_,
		_w6290_,
		_w6292_,
		_w6293_,
		_w6294_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name6261 (
		_w5868_,
		_w5994_,
		_w5995_,
		_w6133_,
		_w6295_
	);
	LUT4 #(
		.INIT('h0155)
	) name6262 (
		_w6134_,
		_w6142_,
		_w6294_,
		_w6295_,
		_w6296_
	);
	LUT3 #(
		.INIT('h60)
	) name6263 (
		_w5996_,
		_w5998_,
		_w6127_,
		_w6297_
	);
	LUT3 #(
		.INIT('h96)
	) name6264 (
		_w5996_,
		_w5998_,
		_w6127_,
		_w6298_
	);
	LUT2 #(
		.INIT('h9)
	) name6265 (
		_w6114_,
		_w6119_,
		_w6299_
	);
	LUT4 #(
		.INIT('h2b00)
	) name6266 (
		_w6121_,
		_w6127_,
		_w6296_,
		_w6299_,
		_w6300_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name6267 (
		_w5848_,
		_w6000_,
		_w6001_,
		_w6112_,
		_w6301_
	);
	LUT4 #(
		.INIT('h0155)
	) name6268 (
		_w6113_,
		_w6120_,
		_w6300_,
		_w6301_,
		_w6302_
	);
	LUT3 #(
		.INIT('h60)
	) name6269 (
		_w6002_,
		_w6004_,
		_w6105_,
		_w6303_
	);
	LUT3 #(
		.INIT('h96)
	) name6270 (
		_w6002_,
		_w6004_,
		_w6105_,
		_w6304_
	);
	LUT2 #(
		.INIT('h9)
	) name6271 (
		_w6098_,
		_w6099_,
		_w6305_
	);
	LUT4 #(
		.INIT('hba00)
	) name6272 (
		_w6106_,
		_w6302_,
		_w6304_,
		_w6305_,
		_w6306_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name6273 (
		_w5826_,
		_w6006_,
		_w6007_,
		_w6091_,
		_w6307_
	);
	LUT4 #(
		.INIT('h0155)
	) name6274 (
		_w6092_,
		_w6100_,
		_w6306_,
		_w6307_,
		_w6308_
	);
	LUT3 #(
		.INIT('h60)
	) name6275 (
		_w6008_,
		_w6010_,
		_w6085_,
		_w6309_
	);
	LUT3 #(
		.INIT('h96)
	) name6276 (
		_w6008_,
		_w6010_,
		_w6085_,
		_w6310_
	);
	LUT2 #(
		.INIT('h9)
	) name6277 (
		_w6072_,
		_w6077_,
		_w6311_
	);
	LUT4 #(
		.INIT('h2b00)
	) name6278 (
		_w6079_,
		_w6085_,
		_w6308_,
		_w6311_,
		_w6312_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name6279 (
		_w5806_,
		_w6012_,
		_w6013_,
		_w6070_,
		_w6313_
	);
	LUT4 #(
		.INIT('h0155)
	) name6280 (
		_w6071_,
		_w6078_,
		_w6312_,
		_w6313_,
		_w6314_
	);
	LUT3 #(
		.INIT('h60)
	) name6281 (
		_w6014_,
		_w6016_,
		_w6063_,
		_w6315_
	);
	LUT3 #(
		.INIT('h96)
	) name6282 (
		_w6014_,
		_w6016_,
		_w6063_,
		_w6316_
	);
	LUT2 #(
		.INIT('h9)
	) name6283 (
		_w6051_,
		_w6057_,
		_w6317_
	);
	LUT4 #(
		.INIT('hba00)
	) name6284 (
		_w6064_,
		_w6314_,
		_w6316_,
		_w6317_,
		_w6318_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name6285 (
		_w5784_,
		_w6018_,
		_w6019_,
		_w6049_,
		_w6319_
	);
	LUT4 #(
		.INIT('h0155)
	) name6286 (
		_w6050_,
		_w6058_,
		_w6318_,
		_w6319_,
		_w6320_
	);
	LUT3 #(
		.INIT('h96)
	) name6287 (
		_w6020_,
		_w6021_,
		_w6027_,
		_w6321_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6288 (
		_w486_,
		_w487_,
		_w509_,
		_w5524_,
		_w6322_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6289 (
		_w121_,
		_w418_,
		_w422_,
		_w6031_,
		_w6323_
	);
	LUT4 #(
		.INIT('h6006)
	) name6290 (
		\a[2] ,
		\a[3] ,
		\a[4] ,
		\a[5] ,
		_w6324_
	);
	LUT3 #(
		.INIT('h2a)
	) name6291 (
		_w6324_,
		_w352_,
		_w373_,
		_w6325_
	);
	LUT3 #(
		.INIT('h01)
	) name6292 (
		_w6322_,
		_w6323_,
		_w6325_,
		_w6326_
	);
	LUT4 #(
		.INIT('h95aa)
	) name6293 (
		\a[5] ,
		_w2535_,
		_w35_,
		_w6326_,
		_w6327_
	);
	LUT3 #(
		.INIT('hb2)
	) name6294 (
		_w6320_,
		_w6321_,
		_w6327_,
		_w6328_
	);
	LUT2 #(
		.INIT('h6)
	) name6295 (
		_w6037_,
		_w6039_,
		_w6329_
	);
	LUT4 #(
		.INIT('h4d00)
	) name6296 (
		_w6320_,
		_w6321_,
		_w6327_,
		_w6329_,
		_w6330_
	);
	LUT3 #(
		.INIT('h96)
	) name6297 (
		_w6320_,
		_w6321_,
		_w6327_,
		_w6331_
	);
	LUT2 #(
		.INIT('h1)
	) name6298 (
		\a[0] ,
		\a[1] ,
		_w6332_
	);
	LUT2 #(
		.INIT('h9)
	) name6299 (
		\a[1] ,
		\a[2] ,
		_w6333_
	);
	LUT3 #(
		.INIT('h10)
	) name6300 (
		\a[0] ,
		\a[1] ,
		\a[2] ,
		_w6334_
	);
	LUT3 #(
		.INIT('h28)
	) name6301 (
		\a[0] ,
		\a[1] ,
		\a[2] ,
		_w6335_
	);
	LUT4 #(
		.INIT('h5150)
	) name6302 (
		_w374_,
		_w2361_,
		_w6334_,
		_w6335_,
		_w6336_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6303 (
		_w486_,
		_w487_,
		_w509_,
		_w6031_,
		_w6337_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name6304 (
		_w6324_,
		_w121_,
		_w418_,
		_w422_,
		_w6338_
	);
	LUT3 #(
		.INIT('h70)
	) name6305 (
		_w544_,
		_w558_,
		_w5524_,
		_w6339_
	);
	LUT3 #(
		.INIT('h01)
	) name6306 (
		_w6337_,
		_w6338_,
		_w6339_,
		_w6340_
	);
	LUT4 #(
		.INIT('h6f00)
	) name6307 (
		_w2355_,
		_w2357_,
		_w35_,
		_w6340_,
		_w6341_
	);
	LUT2 #(
		.INIT('h6)
	) name6308 (
		\a[5] ,
		_w6341_,
		_w6342_
	);
	LUT3 #(
		.INIT('h06)
	) name6309 (
		\a[2] ,
		_w6336_,
		_w6342_,
		_w6343_
	);
	LUT3 #(
		.INIT('h90)
	) name6310 (
		\a[2] ,
		_w6336_,
		_w6342_,
		_w6344_
	);
	LUT4 #(
		.INIT('h001e)
	) name6311 (
		_w6058_,
		_w6318_,
		_w6319_,
		_w6344_,
		_w6345_
	);
	LUT2 #(
		.INIT('h1)
	) name6312 (
		_w6343_,
		_w6345_,
		_w6346_
	);
	LUT2 #(
		.INIT('h2)
	) name6313 (
		_w6331_,
		_w6346_,
		_w6347_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name6314 (
		_w6324_,
		_w486_,
		_w487_,
		_w509_,
		_w6348_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6315 (
		_w587_,
		_w608_,
		_w624_,
		_w5524_,
		_w6349_
	);
	LUT3 #(
		.INIT('h70)
	) name6316 (
		_w544_,
		_w558_,
		_w6031_,
		_w6350_
	);
	LUT3 #(
		.INIT('h01)
	) name6317 (
		_w6348_,
		_w6349_,
		_w6350_,
		_w6351_
	);
	LUT4 #(
		.INIT('h95aa)
	) name6318 (
		\a[5] ,
		_w2526_,
		_w35_,
		_w6351_,
		_w6352_
	);
	LUT4 #(
		.INIT('h54ab)
	) name6319 (
		_w6064_,
		_w6314_,
		_w6315_,
		_w6317_,
		_w6353_
	);
	LUT2 #(
		.INIT('h4)
	) name6320 (
		_w6352_,
		_w6353_,
		_w6354_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6321 (
		_w587_,
		_w608_,
		_w624_,
		_w6031_,
		_w6355_
	);
	LUT3 #(
		.INIT('h70)
	) name6322 (
		_w666_,
		_w694_,
		_w5524_,
		_w6356_
	);
	LUT3 #(
		.INIT('h2a)
	) name6323 (
		_w6324_,
		_w544_,
		_w558_,
		_w6357_
	);
	LUT3 #(
		.INIT('h01)
	) name6324 (
		_w6356_,
		_w6357_,
		_w6355_,
		_w6358_
	);
	LUT4 #(
		.INIT('h6f00)
	) name6325 (
		_w2351_,
		_w2353_,
		_w35_,
		_w6358_,
		_w6359_
	);
	LUT2 #(
		.INIT('h6)
	) name6326 (
		\a[5] ,
		_w6359_,
		_w6360_
	);
	LUT2 #(
		.INIT('h9)
	) name6327 (
		_w6314_,
		_w6316_,
		_w6361_
	);
	LUT3 #(
		.INIT('h09)
	) name6328 (
		_w6314_,
		_w6316_,
		_w6360_,
		_w6362_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name6329 (
		_w6324_,
		_w587_,
		_w608_,
		_w624_,
		_w6363_
	);
	LUT3 #(
		.INIT('h70)
	) name6330 (
		_w725_,
		_w764_,
		_w5524_,
		_w6364_
	);
	LUT3 #(
		.INIT('h70)
	) name6331 (
		_w666_,
		_w694_,
		_w6031_,
		_w6365_
	);
	LUT3 #(
		.INIT('h01)
	) name6332 (
		_w6364_,
		_w6365_,
		_w6363_,
		_w6366_
	);
	LUT4 #(
		.INIT('h95aa)
	) name6333 (
		\a[5] ,
		_w2598_,
		_w35_,
		_w6366_,
		_w6367_
	);
	LUT4 #(
		.INIT('h001e)
	) name6334 (
		_w6078_,
		_w6312_,
		_w6313_,
		_w6367_,
		_w6368_
	);
	LUT3 #(
		.INIT('h70)
	) name6335 (
		_w725_,
		_w764_,
		_w6031_,
		_w6369_
	);
	LUT3 #(
		.INIT('h70)
	) name6336 (
		_w801_,
		_w851_,
		_w5524_,
		_w6370_
	);
	LUT3 #(
		.INIT('h2a)
	) name6337 (
		_w6324_,
		_w666_,
		_w694_,
		_w6371_
	);
	LUT3 #(
		.INIT('h01)
	) name6338 (
		_w6370_,
		_w6371_,
		_w6369_,
		_w6372_
	);
	LUT4 #(
		.INIT('h6f00)
	) name6339 (
		_w2347_,
		_w2349_,
		_w35_,
		_w6372_,
		_w6373_
	);
	LUT2 #(
		.INIT('h6)
	) name6340 (
		\a[5] ,
		_w6373_,
		_w6374_
	);
	LUT4 #(
		.INIT('h54ab)
	) name6341 (
		_w6086_,
		_w6308_,
		_w6309_,
		_w6311_,
		_w6375_
	);
	LUT2 #(
		.INIT('h4)
	) name6342 (
		_w6374_,
		_w6375_,
		_w6376_
	);
	LUT3 #(
		.INIT('h2a)
	) name6343 (
		_w6324_,
		_w725_,
		_w764_,
		_w6377_
	);
	LUT3 #(
		.INIT('h70)
	) name6344 (
		_w801_,
		_w851_,
		_w6031_,
		_w6378_
	);
	LUT3 #(
		.INIT('h70)
	) name6345 (
		_w871_,
		_w927_,
		_w5524_,
		_w6379_
	);
	LUT3 #(
		.INIT('h01)
	) name6346 (
		_w6378_,
		_w6379_,
		_w6377_,
		_w6380_
	);
	LUT4 #(
		.INIT('h95aa)
	) name6347 (
		\a[5] ,
		_w2724_,
		_w35_,
		_w6380_,
		_w6381_
	);
	LUT3 #(
		.INIT('h09)
	) name6348 (
		_w6308_,
		_w6310_,
		_w6381_,
		_w6382_
	);
	LUT3 #(
		.INIT('h70)
	) name6349 (
		_w763_,
		_w983_,
		_w5524_,
		_w6383_
	);
	LUT3 #(
		.INIT('h70)
	) name6350 (
		_w871_,
		_w927_,
		_w6031_,
		_w6384_
	);
	LUT3 #(
		.INIT('h2a)
	) name6351 (
		_w6324_,
		_w801_,
		_w851_,
		_w6385_
	);
	LUT3 #(
		.INIT('h01)
	) name6352 (
		_w6384_,
		_w6385_,
		_w6383_,
		_w6386_
	);
	LUT4 #(
		.INIT('h6f00)
	) name6353 (
		_w2343_,
		_w2345_,
		_w35_,
		_w6386_,
		_w6387_
	);
	LUT2 #(
		.INIT('h6)
	) name6354 (
		\a[5] ,
		_w6387_,
		_w6388_
	);
	LUT4 #(
		.INIT('h001e)
	) name6355 (
		_w6100_,
		_w6306_,
		_w6307_,
		_w6388_,
		_w6389_
	);
	LUT4 #(
		.INIT('h54ab)
	) name6356 (
		_w6106_,
		_w6302_,
		_w6303_,
		_w6305_,
		_w6390_
	);
	LUT3 #(
		.INIT('h70)
	) name6357 (
		_w1009_,
		_w1050_,
		_w5524_,
		_w6391_
	);
	LUT3 #(
		.INIT('h2a)
	) name6358 (
		_w6324_,
		_w871_,
		_w927_,
		_w6392_
	);
	LUT3 #(
		.INIT('h70)
	) name6359 (
		_w763_,
		_w983_,
		_w6031_,
		_w6393_
	);
	LUT3 #(
		.INIT('h01)
	) name6360 (
		_w6392_,
		_w6393_,
		_w6391_,
		_w6394_
	);
	LUT4 #(
		.INIT('h95aa)
	) name6361 (
		\a[5] ,
		_w2839_,
		_w35_,
		_w6394_,
		_w6395_
	);
	LUT2 #(
		.INIT('h2)
	) name6362 (
		_w6390_,
		_w6395_,
		_w6396_
	);
	LUT2 #(
		.INIT('h9)
	) name6363 (
		_w6302_,
		_w6304_,
		_w6397_
	);
	LUT3 #(
		.INIT('h70)
	) name6364 (
		_w1071_,
		_w1102_,
		_w5524_,
		_w6398_
	);
	LUT3 #(
		.INIT('h2a)
	) name6365 (
		_w6324_,
		_w763_,
		_w983_,
		_w6399_
	);
	LUT3 #(
		.INIT('h70)
	) name6366 (
		_w1009_,
		_w1050_,
		_w6031_,
		_w6400_
	);
	LUT3 #(
		.INIT('h01)
	) name6367 (
		_w6399_,
		_w6400_,
		_w6398_,
		_w6401_
	);
	LUT4 #(
		.INIT('h6f00)
	) name6368 (
		_w2339_,
		_w2341_,
		_w35_,
		_w6401_,
		_w6402_
	);
	LUT2 #(
		.INIT('h6)
	) name6369 (
		\a[5] ,
		_w6402_,
		_w6403_
	);
	LUT3 #(
		.INIT('h09)
	) name6370 (
		_w6302_,
		_w6304_,
		_w6403_,
		_w6404_
	);
	LUT3 #(
		.INIT('h70)
	) name6371 (
		_w1136_,
		_w1187_,
		_w5524_,
		_w6405_
	);
	LUT3 #(
		.INIT('h2a)
	) name6372 (
		_w6324_,
		_w1009_,
		_w1050_,
		_w6406_
	);
	LUT3 #(
		.INIT('h70)
	) name6373 (
		_w1071_,
		_w1102_,
		_w6031_,
		_w6407_
	);
	LUT3 #(
		.INIT('h01)
	) name6374 (
		_w6406_,
		_w6407_,
		_w6405_,
		_w6408_
	);
	LUT4 #(
		.INIT('h95aa)
	) name6375 (
		\a[5] ,
		_w2936_,
		_w35_,
		_w6408_,
		_w6409_
	);
	LUT4 #(
		.INIT('h001e)
	) name6376 (
		_w6120_,
		_w6300_,
		_w6301_,
		_w6409_,
		_w6410_
	);
	LUT3 #(
		.INIT('h70)
	) name6377 (
		_w1136_,
		_w1187_,
		_w6031_,
		_w6411_
	);
	LUT3 #(
		.INIT('h2a)
	) name6378 (
		_w6324_,
		_w1071_,
		_w1102_,
		_w6412_
	);
	LUT3 #(
		.INIT('h70)
	) name6379 (
		_w1202_,
		_w1233_,
		_w5524_,
		_w6413_
	);
	LUT3 #(
		.INIT('h01)
	) name6380 (
		_w6412_,
		_w6413_,
		_w6411_,
		_w6414_
	);
	LUT4 #(
		.INIT('h6f00)
	) name6381 (
		_w2335_,
		_w2337_,
		_w35_,
		_w6414_,
		_w6415_
	);
	LUT2 #(
		.INIT('h6)
	) name6382 (
		\a[5] ,
		_w6415_,
		_w6416_
	);
	LUT4 #(
		.INIT('h54ab)
	) name6383 (
		_w6128_,
		_w6296_,
		_w6297_,
		_w6299_,
		_w6417_
	);
	LUT2 #(
		.INIT('h4)
	) name6384 (
		_w6416_,
		_w6417_,
		_w6418_
	);
	LUT3 #(
		.INIT('h70)
	) name6385 (
		_w1202_,
		_w1233_,
		_w6031_,
		_w6419_
	);
	LUT3 #(
		.INIT('h70)
	) name6386 (
		_w1253_,
		_w1294_,
		_w5524_,
		_w6420_
	);
	LUT3 #(
		.INIT('h2a)
	) name6387 (
		_w6324_,
		_w1136_,
		_w1187_,
		_w6421_
	);
	LUT3 #(
		.INIT('h01)
	) name6388 (
		_w6420_,
		_w6421_,
		_w6419_,
		_w6422_
	);
	LUT4 #(
		.INIT('h95aa)
	) name6389 (
		\a[5] ,
		_w3067_,
		_w35_,
		_w6422_,
		_w6423_
	);
	LUT3 #(
		.INIT('h09)
	) name6390 (
		_w6296_,
		_w6298_,
		_w6423_,
		_w6424_
	);
	LUT3 #(
		.INIT('h2a)
	) name6391 (
		_w6324_,
		_w1202_,
		_w1233_,
		_w6425_
	);
	LUT3 #(
		.INIT('h70)
	) name6392 (
		_w1325_,
		_w1367_,
		_w5524_,
		_w6426_
	);
	LUT3 #(
		.INIT('h70)
	) name6393 (
		_w1253_,
		_w1294_,
		_w6031_,
		_w6427_
	);
	LUT3 #(
		.INIT('h01)
	) name6394 (
		_w6426_,
		_w6427_,
		_w6425_,
		_w6428_
	);
	LUT4 #(
		.INIT('h6f00)
	) name6395 (
		_w2331_,
		_w2333_,
		_w35_,
		_w6428_,
		_w6429_
	);
	LUT2 #(
		.INIT('h6)
	) name6396 (
		\a[5] ,
		_w6429_,
		_w6430_
	);
	LUT4 #(
		.INIT('h001e)
	) name6397 (
		_w6142_,
		_w6294_,
		_w6295_,
		_w6430_,
		_w6431_
	);
	LUT4 #(
		.INIT('h54ab)
	) name6398 (
		_w6148_,
		_w6290_,
		_w6291_,
		_w6293_,
		_w6432_
	);
	LUT3 #(
		.INIT('h70)
	) name6399 (
		_w1381_,
		_w1398_,
		_w5524_,
		_w6433_
	);
	LUT3 #(
		.INIT('h70)
	) name6400 (
		_w1325_,
		_w1367_,
		_w6031_,
		_w6434_
	);
	LUT3 #(
		.INIT('h2a)
	) name6401 (
		_w6324_,
		_w1253_,
		_w1294_,
		_w6435_
	);
	LUT3 #(
		.INIT('h01)
	) name6402 (
		_w6434_,
		_w6435_,
		_w6433_,
		_w6436_
	);
	LUT4 #(
		.INIT('h95aa)
	) name6403 (
		\a[5] ,
		_w3182_,
		_w35_,
		_w6436_,
		_w6437_
	);
	LUT2 #(
		.INIT('h2)
	) name6404 (
		_w6432_,
		_w6437_,
		_w6438_
	);
	LUT2 #(
		.INIT('h9)
	) name6405 (
		_w6290_,
		_w6292_,
		_w6439_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6406 (
		_w1454_,
		_w1426_,
		_w1478_,
		_w5524_,
		_w6440_
	);
	LUT3 #(
		.INIT('h2a)
	) name6407 (
		_w6324_,
		_w1325_,
		_w1367_,
		_w6441_
	);
	LUT3 #(
		.INIT('h70)
	) name6408 (
		_w1381_,
		_w1398_,
		_w6031_,
		_w6442_
	);
	LUT3 #(
		.INIT('h01)
	) name6409 (
		_w6441_,
		_w6442_,
		_w6440_,
		_w6443_
	);
	LUT4 #(
		.INIT('h6f00)
	) name6410 (
		_w2327_,
		_w2329_,
		_w35_,
		_w6443_,
		_w6444_
	);
	LUT2 #(
		.INIT('h6)
	) name6411 (
		\a[5] ,
		_w6444_,
		_w6445_
	);
	LUT3 #(
		.INIT('h09)
	) name6412 (
		_w6290_,
		_w6292_,
		_w6445_,
		_w6446_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6413 (
		_w1454_,
		_w1426_,
		_w1478_,
		_w6031_,
		_w6447_
	);
	LUT3 #(
		.INIT('h2a)
	) name6414 (
		_w6324_,
		_w1381_,
		_w1398_,
		_w6448_
	);
	LUT3 #(
		.INIT('h70)
	) name6415 (
		_w1501_,
		_w1545_,
		_w5524_,
		_w6449_
	);
	LUT3 #(
		.INIT('h01)
	) name6416 (
		_w6448_,
		_w6449_,
		_w6447_,
		_w6450_
	);
	LUT4 #(
		.INIT('h95aa)
	) name6417 (
		\a[5] ,
		_w3362_,
		_w35_,
		_w6450_,
		_w6451_
	);
	LUT4 #(
		.INIT('h001e)
	) name6418 (
		_w6162_,
		_w6288_,
		_w6289_,
		_w6451_,
		_w6452_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name6419 (
		_w6324_,
		_w1454_,
		_w1426_,
		_w1478_,
		_w6453_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6420 (
		_w1584_,
		_w1569_,
		_w1606_,
		_w5524_,
		_w6454_
	);
	LUT3 #(
		.INIT('h70)
	) name6421 (
		_w1501_,
		_w1545_,
		_w6031_,
		_w6455_
	);
	LUT3 #(
		.INIT('h01)
	) name6422 (
		_w6454_,
		_w6455_,
		_w6453_,
		_w6456_
	);
	LUT4 #(
		.INIT('h6f00)
	) name6423 (
		_w2323_,
		_w2325_,
		_w35_,
		_w6456_,
		_w6457_
	);
	LUT2 #(
		.INIT('h6)
	) name6424 (
		\a[5] ,
		_w6457_,
		_w6458_
	);
	LUT4 #(
		.INIT('h54ab)
	) name6425 (
		_w6170_,
		_w6284_,
		_w6285_,
		_w6287_,
		_w6459_
	);
	LUT2 #(
		.INIT('h4)
	) name6426 (
		_w6458_,
		_w6459_,
		_w6460_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6427 (
		_w1584_,
		_w1569_,
		_w1606_,
		_w6031_,
		_w6461_
	);
	LUT3 #(
		.INIT('h2a)
	) name6428 (
		_w6324_,
		_w1501_,
		_w1545_,
		_w6462_
	);
	LUT3 #(
		.INIT('h70)
	) name6429 (
		_w1620_,
		_w1661_,
		_w5524_,
		_w6463_
	);
	LUT3 #(
		.INIT('h01)
	) name6430 (
		_w6461_,
		_w6462_,
		_w6463_,
		_w6464_
	);
	LUT4 #(
		.INIT('h95aa)
	) name6431 (
		\a[5] ,
		_w3495_,
		_w35_,
		_w6464_,
		_w6465_
	);
	LUT3 #(
		.INIT('h09)
	) name6432 (
		_w6284_,
		_w6286_,
		_w6465_,
		_w6466_
	);
	LUT3 #(
		.INIT('h70)
	) name6433 (
		_w1692_,
		_w1723_,
		_w5524_,
		_w6467_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name6434 (
		_w6324_,
		_w1584_,
		_w1569_,
		_w1606_,
		_w6468_
	);
	LUT3 #(
		.INIT('h70)
	) name6435 (
		_w1620_,
		_w1661_,
		_w6031_,
		_w6469_
	);
	LUT3 #(
		.INIT('h01)
	) name6436 (
		_w6468_,
		_w6469_,
		_w6467_,
		_w6470_
	);
	LUT4 #(
		.INIT('h6f00)
	) name6437 (
		_w2319_,
		_w2321_,
		_w35_,
		_w6470_,
		_w6471_
	);
	LUT2 #(
		.INIT('h6)
	) name6438 (
		\a[5] ,
		_w6471_,
		_w6472_
	);
	LUT4 #(
		.INIT('h001e)
	) name6439 (
		_w6184_,
		_w6282_,
		_w6283_,
		_w6472_,
		_w6473_
	);
	LUT4 #(
		.INIT('h54ab)
	) name6440 (
		_w6190_,
		_w6278_,
		_w6279_,
		_w6281_,
		_w6474_
	);
	LUT3 #(
		.INIT('h70)
	) name6441 (
		_w1692_,
		_w1723_,
		_w6031_,
		_w6475_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6442 (
		_w1751_,
		_w1742_,
		_w1771_,
		_w5524_,
		_w6476_
	);
	LUT3 #(
		.INIT('h2a)
	) name6443 (
		_w6324_,
		_w1620_,
		_w1661_,
		_w6477_
	);
	LUT3 #(
		.INIT('h01)
	) name6444 (
		_w6476_,
		_w6477_,
		_w6475_,
		_w6478_
	);
	LUT4 #(
		.INIT('h95aa)
	) name6445 (
		\a[5] ,
		_w3599_,
		_w35_,
		_w6478_,
		_w6479_
	);
	LUT2 #(
		.INIT('h2)
	) name6446 (
		_w6474_,
		_w6479_,
		_w6480_
	);
	LUT2 #(
		.INIT('h9)
	) name6447 (
		_w6278_,
		_w6280_,
		_w6481_
	);
	LUT3 #(
		.INIT('h2a)
	) name6448 (
		_w6324_,
		_w1692_,
		_w1723_,
		_w6482_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6449 (
		_w1751_,
		_w1742_,
		_w1771_,
		_w6031_,
		_w6483_
	);
	LUT3 #(
		.INIT('h70)
	) name6450 (
		_w1795_,
		_w1796_,
		_w5524_,
		_w6484_
	);
	LUT3 #(
		.INIT('h01)
	) name6451 (
		_w6483_,
		_w6484_,
		_w6482_,
		_w6485_
	);
	LUT4 #(
		.INIT('h6f00)
	) name6452 (
		_w2315_,
		_w2317_,
		_w35_,
		_w6485_,
		_w6486_
	);
	LUT2 #(
		.INIT('h6)
	) name6453 (
		\a[5] ,
		_w6486_,
		_w6487_
	);
	LUT3 #(
		.INIT('h09)
	) name6454 (
		_w6278_,
		_w6280_,
		_w6487_,
		_w6488_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name6455 (
		_w6324_,
		_w1751_,
		_w1742_,
		_w1771_,
		_w6489_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6456 (
		_w1817_,
		_w1799_,
		_w1840_,
		_w5524_,
		_w6490_
	);
	LUT3 #(
		.INIT('h70)
	) name6457 (
		_w1795_,
		_w1796_,
		_w6031_,
		_w6491_
	);
	LUT3 #(
		.INIT('h01)
	) name6458 (
		_w6490_,
		_w6491_,
		_w6489_,
		_w6492_
	);
	LUT4 #(
		.INIT('h95aa)
	) name6459 (
		\a[5] ,
		_w3909_,
		_w35_,
		_w6492_,
		_w6493_
	);
	LUT4 #(
		.INIT('h001e)
	) name6460 (
		_w6205_,
		_w6275_,
		_w6277_,
		_w6493_,
		_w6494_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6461 (
		_w1817_,
		_w1799_,
		_w1840_,
		_w6031_,
		_w6495_
	);
	LUT3 #(
		.INIT('h2a)
	) name6462 (
		_w6324_,
		_w1795_,
		_w1796_,
		_w6496_
	);
	LUT3 #(
		.INIT('h70)
	) name6463 (
		_w1863_,
		_w1875_,
		_w5524_,
		_w6497_
	);
	LUT3 #(
		.INIT('h01)
	) name6464 (
		_w6496_,
		_w6497_,
		_w6495_,
		_w6498_
	);
	LUT4 #(
		.INIT('h6f00)
	) name6465 (
		_w2311_,
		_w2313_,
		_w35_,
		_w6498_,
		_w6499_
	);
	LUT2 #(
		.INIT('h6)
	) name6466 (
		\a[5] ,
		_w6499_,
		_w6500_
	);
	LUT4 #(
		.INIT('h54ab)
	) name6467 (
		_w6213_,
		_w6271_,
		_w6272_,
		_w6274_,
		_w6501_
	);
	LUT2 #(
		.INIT('h4)
	) name6468 (
		_w6500_,
		_w6501_,
		_w6502_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name6469 (
		_w6324_,
		_w1817_,
		_w1799_,
		_w1840_,
		_w6503_
	);
	LUT3 #(
		.INIT('h70)
	) name6470 (
		_w1898_,
		_w1928_,
		_w5524_,
		_w6504_
	);
	LUT3 #(
		.INIT('h70)
	) name6471 (
		_w1863_,
		_w1875_,
		_w6031_,
		_w6505_
	);
	LUT3 #(
		.INIT('h01)
	) name6472 (
		_w6504_,
		_w6505_,
		_w6503_,
		_w6506_
	);
	LUT4 #(
		.INIT('h95aa)
	) name6473 (
		\a[5] ,
		_w3972_,
		_w35_,
		_w6506_,
		_w6507_
	);
	LUT3 #(
		.INIT('h09)
	) name6474 (
		_w6271_,
		_w6273_,
		_w6507_,
		_w6508_
	);
	LUT3 #(
		.INIT('h1e)
	) name6475 (
		_w6227_,
		_w6268_,
		_w6270_,
		_w6509_
	);
	LUT3 #(
		.INIT('h70)
	) name6476 (
		_w1501_,
		_w1949_,
		_w5524_,
		_w6510_
	);
	LUT3 #(
		.INIT('h70)
	) name6477 (
		_w1898_,
		_w1928_,
		_w6031_,
		_w6511_
	);
	LUT3 #(
		.INIT('h2a)
	) name6478 (
		_w6324_,
		_w1863_,
		_w1875_,
		_w6512_
	);
	LUT3 #(
		.INIT('h01)
	) name6479 (
		_w6511_,
		_w6512_,
		_w6510_,
		_w6513_
	);
	LUT4 #(
		.INIT('h6f00)
	) name6480 (
		_w2307_,
		_w2309_,
		_w35_,
		_w6513_,
		_w6514_
	);
	LUT2 #(
		.INIT('h6)
	) name6481 (
		\a[5] ,
		_w6514_,
		_w6515_
	);
	LUT2 #(
		.INIT('h2)
	) name6482 (
		_w6509_,
		_w6515_,
		_w6516_
	);
	LUT4 #(
		.INIT('h54ab)
	) name6483 (
		_w6235_,
		_w6264_,
		_w6265_,
		_w6267_,
		_w6517_
	);
	LUT3 #(
		.INIT('h70)
	) name6484 (
		_w1973_,
		_w1997_,
		_w5524_,
		_w6518_
	);
	LUT3 #(
		.INIT('h2a)
	) name6485 (
		_w6324_,
		_w1898_,
		_w1928_,
		_w6519_
	);
	LUT3 #(
		.INIT('h70)
	) name6486 (
		_w1501_,
		_w1949_,
		_w6031_,
		_w6520_
	);
	LUT3 #(
		.INIT('h01)
	) name6487 (
		_w6519_,
		_w6520_,
		_w6518_,
		_w6521_
	);
	LUT4 #(
		.INIT('h95aa)
	) name6488 (
		\a[5] ,
		_w4126_,
		_w35_,
		_w6521_,
		_w6522_
	);
	LUT2 #(
		.INIT('h2)
	) name6489 (
		_w6517_,
		_w6522_,
		_w6523_
	);
	LUT2 #(
		.INIT('h9)
	) name6490 (
		_w6264_,
		_w6266_,
		_w6524_
	);
	LUT3 #(
		.INIT('h70)
	) name6491 (
		_w1973_,
		_w1997_,
		_w6031_,
		_w6525_
	);
	LUT3 #(
		.INIT('h2a)
	) name6492 (
		_w6324_,
		_w1501_,
		_w1949_,
		_w6526_
	);
	LUT3 #(
		.INIT('h70)
	) name6493 (
		_w2023_,
		_w2055_,
		_w5524_,
		_w6527_
	);
	LUT3 #(
		.INIT('h01)
	) name6494 (
		_w6526_,
		_w6527_,
		_w6525_,
		_w6528_
	);
	LUT4 #(
		.INIT('h6f00)
	) name6495 (
		_w2303_,
		_w2305_,
		_w35_,
		_w6528_,
		_w6529_
	);
	LUT2 #(
		.INIT('h6)
	) name6496 (
		\a[5] ,
		_w6529_,
		_w6530_
	);
	LUT4 #(
		.INIT('h8241)
	) name6497 (
		\a[5] ,
		_w6264_,
		_w6266_,
		_w6529_,
		_w6531_
	);
	LUT3 #(
		.INIT('h2a)
	) name6498 (
		_w6324_,
		_w1973_,
		_w1997_,
		_w6532_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6499 (
		_w1874_,
		_w2076_,
		_w2099_,
		_w5524_,
		_w6533_
	);
	LUT3 #(
		.INIT('h70)
	) name6500 (
		_w2023_,
		_w2055_,
		_w6031_,
		_w6534_
	);
	LUT3 #(
		.INIT('h01)
	) name6501 (
		_w6533_,
		_w6534_,
		_w6532_,
		_w6535_
	);
	LUT4 #(
		.INIT('h95aa)
	) name6502 (
		\a[5] ,
		_w4151_,
		_w35_,
		_w6535_,
		_w6536_
	);
	LUT2 #(
		.INIT('h9)
	) name6503 (
		_w6261_,
		_w6263_,
		_w6537_
	);
	LUT2 #(
		.INIT('h4)
	) name6504 (
		_w6536_,
		_w6537_,
		_w6538_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6505 (
		_w1874_,
		_w2076_,
		_w2099_,
		_w6031_,
		_w6539_
	);
	LUT3 #(
		.INIT('h70)
	) name6506 (
		_w2124_,
		_w2133_,
		_w5524_,
		_w6540_
	);
	LUT3 #(
		.INIT('h2a)
	) name6507 (
		_w6324_,
		_w2023_,
		_w2055_,
		_w6541_
	);
	LUT3 #(
		.INIT('h01)
	) name6508 (
		_w6539_,
		_w6540_,
		_w6541_,
		_w6542_
	);
	LUT4 #(
		.INIT('h6f00)
	) name6509 (
		_w2299_,
		_w2301_,
		_w35_,
		_w6542_,
		_w6543_
	);
	LUT3 #(
		.INIT('h69)
	) name6510 (
		_w5953_,
		_w6255_,
		_w6260_,
		_w6544_
	);
	LUT3 #(
		.INIT('h90)
	) name6511 (
		\a[5] ,
		_w6543_,
		_w6544_,
		_w6545_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name6512 (
		_w6324_,
		_w1874_,
		_w2076_,
		_w2099_,
		_w6546_
	);
	LUT3 #(
		.INIT('h70)
	) name6513 (
		_w2124_,
		_w2133_,
		_w6031_,
		_w6547_
	);
	LUT3 #(
		.INIT('h70)
	) name6514 (
		_w2155_,
		_w2156_,
		_w5524_,
		_w6548_
	);
	LUT3 #(
		.INIT('h01)
	) name6515 (
		_w6546_,
		_w6547_,
		_w6548_,
		_w6549_
	);
	LUT4 #(
		.INIT('h95aa)
	) name6516 (
		\a[5] ,
		_w4209_,
		_w35_,
		_w6549_,
		_w6550_
	);
	LUT3 #(
		.INIT('h8a)
	) name6517 (
		\a[8] ,
		_w6247_,
		_w6246_,
		_w6551_
	);
	LUT2 #(
		.INIT('h9)
	) name6518 (
		_w6254_,
		_w6551_,
		_w6552_
	);
	LUT2 #(
		.INIT('h4)
	) name6519 (
		_w6550_,
		_w6552_,
		_w6553_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6520 (
		_w2193_,
		_w2183_,
		_w2213_,
		_w5524_,
		_w6554_
	);
	LUT3 #(
		.INIT('h70)
	) name6521 (
		_w2155_,
		_w2156_,
		_w6031_,
		_w6555_
	);
	LUT3 #(
		.INIT('h2a)
	) name6522 (
		_w6324_,
		_w2124_,
		_w2133_,
		_w6556_
	);
	LUT3 #(
		.INIT('h01)
	) name6523 (
		_w6554_,
		_w6555_,
		_w6556_,
		_w6557_
	);
	LUT4 #(
		.INIT('h6f00)
	) name6524 (
		_w2295_,
		_w2297_,
		_w35_,
		_w6557_,
		_w6558_
	);
	LUT4 #(
		.INIT('h002a)
	) name6525 (
		\a[8] ,
		_w2228_,
		_w2262_,
		_w4874_,
		_w6559_
	);
	LUT2 #(
		.INIT('h9)
	) name6526 (
		_w6246_,
		_w6559_,
		_w6560_
	);
	LUT3 #(
		.INIT('h90)
	) name6527 (
		\a[5] ,
		_w6558_,
		_w6560_,
		_w6561_
	);
	LUT3 #(
		.INIT('h70)
	) name6528 (
		_w2228_,
		_w2262_,
		_w6031_,
		_w6562_
	);
	LUT3 #(
		.INIT('h2a)
	) name6529 (
		_w6324_,
		_w2273_,
		_w2293_,
		_w6563_
	);
	LUT4 #(
		.INIT('h000b)
	) name6530 (
		_w4599_,
		_w35_,
		_w6562_,
		_w6563_,
		_w6564_
	);
	LUT3 #(
		.INIT('h15)
	) name6531 (
		_w34_,
		_w2228_,
		_w2262_,
		_w6565_
	);
	LUT4 #(
		.INIT('ha888)
	) name6532 (
		\a[5] ,
		_w34_,
		_w2228_,
		_w2262_,
		_w6566_
	);
	LUT3 #(
		.INIT('h90)
	) name6533 (
		_w2214_,
		_w4258_,
		_w35_,
		_w6567_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name6534 (
		_w6324_,
		_w2193_,
		_w2183_,
		_w2213_,
		_w6568_
	);
	LUT3 #(
		.INIT('h70)
	) name6535 (
		_w2228_,
		_w2262_,
		_w5524_,
		_w6569_
	);
	LUT3 #(
		.INIT('h70)
	) name6536 (
		_w2273_,
		_w2293_,
		_w6031_,
		_w6570_
	);
	LUT3 #(
		.INIT('h01)
	) name6537 (
		_w6569_,
		_w6570_,
		_w6568_,
		_w6571_
	);
	LUT2 #(
		.INIT('h4)
	) name6538 (
		_w6567_,
		_w6571_,
		_w6572_
	);
	LUT4 #(
		.INIT('h0800)
	) name6539 (
		_w6564_,
		_w6566_,
		_w6567_,
		_w6571_,
		_w6573_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6540 (
		_w2193_,
		_w2183_,
		_w2213_,
		_w6031_,
		_w6574_
	);
	LUT3 #(
		.INIT('h2a)
	) name6541 (
		_w6324_,
		_w2155_,
		_w2156_,
		_w6575_
	);
	LUT3 #(
		.INIT('h70)
	) name6542 (
		_w2273_,
		_w2293_,
		_w5524_,
		_w6576_
	);
	LUT3 #(
		.INIT('h01)
	) name6543 (
		_w6574_,
		_w6575_,
		_w6576_,
		_w6577_
	);
	LUT4 #(
		.INIT('h95aa)
	) name6544 (
		\a[5] ,
		_w4293_,
		_w35_,
		_w6577_,
		_w6578_
	);
	LUT3 #(
		.INIT('h71)
	) name6545 (
		_w6247_,
		_w6573_,
		_w6578_,
		_w6579_
	);
	LUT3 #(
		.INIT('h06)
	) name6546 (
		\a[5] ,
		_w6558_,
		_w6560_,
		_w6580_
	);
	LUT3 #(
		.INIT('h69)
	) name6547 (
		\a[5] ,
		_w6558_,
		_w6560_,
		_w6581_
	);
	LUT3 #(
		.INIT('h54)
	) name6548 (
		_w6561_,
		_w6579_,
		_w6580_,
		_w6582_
	);
	LUT2 #(
		.INIT('h2)
	) name6549 (
		_w6550_,
		_w6552_,
		_w6583_
	);
	LUT2 #(
		.INIT('h9)
	) name6550 (
		_w6550_,
		_w6552_,
		_w6584_
	);
	LUT3 #(
		.INIT('h69)
	) name6551 (
		\a[5] ,
		_w6543_,
		_w6544_,
		_w6585_
	);
	LUT4 #(
		.INIT('h4d00)
	) name6552 (
		_w6550_,
		_w6552_,
		_w6582_,
		_w6585_,
		_w6586_
	);
	LUT2 #(
		.INIT('h2)
	) name6553 (
		_w6536_,
		_w6537_,
		_w6587_
	);
	LUT2 #(
		.INIT('h9)
	) name6554 (
		_w6536_,
		_w6537_,
		_w6588_
	);
	LUT4 #(
		.INIT('h5501)
	) name6555 (
		_w6538_,
		_w6545_,
		_w6586_,
		_w6587_,
		_w6589_
	);
	LUT4 #(
		.INIT('h1428)
	) name6556 (
		\a[5] ,
		_w6264_,
		_w6266_,
		_w6529_,
		_w6590_
	);
	LUT4 #(
		.INIT('h6996)
	) name6557 (
		\a[5] ,
		_w6264_,
		_w6266_,
		_w6529_,
		_w6591_
	);
	LUT2 #(
		.INIT('h9)
	) name6558 (
		_w6517_,
		_w6522_,
		_w6592_
	);
	LUT4 #(
		.INIT('h2b00)
	) name6559 (
		_w6524_,
		_w6530_,
		_w6589_,
		_w6592_,
		_w6593_
	);
	LUT2 #(
		.INIT('h4)
	) name6560 (
		_w6509_,
		_w6515_,
		_w6594_
	);
	LUT2 #(
		.INIT('h9)
	) name6561 (
		_w6509_,
		_w6515_,
		_w6595_
	);
	LUT4 #(
		.INIT('h5501)
	) name6562 (
		_w6516_,
		_w6523_,
		_w6593_,
		_w6594_,
		_w6596_
	);
	LUT3 #(
		.INIT('h60)
	) name6563 (
		_w6271_,
		_w6273_,
		_w6507_,
		_w6597_
	);
	LUT3 #(
		.INIT('h96)
	) name6564 (
		_w6271_,
		_w6273_,
		_w6507_,
		_w6598_
	);
	LUT2 #(
		.INIT('h9)
	) name6565 (
		_w6500_,
		_w6501_,
		_w6599_
	);
	LUT4 #(
		.INIT('hba00)
	) name6566 (
		_w6508_,
		_w6596_,
		_w6598_,
		_w6599_,
		_w6600_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name6567 (
		_w6205_,
		_w6275_,
		_w6277_,
		_w6493_,
		_w6601_
	);
	LUT4 #(
		.INIT('h0155)
	) name6568 (
		_w6494_,
		_w6502_,
		_w6600_,
		_w6601_,
		_w6602_
	);
	LUT3 #(
		.INIT('h60)
	) name6569 (
		_w6278_,
		_w6280_,
		_w6487_,
		_w6603_
	);
	LUT3 #(
		.INIT('h96)
	) name6570 (
		_w6278_,
		_w6280_,
		_w6487_,
		_w6604_
	);
	LUT2 #(
		.INIT('h9)
	) name6571 (
		_w6474_,
		_w6479_,
		_w6605_
	);
	LUT4 #(
		.INIT('h2b00)
	) name6572 (
		_w6481_,
		_w6487_,
		_w6602_,
		_w6605_,
		_w6606_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name6573 (
		_w6184_,
		_w6282_,
		_w6283_,
		_w6472_,
		_w6607_
	);
	LUT4 #(
		.INIT('h0155)
	) name6574 (
		_w6473_,
		_w6480_,
		_w6606_,
		_w6607_,
		_w6608_
	);
	LUT3 #(
		.INIT('h60)
	) name6575 (
		_w6284_,
		_w6286_,
		_w6465_,
		_w6609_
	);
	LUT3 #(
		.INIT('h96)
	) name6576 (
		_w6284_,
		_w6286_,
		_w6465_,
		_w6610_
	);
	LUT2 #(
		.INIT('h9)
	) name6577 (
		_w6458_,
		_w6459_,
		_w6611_
	);
	LUT4 #(
		.INIT('hba00)
	) name6578 (
		_w6466_,
		_w6608_,
		_w6610_,
		_w6611_,
		_w6612_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name6579 (
		_w6162_,
		_w6288_,
		_w6289_,
		_w6451_,
		_w6613_
	);
	LUT4 #(
		.INIT('h0155)
	) name6580 (
		_w6452_,
		_w6460_,
		_w6612_,
		_w6613_,
		_w6614_
	);
	LUT3 #(
		.INIT('h60)
	) name6581 (
		_w6290_,
		_w6292_,
		_w6445_,
		_w6615_
	);
	LUT3 #(
		.INIT('h96)
	) name6582 (
		_w6290_,
		_w6292_,
		_w6445_,
		_w6616_
	);
	LUT2 #(
		.INIT('h9)
	) name6583 (
		_w6432_,
		_w6437_,
		_w6617_
	);
	LUT4 #(
		.INIT('h2b00)
	) name6584 (
		_w6439_,
		_w6445_,
		_w6614_,
		_w6617_,
		_w6618_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name6585 (
		_w6142_,
		_w6294_,
		_w6295_,
		_w6430_,
		_w6619_
	);
	LUT4 #(
		.INIT('h0155)
	) name6586 (
		_w6431_,
		_w6438_,
		_w6618_,
		_w6619_,
		_w6620_
	);
	LUT3 #(
		.INIT('h60)
	) name6587 (
		_w6296_,
		_w6298_,
		_w6423_,
		_w6621_
	);
	LUT3 #(
		.INIT('h96)
	) name6588 (
		_w6296_,
		_w6298_,
		_w6423_,
		_w6622_
	);
	LUT2 #(
		.INIT('h9)
	) name6589 (
		_w6416_,
		_w6417_,
		_w6623_
	);
	LUT4 #(
		.INIT('hba00)
	) name6590 (
		_w6424_,
		_w6620_,
		_w6622_,
		_w6623_,
		_w6624_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name6591 (
		_w6120_,
		_w6300_,
		_w6301_,
		_w6409_,
		_w6625_
	);
	LUT4 #(
		.INIT('h0155)
	) name6592 (
		_w6410_,
		_w6418_,
		_w6624_,
		_w6625_,
		_w6626_
	);
	LUT3 #(
		.INIT('h60)
	) name6593 (
		_w6302_,
		_w6304_,
		_w6403_,
		_w6627_
	);
	LUT3 #(
		.INIT('h96)
	) name6594 (
		_w6302_,
		_w6304_,
		_w6403_,
		_w6628_
	);
	LUT2 #(
		.INIT('h9)
	) name6595 (
		_w6390_,
		_w6395_,
		_w6629_
	);
	LUT4 #(
		.INIT('h2b00)
	) name6596 (
		_w6397_,
		_w6403_,
		_w6626_,
		_w6629_,
		_w6630_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name6597 (
		_w6100_,
		_w6306_,
		_w6307_,
		_w6388_,
		_w6631_
	);
	LUT4 #(
		.INIT('h0155)
	) name6598 (
		_w6389_,
		_w6396_,
		_w6630_,
		_w6631_,
		_w6632_
	);
	LUT3 #(
		.INIT('h60)
	) name6599 (
		_w6308_,
		_w6310_,
		_w6381_,
		_w6633_
	);
	LUT3 #(
		.INIT('h96)
	) name6600 (
		_w6308_,
		_w6310_,
		_w6381_,
		_w6634_
	);
	LUT2 #(
		.INIT('h9)
	) name6601 (
		_w6374_,
		_w6375_,
		_w6635_
	);
	LUT4 #(
		.INIT('hba00)
	) name6602 (
		_w6382_,
		_w6632_,
		_w6634_,
		_w6635_,
		_w6636_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name6603 (
		_w6078_,
		_w6312_,
		_w6313_,
		_w6367_,
		_w6637_
	);
	LUT4 #(
		.INIT('h0155)
	) name6604 (
		_w6368_,
		_w6376_,
		_w6636_,
		_w6637_,
		_w6638_
	);
	LUT3 #(
		.INIT('h60)
	) name6605 (
		_w6314_,
		_w6316_,
		_w6360_,
		_w6639_
	);
	LUT3 #(
		.INIT('h96)
	) name6606 (
		_w6314_,
		_w6316_,
		_w6360_,
		_w6640_
	);
	LUT2 #(
		.INIT('h9)
	) name6607 (
		_w6352_,
		_w6353_,
		_w6641_
	);
	LUT4 #(
		.INIT('h4d00)
	) name6608 (
		_w6360_,
		_w6361_,
		_w6638_,
		_w6641_,
		_w6642_
	);
	LUT3 #(
		.INIT('h69)
	) name6609 (
		\a[2] ,
		_w6336_,
		_w6342_,
		_w6643_
	);
	LUT4 #(
		.INIT('he11e)
	) name6610 (
		_w6058_,
		_w6318_,
		_w6319_,
		_w6643_,
		_w6644_
	);
	LUT3 #(
		.INIT('he0)
	) name6611 (
		_w6354_,
		_w6642_,
		_w6644_,
		_w6645_
	);
	LUT3 #(
		.INIT('h1e)
	) name6612 (
		_w6354_,
		_w6642_,
		_w6644_,
		_w6646_
	);
	LUT4 #(
		.INIT('h54ab)
	) name6613 (
		_w6362_,
		_w6638_,
		_w6639_,
		_w6641_,
		_w6647_
	);
	LUT4 #(
		.INIT('hf400)
	) name6614 (
		_w374_,
		_w2361_,
		_w2404_,
		_w6335_,
		_w6648_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6615 (
		_w121_,
		_w418_,
		_w422_,
		_w6334_,
		_w6649_
	);
	LUT2 #(
		.INIT('h4)
	) name6616 (
		\a[0] ,
		\a[1] ,
		_w6650_
	);
	LUT3 #(
		.INIT('h70)
	) name6617 (
		_w352_,
		_w373_,
		_w6650_,
		_w6651_
	);
	LUT2 #(
		.INIT('h1)
	) name6618 (
		_w6649_,
		_w6651_,
		_w6652_
	);
	LUT3 #(
		.INIT('h9a)
	) name6619 (
		\a[2] ,
		_w6648_,
		_w6652_,
		_w6653_
	);
	LUT2 #(
		.INIT('h2)
	) name6620 (
		_w6647_,
		_w6653_,
		_w6654_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6621 (
		_w486_,
		_w487_,
		_w509_,
		_w6334_,
		_w6655_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6622 (
		_w121_,
		_w418_,
		_w422_,
		_w6650_,
		_w6656_
	);
	LUT3 #(
		.INIT('h82)
	) name6623 (
		\a[0] ,
		\a[1] ,
		\a[2] ,
		_w6657_
	);
	LUT3 #(
		.INIT('h70)
	) name6624 (
		_w352_,
		_w373_,
		_w6657_,
		_w6658_
	);
	LUT3 #(
		.INIT('h01)
	) name6625 (
		_w6655_,
		_w6656_,
		_w6658_,
		_w6659_
	);
	LUT4 #(
		.INIT('h95aa)
	) name6626 (
		\a[2] ,
		_w2535_,
		_w6335_,
		_w6659_,
		_w6660_
	);
	LUT3 #(
		.INIT('h09)
	) name6627 (
		_w6638_,
		_w6640_,
		_w6660_,
		_w6661_
	);
	LUT3 #(
		.INIT('h1e)
	) name6628 (
		_w6376_,
		_w6636_,
		_w6637_,
		_w6662_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6629 (
		_w486_,
		_w487_,
		_w509_,
		_w6650_,
		_w6663_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6630 (
		_w121_,
		_w418_,
		_w422_,
		_w6657_,
		_w6664_
	);
	LUT3 #(
		.INIT('h70)
	) name6631 (
		_w544_,
		_w558_,
		_w6334_,
		_w6665_
	);
	LUT3 #(
		.INIT('h01)
	) name6632 (
		_w6663_,
		_w6664_,
		_w6665_,
		_w6666_
	);
	LUT4 #(
		.INIT('h6f00)
	) name6633 (
		_w2355_,
		_w2357_,
		_w6335_,
		_w6666_,
		_w6667_
	);
	LUT2 #(
		.INIT('h6)
	) name6634 (
		\a[2] ,
		_w6667_,
		_w6668_
	);
	LUT4 #(
		.INIT('h001e)
	) name6635 (
		_w6376_,
		_w6636_,
		_w6637_,
		_w6668_,
		_w6669_
	);
	LUT4 #(
		.INIT('h54ab)
	) name6636 (
		_w6382_,
		_w6632_,
		_w6633_,
		_w6635_,
		_w6670_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6637 (
		_w486_,
		_w487_,
		_w509_,
		_w6657_,
		_w6671_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6638 (
		_w587_,
		_w608_,
		_w624_,
		_w6334_,
		_w6672_
	);
	LUT3 #(
		.INIT('h70)
	) name6639 (
		_w544_,
		_w558_,
		_w6650_,
		_w6673_
	);
	LUT3 #(
		.INIT('h01)
	) name6640 (
		_w6671_,
		_w6672_,
		_w6673_,
		_w6674_
	);
	LUT4 #(
		.INIT('h95aa)
	) name6641 (
		\a[2] ,
		_w2526_,
		_w6335_,
		_w6674_,
		_w6675_
	);
	LUT2 #(
		.INIT('h2)
	) name6642 (
		_w6670_,
		_w6675_,
		_w6676_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6643 (
		_w587_,
		_w608_,
		_w624_,
		_w6650_,
		_w6677_
	);
	LUT3 #(
		.INIT('h70)
	) name6644 (
		_w666_,
		_w694_,
		_w6334_,
		_w6678_
	);
	LUT3 #(
		.INIT('h70)
	) name6645 (
		_w544_,
		_w558_,
		_w6657_,
		_w6679_
	);
	LUT3 #(
		.INIT('h01)
	) name6646 (
		_w6678_,
		_w6679_,
		_w6677_,
		_w6680_
	);
	LUT4 #(
		.INIT('h6f00)
	) name6647 (
		_w2351_,
		_w2353_,
		_w6335_,
		_w6680_,
		_w6681_
	);
	LUT2 #(
		.INIT('h6)
	) name6648 (
		\a[2] ,
		_w6681_,
		_w6682_
	);
	LUT3 #(
		.INIT('h09)
	) name6649 (
		_w6632_,
		_w6634_,
		_w6682_,
		_w6683_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6650 (
		_w587_,
		_w608_,
		_w624_,
		_w6657_,
		_w6684_
	);
	LUT3 #(
		.INIT('h70)
	) name6651 (
		_w725_,
		_w764_,
		_w6334_,
		_w6685_
	);
	LUT3 #(
		.INIT('h70)
	) name6652 (
		_w666_,
		_w694_,
		_w6650_,
		_w6686_
	);
	LUT3 #(
		.INIT('h01)
	) name6653 (
		_w6685_,
		_w6686_,
		_w6684_,
		_w6687_
	);
	LUT4 #(
		.INIT('h95aa)
	) name6654 (
		\a[2] ,
		_w2598_,
		_w6335_,
		_w6687_,
		_w6688_
	);
	LUT4 #(
		.INIT('he100)
	) name6655 (
		_w6396_,
		_w6630_,
		_w6631_,
		_w6688_,
		_w6689_
	);
	LUT4 #(
		.INIT('h54ab)
	) name6656 (
		_w6404_,
		_w6626_,
		_w6627_,
		_w6629_,
		_w6690_
	);
	LUT2 #(
		.INIT('h9)
	) name6657 (
		_w6626_,
		_w6628_,
		_w6691_
	);
	LUT3 #(
		.INIT('h1e)
	) name6658 (
		_w6418_,
		_w6624_,
		_w6625_,
		_w6692_
	);
	LUT4 #(
		.INIT('h54ab)
	) name6659 (
		_w6424_,
		_w6620_,
		_w6621_,
		_w6623_,
		_w6693_
	);
	LUT3 #(
		.INIT('h70)
	) name6660 (
		_w1071_,
		_w1102_,
		_w6334_,
		_w6694_
	);
	LUT3 #(
		.INIT('h70)
	) name6661 (
		_w763_,
		_w983_,
		_w6657_,
		_w6695_
	);
	LUT3 #(
		.INIT('h70)
	) name6662 (
		_w1009_,
		_w1050_,
		_w6650_,
		_w6696_
	);
	LUT3 #(
		.INIT('h01)
	) name6663 (
		_w6695_,
		_w6696_,
		_w6694_,
		_w6697_
	);
	LUT4 #(
		.INIT('h6f00)
	) name6664 (
		_w2339_,
		_w2341_,
		_w6335_,
		_w6697_,
		_w6698_
	);
	LUT2 #(
		.INIT('h6)
	) name6665 (
		\a[2] ,
		_w6698_,
		_w6699_
	);
	LUT3 #(
		.INIT('h60)
	) name6666 (
		_w6620_,
		_w6622_,
		_w6699_,
		_w6700_
	);
	LUT3 #(
		.INIT('h1e)
	) name6667 (
		_w6438_,
		_w6618_,
		_w6619_,
		_w6701_
	);
	LUT4 #(
		.INIT('h54ab)
	) name6668 (
		_w6446_,
		_w6614_,
		_w6615_,
		_w6617_,
		_w6702_
	);
	LUT2 #(
		.INIT('h9)
	) name6669 (
		_w6614_,
		_w6616_,
		_w6703_
	);
	LUT3 #(
		.INIT('h1e)
	) name6670 (
		_w6460_,
		_w6612_,
		_w6613_,
		_w6704_
	);
	LUT4 #(
		.INIT('h54ab)
	) name6671 (
		_w6466_,
		_w6608_,
		_w6609_,
		_w6611_,
		_w6705_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6672 (
		_w1454_,
		_w1426_,
		_w1478_,
		_w6334_,
		_w6706_
	);
	LUT3 #(
		.INIT('h70)
	) name6673 (
		_w1325_,
		_w1367_,
		_w6657_,
		_w6707_
	);
	LUT3 #(
		.INIT('h70)
	) name6674 (
		_w1381_,
		_w1398_,
		_w6650_,
		_w6708_
	);
	LUT3 #(
		.INIT('h01)
	) name6675 (
		_w6707_,
		_w6708_,
		_w6706_,
		_w6709_
	);
	LUT4 #(
		.INIT('h6f00)
	) name6676 (
		_w2327_,
		_w2329_,
		_w6335_,
		_w6709_,
		_w6710_
	);
	LUT2 #(
		.INIT('h6)
	) name6677 (
		\a[2] ,
		_w6710_,
		_w6711_
	);
	LUT3 #(
		.INIT('h60)
	) name6678 (
		_w6608_,
		_w6610_,
		_w6711_,
		_w6712_
	);
	LUT3 #(
		.INIT('h1e)
	) name6679 (
		_w6480_,
		_w6606_,
		_w6607_,
		_w6713_
	);
	LUT4 #(
		.INIT('h54ab)
	) name6680 (
		_w6488_,
		_w6602_,
		_w6603_,
		_w6605_,
		_w6714_
	);
	LUT2 #(
		.INIT('h9)
	) name6681 (
		_w6602_,
		_w6604_,
		_w6715_
	);
	LUT3 #(
		.INIT('h1e)
	) name6682 (
		_w6502_,
		_w6600_,
		_w6601_,
		_w6716_
	);
	LUT4 #(
		.INIT('h54ab)
	) name6683 (
		_w6508_,
		_w6596_,
		_w6597_,
		_w6599_,
		_w6717_
	);
	LUT3 #(
		.INIT('h70)
	) name6684 (
		_w1692_,
		_w1723_,
		_w6657_,
		_w6718_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6685 (
		_w1751_,
		_w1742_,
		_w1771_,
		_w6650_,
		_w6719_
	);
	LUT3 #(
		.INIT('h70)
	) name6686 (
		_w1795_,
		_w1796_,
		_w6334_,
		_w6720_
	);
	LUT3 #(
		.INIT('h01)
	) name6687 (
		_w6719_,
		_w6720_,
		_w6718_,
		_w6721_
	);
	LUT4 #(
		.INIT('h6f00)
	) name6688 (
		_w2315_,
		_w2317_,
		_w6335_,
		_w6721_,
		_w6722_
	);
	LUT2 #(
		.INIT('h6)
	) name6689 (
		\a[2] ,
		_w6722_,
		_w6723_
	);
	LUT3 #(
		.INIT('h60)
	) name6690 (
		_w6596_,
		_w6598_,
		_w6723_,
		_w6724_
	);
	LUT3 #(
		.INIT('h1e)
	) name6691 (
		_w6523_,
		_w6593_,
		_w6595_,
		_w6725_
	);
	LUT4 #(
		.INIT('h54ab)
	) name6692 (
		_w6531_,
		_w6589_,
		_w6590_,
		_w6592_,
		_w6726_
	);
	LUT2 #(
		.INIT('h9)
	) name6693 (
		_w6589_,
		_w6591_,
		_w6727_
	);
	LUT3 #(
		.INIT('h1e)
	) name6694 (
		_w6545_,
		_w6586_,
		_w6588_,
		_w6728_
	);
	LUT4 #(
		.INIT('h54ab)
	) name6695 (
		_w6553_,
		_w6582_,
		_w6583_,
		_w6585_,
		_w6729_
	);
	LUT3 #(
		.INIT('h70)
	) name6696 (
		_w1973_,
		_w1997_,
		_w6650_,
		_w6730_
	);
	LUT3 #(
		.INIT('h70)
	) name6697 (
		_w1501_,
		_w1949_,
		_w6657_,
		_w6731_
	);
	LUT3 #(
		.INIT('h70)
	) name6698 (
		_w2023_,
		_w2055_,
		_w6334_,
		_w6732_
	);
	LUT3 #(
		.INIT('h01)
	) name6699 (
		_w6730_,
		_w6731_,
		_w6732_,
		_w6733_
	);
	LUT4 #(
		.INIT('h6f00)
	) name6700 (
		_w2303_,
		_w2305_,
		_w6335_,
		_w6733_,
		_w6734_
	);
	LUT4 #(
		.INIT('h1428)
	) name6701 (
		\a[2] ,
		_w6582_,
		_w6584_,
		_w6734_,
		_w6735_
	);
	LUT4 #(
		.INIT('h8241)
	) name6702 (
		\a[2] ,
		_w6582_,
		_w6584_,
		_w6734_,
		_w6736_
	);
	LUT2 #(
		.INIT('h9)
	) name6703 (
		_w6579_,
		_w6581_,
		_w6737_
	);
	LUT3 #(
		.INIT('h70)
	) name6704 (
		_w1973_,
		_w1997_,
		_w6657_,
		_w6738_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6705 (
		_w1874_,
		_w2076_,
		_w2099_,
		_w6334_,
		_w6739_
	);
	LUT3 #(
		.INIT('h70)
	) name6706 (
		_w2023_,
		_w2055_,
		_w6650_,
		_w6740_
	);
	LUT3 #(
		.INIT('h01)
	) name6707 (
		_w6739_,
		_w6738_,
		_w6740_,
		_w6741_
	);
	LUT4 #(
		.INIT('h6a55)
	) name6708 (
		\a[2] ,
		_w4151_,
		_w6335_,
		_w6741_,
		_w6742_
	);
	LUT2 #(
		.INIT('h1)
	) name6709 (
		_w6737_,
		_w6742_,
		_w6743_
	);
	LUT2 #(
		.INIT('h8)
	) name6710 (
		_w6737_,
		_w6742_,
		_w6744_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6711 (
		_w1874_,
		_w2076_,
		_w2099_,
		_w6650_,
		_w6745_
	);
	LUT3 #(
		.INIT('h70)
	) name6712 (
		_w2124_,
		_w2133_,
		_w6334_,
		_w6746_
	);
	LUT3 #(
		.INIT('h70)
	) name6713 (
		_w2023_,
		_w2055_,
		_w6657_,
		_w6747_
	);
	LUT3 #(
		.INIT('h01)
	) name6714 (
		_w6745_,
		_w6746_,
		_w6747_,
		_w6748_
	);
	LUT4 #(
		.INIT('h6f00)
	) name6715 (
		_w2299_,
		_w2301_,
		_w6335_,
		_w6748_,
		_w6749_
	);
	LUT3 #(
		.INIT('h69)
	) name6716 (
		_w6247_,
		_w6573_,
		_w6578_,
		_w6750_
	);
	LUT3 #(
		.INIT('h06)
	) name6717 (
		\a[2] ,
		_w6749_,
		_w6750_,
		_w6751_
	);
	LUT3 #(
		.INIT('h90)
	) name6718 (
		\a[2] ,
		_w6749_,
		_w6750_,
		_w6752_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6719 (
		_w1874_,
		_w2076_,
		_w2099_,
		_w6657_,
		_w6753_
	);
	LUT3 #(
		.INIT('h70)
	) name6720 (
		_w2124_,
		_w2133_,
		_w6650_,
		_w6754_
	);
	LUT3 #(
		.INIT('h70)
	) name6721 (
		_w2155_,
		_w2156_,
		_w6334_,
		_w6755_
	);
	LUT3 #(
		.INIT('h01)
	) name6722 (
		_w6754_,
		_w6755_,
		_w6753_,
		_w6756_
	);
	LUT4 #(
		.INIT('h95aa)
	) name6723 (
		\a[2] ,
		_w4209_,
		_w6335_,
		_w6756_,
		_w6757_
	);
	LUT3 #(
		.INIT('h8a)
	) name6724 (
		\a[5] ,
		_w6565_,
		_w6564_,
		_w6758_
	);
	LUT2 #(
		.INIT('h9)
	) name6725 (
		_w6572_,
		_w6758_,
		_w6759_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6726 (
		_w2193_,
		_w2183_,
		_w2213_,
		_w6334_,
		_w6760_
	);
	LUT3 #(
		.INIT('h70)
	) name6727 (
		_w2155_,
		_w2156_,
		_w6650_,
		_w6761_
	);
	LUT3 #(
		.INIT('h70)
	) name6728 (
		_w2124_,
		_w2133_,
		_w6657_,
		_w6762_
	);
	LUT3 #(
		.INIT('h01)
	) name6729 (
		_w6760_,
		_w6761_,
		_w6762_,
		_w6763_
	);
	LUT4 #(
		.INIT('h6f00)
	) name6730 (
		_w2295_,
		_w2297_,
		_w6335_,
		_w6763_,
		_w6764_
	);
	LUT4 #(
		.INIT('h0222)
	) name6731 (
		\a[5] ,
		_w34_,
		_w2228_,
		_w2262_,
		_w6765_
	);
	LUT2 #(
		.INIT('h9)
	) name6732 (
		_w6564_,
		_w6765_,
		_w6766_
	);
	LUT3 #(
		.INIT('h06)
	) name6733 (
		\a[2] ,
		_w6764_,
		_w6766_,
		_w6767_
	);
	LUT3 #(
		.INIT('h90)
	) name6734 (
		\a[2] ,
		_w6764_,
		_w6766_,
		_w6768_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6735 (
		_w2193_,
		_w2183_,
		_w2213_,
		_w6650_,
		_w6769_
	);
	LUT3 #(
		.INIT('h70)
	) name6736 (
		_w2155_,
		_w2156_,
		_w6657_,
		_w6770_
	);
	LUT3 #(
		.INIT('h70)
	) name6737 (
		_w2273_,
		_w2293_,
		_w6334_,
		_w6771_
	);
	LUT3 #(
		.INIT('h01)
	) name6738 (
		_w6769_,
		_w6770_,
		_w6771_,
		_w6772_
	);
	LUT3 #(
		.INIT('h70)
	) name6739 (
		_w4293_,
		_w6335_,
		_w6772_,
		_w6773_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name6740 (
		\a[0] ,
		_w2193_,
		_w2183_,
		_w2213_,
		_w6774_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name6741 (
		_w2263_,
		_w2294_,
		_w6332_,
		_w6774_,
		_w6775_
	);
	LUT4 #(
		.INIT('hac84)
	) name6742 (
		\a[2] ,
		_w6565_,
		_w6773_,
		_w6775_,
		_w6776_
	);
	LUT3 #(
		.INIT('h54)
	) name6743 (
		_w6767_,
		_w6768_,
		_w6776_,
		_w6777_
	);
	LUT4 #(
		.INIT('h0445)
	) name6744 (
		_w6752_,
		_w6757_,
		_w6759_,
		_w6777_,
		_w6778_
	);
	LUT4 #(
		.INIT('h4445)
	) name6745 (
		_w6743_,
		_w6744_,
		_w6751_,
		_w6778_,
		_w6779_
	);
	LUT3 #(
		.INIT('h54)
	) name6746 (
		_w6735_,
		_w6736_,
		_w6779_,
		_w6780_
	);
	LUT3 #(
		.INIT('h70)
	) name6747 (
		_w1973_,
		_w1997_,
		_w6334_,
		_w6781_
	);
	LUT3 #(
		.INIT('h70)
	) name6748 (
		_w1898_,
		_w1928_,
		_w6657_,
		_w6782_
	);
	LUT3 #(
		.INIT('h70)
	) name6749 (
		_w1501_,
		_w1949_,
		_w6650_,
		_w6783_
	);
	LUT3 #(
		.INIT('h01)
	) name6750 (
		_w6782_,
		_w6783_,
		_w6781_,
		_w6784_
	);
	LUT4 #(
		.INIT('h95aa)
	) name6751 (
		\a[2] ,
		_w4126_,
		_w6335_,
		_w6784_,
		_w6785_
	);
	LUT4 #(
		.INIT('h1501)
	) name6752 (
		_w6728_,
		_w6729_,
		_w6780_,
		_w6785_,
		_w6786_
	);
	LUT4 #(
		.INIT('h80a8)
	) name6753 (
		_w6728_,
		_w6729_,
		_w6780_,
		_w6785_,
		_w6787_
	);
	LUT3 #(
		.INIT('h70)
	) name6754 (
		_w1501_,
		_w1949_,
		_w6334_,
		_w6788_
	);
	LUT3 #(
		.INIT('h70)
	) name6755 (
		_w1898_,
		_w1928_,
		_w6650_,
		_w6789_
	);
	LUT3 #(
		.INIT('h70)
	) name6756 (
		_w1863_,
		_w1875_,
		_w6657_,
		_w6790_
	);
	LUT3 #(
		.INIT('h01)
	) name6757 (
		_w6789_,
		_w6790_,
		_w6788_,
		_w6791_
	);
	LUT4 #(
		.INIT('h6f00)
	) name6758 (
		_w2307_,
		_w2309_,
		_w6335_,
		_w6791_,
		_w6792_
	);
	LUT2 #(
		.INIT('h6)
	) name6759 (
		\a[2] ,
		_w6792_,
		_w6793_
	);
	LUT3 #(
		.INIT('h45)
	) name6760 (
		_w6786_,
		_w6787_,
		_w6793_,
		_w6794_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6761 (
		_w1817_,
		_w1799_,
		_w1840_,
		_w6657_,
		_w6795_
	);
	LUT3 #(
		.INIT('h70)
	) name6762 (
		_w1898_,
		_w1928_,
		_w6334_,
		_w6796_
	);
	LUT3 #(
		.INIT('h70)
	) name6763 (
		_w1863_,
		_w1875_,
		_w6650_,
		_w6797_
	);
	LUT3 #(
		.INIT('h01)
	) name6764 (
		_w6796_,
		_w6797_,
		_w6795_,
		_w6798_
	);
	LUT4 #(
		.INIT('h6a55)
	) name6765 (
		\a[2] ,
		_w3972_,
		_w6335_,
		_w6798_,
		_w6799_
	);
	LUT4 #(
		.INIT('ha880)
	) name6766 (
		_w6726_,
		_w6727_,
		_w6794_,
		_w6799_,
		_w6800_
	);
	LUT4 #(
		.INIT('h0115)
	) name6767 (
		_w6726_,
		_w6727_,
		_w6794_,
		_w6799_,
		_w6801_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6768 (
		_w1817_,
		_w1799_,
		_w1840_,
		_w6650_,
		_w6802_
	);
	LUT3 #(
		.INIT('h70)
	) name6769 (
		_w1795_,
		_w1796_,
		_w6657_,
		_w6803_
	);
	LUT3 #(
		.INIT('h70)
	) name6770 (
		_w1863_,
		_w1875_,
		_w6334_,
		_w6804_
	);
	LUT3 #(
		.INIT('h01)
	) name6771 (
		_w6803_,
		_w6804_,
		_w6802_,
		_w6805_
	);
	LUT4 #(
		.INIT('h6f00)
	) name6772 (
		_w2311_,
		_w2313_,
		_w6335_,
		_w6805_,
		_w6806_
	);
	LUT2 #(
		.INIT('h9)
	) name6773 (
		\a[2] ,
		_w6806_,
		_w6807_
	);
	LUT3 #(
		.INIT('h45)
	) name6774 (
		_w6800_,
		_w6801_,
		_w6807_,
		_w6808_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6775 (
		_w1751_,
		_w1742_,
		_w1771_,
		_w6657_,
		_w6809_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6776 (
		_w1817_,
		_w1799_,
		_w1840_,
		_w6334_,
		_w6810_
	);
	LUT3 #(
		.INIT('h70)
	) name6777 (
		_w1795_,
		_w1796_,
		_w6650_,
		_w6811_
	);
	LUT3 #(
		.INIT('h01)
	) name6778 (
		_w6810_,
		_w6811_,
		_w6809_,
		_w6812_
	);
	LUT4 #(
		.INIT('h6a55)
	) name6779 (
		\a[2] ,
		_w3909_,
		_w6335_,
		_w6812_,
		_w6813_
	);
	LUT3 #(
		.INIT('h09)
	) name6780 (
		_w6596_,
		_w6598_,
		_w6723_,
		_w6814_
	);
	LUT4 #(
		.INIT('h040d)
	) name6781 (
		_w6725_,
		_w6808_,
		_w6814_,
		_w6813_,
		_w6815_
	);
	LUT3 #(
		.INIT('h70)
	) name6782 (
		_w1692_,
		_w1723_,
		_w6650_,
		_w6816_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6783 (
		_w1751_,
		_w1742_,
		_w1771_,
		_w6334_,
		_w6817_
	);
	LUT3 #(
		.INIT('h70)
	) name6784 (
		_w1620_,
		_w1661_,
		_w6657_,
		_w6818_
	);
	LUT3 #(
		.INIT('h01)
	) name6785 (
		_w6817_,
		_w6818_,
		_w6816_,
		_w6819_
	);
	LUT4 #(
		.INIT('h95aa)
	) name6786 (
		\a[2] ,
		_w3599_,
		_w6335_,
		_w6819_,
		_w6820_
	);
	LUT4 #(
		.INIT('h02ab)
	) name6787 (
		_w6717_,
		_w6724_,
		_w6815_,
		_w6820_,
		_w6821_
	);
	LUT3 #(
		.INIT('h70)
	) name6788 (
		_w1692_,
		_w1723_,
		_w6334_,
		_w6822_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6789 (
		_w1584_,
		_w1569_,
		_w1606_,
		_w6657_,
		_w6823_
	);
	LUT3 #(
		.INIT('h70)
	) name6790 (
		_w1620_,
		_w1661_,
		_w6650_,
		_w6824_
	);
	LUT3 #(
		.INIT('h01)
	) name6791 (
		_w6823_,
		_w6824_,
		_w6822_,
		_w6825_
	);
	LUT4 #(
		.INIT('h6f00)
	) name6792 (
		_w2319_,
		_w2321_,
		_w6335_,
		_w6825_,
		_w6826_
	);
	LUT2 #(
		.INIT('h6)
	) name6793 (
		\a[2] ,
		_w6826_,
		_w6827_
	);
	LUT3 #(
		.INIT('h8e)
	) name6794 (
		_w6716_,
		_w6821_,
		_w6827_,
		_w6828_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6795 (
		_w1584_,
		_w1569_,
		_w1606_,
		_w6650_,
		_w6829_
	);
	LUT3 #(
		.INIT('h70)
	) name6796 (
		_w1501_,
		_w1545_,
		_w6657_,
		_w6830_
	);
	LUT3 #(
		.INIT('h70)
	) name6797 (
		_w1620_,
		_w1661_,
		_w6334_,
		_w6831_
	);
	LUT3 #(
		.INIT('h01)
	) name6798 (
		_w6829_,
		_w6830_,
		_w6831_,
		_w6832_
	);
	LUT4 #(
		.INIT('h6a55)
	) name6799 (
		\a[2] ,
		_w3495_,
		_w6335_,
		_w6832_,
		_w6833_
	);
	LUT4 #(
		.INIT('ha880)
	) name6800 (
		_w6714_,
		_w6715_,
		_w6828_,
		_w6833_,
		_w6834_
	);
	LUT4 #(
		.INIT('h0115)
	) name6801 (
		_w6714_,
		_w6715_,
		_w6828_,
		_w6833_,
		_w6835_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6802 (
		_w1454_,
		_w1426_,
		_w1478_,
		_w6657_,
		_w6836_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6803 (
		_w1584_,
		_w1569_,
		_w1606_,
		_w6334_,
		_w6837_
	);
	LUT3 #(
		.INIT('h70)
	) name6804 (
		_w1501_,
		_w1545_,
		_w6650_,
		_w6838_
	);
	LUT3 #(
		.INIT('h01)
	) name6805 (
		_w6837_,
		_w6838_,
		_w6836_,
		_w6839_
	);
	LUT4 #(
		.INIT('h6f00)
	) name6806 (
		_w2323_,
		_w2325_,
		_w6335_,
		_w6839_,
		_w6840_
	);
	LUT2 #(
		.INIT('h9)
	) name6807 (
		\a[2] ,
		_w6840_,
		_w6841_
	);
	LUT3 #(
		.INIT('h45)
	) name6808 (
		_w6834_,
		_w6835_,
		_w6841_,
		_w6842_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6809 (
		_w1454_,
		_w1426_,
		_w1478_,
		_w6650_,
		_w6843_
	);
	LUT3 #(
		.INIT('h70)
	) name6810 (
		_w1381_,
		_w1398_,
		_w6657_,
		_w6844_
	);
	LUT3 #(
		.INIT('h70)
	) name6811 (
		_w1501_,
		_w1545_,
		_w6334_,
		_w6845_
	);
	LUT3 #(
		.INIT('h01)
	) name6812 (
		_w6844_,
		_w6845_,
		_w6843_,
		_w6846_
	);
	LUT4 #(
		.INIT('h6a55)
	) name6813 (
		\a[2] ,
		_w3362_,
		_w6335_,
		_w6846_,
		_w6847_
	);
	LUT3 #(
		.INIT('h09)
	) name6814 (
		_w6608_,
		_w6610_,
		_w6711_,
		_w6848_
	);
	LUT4 #(
		.INIT('h040d)
	) name6815 (
		_w6713_,
		_w6842_,
		_w6848_,
		_w6847_,
		_w6849_
	);
	LUT3 #(
		.INIT('h70)
	) name6816 (
		_w1381_,
		_w1398_,
		_w6334_,
		_w6850_
	);
	LUT3 #(
		.INIT('h70)
	) name6817 (
		_w1325_,
		_w1367_,
		_w6650_,
		_w6851_
	);
	LUT3 #(
		.INIT('h70)
	) name6818 (
		_w1253_,
		_w1294_,
		_w6657_,
		_w6852_
	);
	LUT3 #(
		.INIT('h01)
	) name6819 (
		_w6851_,
		_w6852_,
		_w6850_,
		_w6853_
	);
	LUT4 #(
		.INIT('h95aa)
	) name6820 (
		\a[2] ,
		_w3182_,
		_w6335_,
		_w6853_,
		_w6854_
	);
	LUT4 #(
		.INIT('h02ab)
	) name6821 (
		_w6705_,
		_w6712_,
		_w6849_,
		_w6854_,
		_w6855_
	);
	LUT3 #(
		.INIT('h70)
	) name6822 (
		_w1202_,
		_w1233_,
		_w6657_,
		_w6856_
	);
	LUT3 #(
		.INIT('h70)
	) name6823 (
		_w1325_,
		_w1367_,
		_w6334_,
		_w6857_
	);
	LUT3 #(
		.INIT('h70)
	) name6824 (
		_w1253_,
		_w1294_,
		_w6650_,
		_w6858_
	);
	LUT3 #(
		.INIT('h01)
	) name6825 (
		_w6857_,
		_w6858_,
		_w6856_,
		_w6859_
	);
	LUT4 #(
		.INIT('h6f00)
	) name6826 (
		_w2331_,
		_w2333_,
		_w6335_,
		_w6859_,
		_w6860_
	);
	LUT2 #(
		.INIT('h6)
	) name6827 (
		\a[2] ,
		_w6860_,
		_w6861_
	);
	LUT3 #(
		.INIT('h8e)
	) name6828 (
		_w6704_,
		_w6855_,
		_w6861_,
		_w6862_
	);
	LUT3 #(
		.INIT('h70)
	) name6829 (
		_w1202_,
		_w1233_,
		_w6650_,
		_w6863_
	);
	LUT3 #(
		.INIT('h70)
	) name6830 (
		_w1253_,
		_w1294_,
		_w6334_,
		_w6864_
	);
	LUT3 #(
		.INIT('h70)
	) name6831 (
		_w1136_,
		_w1187_,
		_w6657_,
		_w6865_
	);
	LUT3 #(
		.INIT('h01)
	) name6832 (
		_w6864_,
		_w6865_,
		_w6863_,
		_w6866_
	);
	LUT4 #(
		.INIT('h6a55)
	) name6833 (
		\a[2] ,
		_w3067_,
		_w6335_,
		_w6866_,
		_w6867_
	);
	LUT4 #(
		.INIT('ha880)
	) name6834 (
		_w6702_,
		_w6703_,
		_w6862_,
		_w6867_,
		_w6868_
	);
	LUT4 #(
		.INIT('h0115)
	) name6835 (
		_w6702_,
		_w6703_,
		_w6862_,
		_w6867_,
		_w6869_
	);
	LUT3 #(
		.INIT('h70)
	) name6836 (
		_w1136_,
		_w1187_,
		_w6650_,
		_w6870_
	);
	LUT3 #(
		.INIT('h70)
	) name6837 (
		_w1071_,
		_w1102_,
		_w6657_,
		_w6871_
	);
	LUT3 #(
		.INIT('h70)
	) name6838 (
		_w1202_,
		_w1233_,
		_w6334_,
		_w6872_
	);
	LUT3 #(
		.INIT('h01)
	) name6839 (
		_w6871_,
		_w6872_,
		_w6870_,
		_w6873_
	);
	LUT4 #(
		.INIT('h6f00)
	) name6840 (
		_w2335_,
		_w2337_,
		_w6335_,
		_w6873_,
		_w6874_
	);
	LUT2 #(
		.INIT('h9)
	) name6841 (
		\a[2] ,
		_w6874_,
		_w6875_
	);
	LUT3 #(
		.INIT('h45)
	) name6842 (
		_w6868_,
		_w6869_,
		_w6875_,
		_w6876_
	);
	LUT3 #(
		.INIT('h70)
	) name6843 (
		_w1136_,
		_w1187_,
		_w6334_,
		_w6877_
	);
	LUT3 #(
		.INIT('h70)
	) name6844 (
		_w1009_,
		_w1050_,
		_w6657_,
		_w6878_
	);
	LUT3 #(
		.INIT('h70)
	) name6845 (
		_w1071_,
		_w1102_,
		_w6650_,
		_w6879_
	);
	LUT3 #(
		.INIT('h01)
	) name6846 (
		_w6878_,
		_w6879_,
		_w6877_,
		_w6880_
	);
	LUT4 #(
		.INIT('h6a55)
	) name6847 (
		\a[2] ,
		_w2936_,
		_w6335_,
		_w6880_,
		_w6881_
	);
	LUT3 #(
		.INIT('h09)
	) name6848 (
		_w6620_,
		_w6622_,
		_w6699_,
		_w6882_
	);
	LUT4 #(
		.INIT('h040d)
	) name6849 (
		_w6701_,
		_w6876_,
		_w6882_,
		_w6881_,
		_w6883_
	);
	LUT3 #(
		.INIT('h70)
	) name6850 (
		_w1009_,
		_w1050_,
		_w6334_,
		_w6884_
	);
	LUT3 #(
		.INIT('h70)
	) name6851 (
		_w871_,
		_w927_,
		_w6657_,
		_w6885_
	);
	LUT3 #(
		.INIT('h70)
	) name6852 (
		_w763_,
		_w983_,
		_w6650_,
		_w6886_
	);
	LUT3 #(
		.INIT('h01)
	) name6853 (
		_w6885_,
		_w6886_,
		_w6884_,
		_w6887_
	);
	LUT4 #(
		.INIT('h95aa)
	) name6854 (
		\a[2] ,
		_w2839_,
		_w6335_,
		_w6887_,
		_w6888_
	);
	LUT4 #(
		.INIT('h02ab)
	) name6855 (
		_w6693_,
		_w6700_,
		_w6883_,
		_w6888_,
		_w6889_
	);
	LUT3 #(
		.INIT('h70)
	) name6856 (
		_w763_,
		_w983_,
		_w6334_,
		_w6890_
	);
	LUT3 #(
		.INIT('h70)
	) name6857 (
		_w871_,
		_w927_,
		_w6650_,
		_w6891_
	);
	LUT3 #(
		.INIT('h70)
	) name6858 (
		_w801_,
		_w851_,
		_w6657_,
		_w6892_
	);
	LUT3 #(
		.INIT('h01)
	) name6859 (
		_w6891_,
		_w6892_,
		_w6890_,
		_w6893_
	);
	LUT4 #(
		.INIT('h6f00)
	) name6860 (
		_w2343_,
		_w2345_,
		_w6335_,
		_w6893_,
		_w6894_
	);
	LUT2 #(
		.INIT('h6)
	) name6861 (
		\a[2] ,
		_w6894_,
		_w6895_
	);
	LUT4 #(
		.INIT('h80a8)
	) name6862 (
		_w6691_,
		_w6692_,
		_w6889_,
		_w6895_,
		_w6896_
	);
	LUT4 #(
		.INIT('h1501)
	) name6863 (
		_w6691_,
		_w6692_,
		_w6889_,
		_w6895_,
		_w6897_
	);
	LUT3 #(
		.INIT('h70)
	) name6864 (
		_w725_,
		_w764_,
		_w6657_,
		_w6898_
	);
	LUT3 #(
		.INIT('h70)
	) name6865 (
		_w801_,
		_w851_,
		_w6650_,
		_w6899_
	);
	LUT3 #(
		.INIT('h70)
	) name6866 (
		_w871_,
		_w927_,
		_w6334_,
		_w6900_
	);
	LUT3 #(
		.INIT('h01)
	) name6867 (
		_w6899_,
		_w6900_,
		_w6898_,
		_w6901_
	);
	LUT4 #(
		.INIT('h6a55)
	) name6868 (
		\a[2] ,
		_w2724_,
		_w6335_,
		_w6901_,
		_w6902_
	);
	LUT3 #(
		.INIT('h45)
	) name6869 (
		_w6896_,
		_w6897_,
		_w6902_,
		_w6903_
	);
	LUT3 #(
		.INIT('h70)
	) name6870 (
		_w725_,
		_w764_,
		_w6650_,
		_w6904_
	);
	LUT3 #(
		.INIT('h70)
	) name6871 (
		_w801_,
		_w851_,
		_w6334_,
		_w6905_
	);
	LUT3 #(
		.INIT('h70)
	) name6872 (
		_w666_,
		_w694_,
		_w6657_,
		_w6906_
	);
	LUT3 #(
		.INIT('h01)
	) name6873 (
		_w6905_,
		_w6906_,
		_w6904_,
		_w6907_
	);
	LUT4 #(
		.INIT('h6f00)
	) name6874 (
		_w2347_,
		_w2349_,
		_w6335_,
		_w6907_,
		_w6908_
	);
	LUT2 #(
		.INIT('h9)
	) name6875 (
		\a[2] ,
		_w6908_,
		_w6909_
	);
	LUT4 #(
		.INIT('h001e)
	) name6876 (
		_w6396_,
		_w6630_,
		_w6631_,
		_w6688_,
		_w6910_
	);
	LUT4 #(
		.INIT('h040d)
	) name6877 (
		_w6690_,
		_w6903_,
		_w6910_,
		_w6909_,
		_w6911_
	);
	LUT3 #(
		.INIT('h60)
	) name6878 (
		_w6632_,
		_w6634_,
		_w6682_,
		_w6912_
	);
	LUT3 #(
		.INIT('h96)
	) name6879 (
		_w6632_,
		_w6634_,
		_w6682_,
		_w6913_
	);
	LUT4 #(
		.INIT('h5554)
	) name6880 (
		_w6683_,
		_w6689_,
		_w6911_,
		_w6912_,
		_w6914_
	);
	LUT2 #(
		.INIT('h4)
	) name6881 (
		_w6670_,
		_w6675_,
		_w6915_
	);
	LUT2 #(
		.INIT('h9)
	) name6882 (
		_w6670_,
		_w6675_,
		_w6916_
	);
	LUT3 #(
		.INIT('h54)
	) name6883 (
		_w6676_,
		_w6914_,
		_w6915_,
		_w6917_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name6884 (
		_w6376_,
		_w6636_,
		_w6637_,
		_w6668_,
		_w6918_
	);
	LUT4 #(
		.INIT('h2b00)
	) name6885 (
		_w6670_,
		_w6675_,
		_w6914_,
		_w6918_,
		_w6919_
	);
	LUT3 #(
		.INIT('h60)
	) name6886 (
		_w6638_,
		_w6640_,
		_w6660_,
		_w6920_
	);
	LUT3 #(
		.INIT('h96)
	) name6887 (
		_w6638_,
		_w6640_,
		_w6660_,
		_w6921_
	);
	LUT4 #(
		.INIT('h5501)
	) name6888 (
		_w6661_,
		_w6669_,
		_w6919_,
		_w6920_,
		_w6922_
	);
	LUT2 #(
		.INIT('h4)
	) name6889 (
		_w6647_,
		_w6653_,
		_w6923_
	);
	LUT2 #(
		.INIT('h9)
	) name6890 (
		_w6647_,
		_w6653_,
		_w6924_
	);
	LUT3 #(
		.INIT('h54)
	) name6891 (
		_w6654_,
		_w6922_,
		_w6923_,
		_w6925_
	);
	LUT4 #(
		.INIT('h088a)
	) name6892 (
		_w6646_,
		_w6647_,
		_w6653_,
		_w6922_,
		_w6926_
	);
	LUT2 #(
		.INIT('h4)
	) name6893 (
		_w6331_,
		_w6346_,
		_w6927_
	);
	LUT2 #(
		.INIT('h9)
	) name6894 (
		_w6331_,
		_w6346_,
		_w6928_
	);
	LUT4 #(
		.INIT('h5501)
	) name6895 (
		_w6347_,
		_w6645_,
		_w6926_,
		_w6927_,
		_w6929_
	);
	LUT4 #(
		.INIT('h00b2)
	) name6896 (
		_w6320_,
		_w6321_,
		_w6327_,
		_w6329_,
		_w6930_
	);
	LUT4 #(
		.INIT('hb24d)
	) name6897 (
		_w6320_,
		_w6321_,
		_w6327_,
		_w6329_,
		_w6931_
	);
	LUT3 #(
		.INIT('h54)
	) name6898 (
		_w6330_,
		_w6929_,
		_w6930_,
		_w6932_
	);
	LUT4 #(
		.INIT('h20a2)
	) name6899 (
		_w6044_,
		_w6328_,
		_w6329_,
		_w6929_,
		_w6933_
	);
	LUT4 #(
		.INIT('h6566)
	) name6900 (
		_w5522_,
		_w5766_,
		_w5767_,
		_w5769_,
		_w6934_
	);
	LUT4 #(
		.INIT('h0155)
	) name6901 (
		_w5770_,
		_w6043_,
		_w6933_,
		_w6934_,
		_w6935_
	);
	LUT2 #(
		.INIT('h2)
	) name6902 (
		_w5519_,
		_w5520_,
		_w6936_
	);
	LUT2 #(
		.INIT('h9)
	) name6903 (
		_w5519_,
		_w5520_,
		_w6937_
	);
	LUT3 #(
		.INIT('h54)
	) name6904 (
		_w5521_,
		_w6935_,
		_w6936_,
		_w6938_
	);
	LUT4 #(
		.INIT('h20a2)
	) name6905 (
		_w5283_,
		_w5519_,
		_w5520_,
		_w6935_,
		_w6939_
	);
	LUT4 #(
		.INIT('h4445)
	) name6906 (
		_w5065_,
		_w5066_,
		_w5282_,
		_w6939_,
		_w6940_
	);
	LUT3 #(
		.INIT('h90)
	) name6907 (
		_w4690_,
		_w4692_,
		_w4871_,
		_w6941_
	);
	LUT3 #(
		.INIT('h69)
	) name6908 (
		_w4690_,
		_w4692_,
		_w4871_,
		_w6942_
	);
	LUT3 #(
		.INIT('h54)
	) name6909 (
		_w4872_,
		_w6940_,
		_w6941_,
		_w6943_
	);
	LUT4 #(
		.INIT('h088a)
	) name6910 (
		_w4696_,
		_w4697_,
		_w4871_,
		_w6940_,
		_w6944_
	);
	LUT2 #(
		.INIT('h4)
	) name6911 (
		_w4456_,
		_w4531_,
		_w6945_
	);
	LUT2 #(
		.INIT('h9)
	) name6912 (
		_w4456_,
		_w4531_,
		_w6946_
	);
	LUT4 #(
		.INIT('h5501)
	) name6913 (
		_w4532_,
		_w4695_,
		_w6944_,
		_w6945_,
		_w6947_
	);
	LUT3 #(
		.INIT('h60)
	) name6914 (
		_w4373_,
		_w4375_,
		_w4453_,
		_w6948_
	);
	LUT3 #(
		.INIT('h96)
	) name6915 (
		_w4373_,
		_w4375_,
		_w4453_,
		_w6949_
	);
	LUT3 #(
		.INIT('h54)
	) name6916 (
		_w4455_,
		_w6947_,
		_w6948_,
		_w6950_
	);
	LUT4 #(
		.INIT('h20a2)
	) name6917 (
		_w4379_,
		_w4453_,
		_w4454_,
		_w6947_,
		_w6951_
	);
	LUT4 #(
		.INIT('h4445)
	) name6918 (
		_w4097_,
		_w4098_,
		_w4378_,
		_w6951_,
		_w6952_
	);
	LUT3 #(
		.INIT('h54)
	) name6919 (
		_w4028_,
		_w4029_,
		_w6952_,
		_w6953_
	);
	LUT4 #(
		.INIT('h022a)
	) name6920 (
		_w3883_,
		_w4025_,
		_w4027_,
		_w6952_,
		_w6954_
	);
	LUT2 #(
		.INIT('h4)
	) name6921 (
		_w3707_,
		_w3770_,
		_w6955_
	);
	LUT2 #(
		.INIT('h9)
	) name6922 (
		_w3707_,
		_w3770_,
		_w6956_
	);
	LUT4 #(
		.INIT('h5501)
	) name6923 (
		_w3771_,
		_w3882_,
		_w6954_,
		_w6955_,
		_w6957_
	);
	LUT3 #(
		.INIT('h54)
	) name6924 (
		_w3704_,
		_w3705_,
		_w6957_,
		_w6958_
	);
	LUT4 #(
		.INIT('h20a2)
	) name6925 (
		_w3651_,
		_w3701_,
		_w3703_,
		_w6957_,
		_w6959_
	);
	LUT4 #(
		.INIT('h4445)
	) name6926 (
		_w3407_,
		_w3408_,
		_w3650_,
		_w6959_,
		_w6960_
	);
	LUT3 #(
		.INIT('h60)
	) name6927 (
		_w3252_,
		_w3254_,
		_w3307_,
		_w6961_
	);
	LUT3 #(
		.INIT('h96)
	) name6928 (
		_w3252_,
		_w3254_,
		_w3307_,
		_w6962_
	);
	LUT3 #(
		.INIT('h54)
	) name6929 (
		_w3308_,
		_w6960_,
		_w6961_,
		_w6963_
	);
	LUT4 #(
		.INIT('h088a)
	) name6930 (
		_w3258_,
		_w3259_,
		_w3307_,
		_w6960_,
		_w6964_
	);
	LUT2 #(
		.INIT('h1)
	) name6931 (
		_w3008_,
		_w3218_,
		_w6965_
	);
	LUT2 #(
		.INIT('h6)
	) name6932 (
		_w3008_,
		_w3218_,
		_w6966_
	);
	LUT4 #(
		.INIT('h5501)
	) name6933 (
		_w3219_,
		_w3257_,
		_w6964_,
		_w6965_,
		_w6967_
	);
	LUT3 #(
		.INIT('h60)
	) name6934 (
		_w2978_,
		_w2980_,
		_w3005_,
		_w6968_
	);
	LUT3 #(
		.INIT('h96)
	) name6935 (
		_w2978_,
		_w2980_,
		_w3005_,
		_w6969_
	);
	LUT3 #(
		.INIT('h54)
	) name6936 (
		_w3007_,
		_w6967_,
		_w6968_,
		_w6970_
	);
	LUT4 #(
		.INIT('h54ab)
	) name6937 (
		_w2972_,
		_w2978_,
		_w2979_,
		_w2982_,
		_w6971_
	);
	LUT4 #(
		.INIT('h4d00)
	) name6938 (
		_w3005_,
		_w3006_,
		_w6967_,
		_w6971_,
		_w6972_
	);
	LUT2 #(
		.INIT('h2)
	) name6939 (
		_w2884_,
		_w2885_,
		_w6973_
	);
	LUT2 #(
		.INIT('h9)
	) name6940 (
		_w2884_,
		_w2885_,
		_w6974_
	);
	LUT4 #(
		.INIT('h5501)
	) name6941 (
		_w2886_,
		_w2983_,
		_w6972_,
		_w6973_,
		_w6975_
	);
	LUT3 #(
		.INIT('h54)
	) name6942 (
		_w2870_,
		_w2871_,
		_w6975_,
		_w6976_
	);
	LUT3 #(
		.INIT('he1)
	) name6943 (
		_w2613_,
		_w2620_,
		_w2621_,
		_w6977_
	);
	LUT4 #(
		.INIT('h4d00)
	) name6944 (
		_w2867_,
		_w2869_,
		_w6975_,
		_w6977_,
		_w6978_
	);
	LUT2 #(
		.INIT('h1)
	) name6945 (
		_w2547_,
		_w2558_,
		_w6979_
	);
	LUT2 #(
		.INIT('h6)
	) name6946 (
		_w2547_,
		_w2558_,
		_w6980_
	);
	LUT4 #(
		.INIT('h5501)
	) name6947 (
		_w2559_,
		_w2622_,
		_w6978_,
		_w6979_,
		_w6981_
	);
	LUT3 #(
		.INIT('h54)
	) name6948 (
		_w2544_,
		_w2545_,
		_w6981_,
		_w6982_
	);
	LUT4 #(
		.INIT('h20a2)
	) name6949 (
		_w2412_,
		_w2541_,
		_w2543_,
		_w6981_,
		_w6983_
	);
	LUT4 #(
		.INIT('h5557)
	) name6950 (
		_w122_,
		_w55_,
		_w52_,
		_w59_,
		_w6984_
	);
	LUT4 #(
		.INIT('h8000)
	) name6951 (
		_w302_,
		_w305_,
		_w1648_,
		_w6984_,
		_w6985_
	);
	LUT2 #(
		.INIT('h8)
	) name6952 (
		_w327_,
		_w6985_,
		_w6986_
	);
	LUT2 #(
		.INIT('h8)
	) name6953 (
		_w416_,
		_w6986_,
		_w6987_
	);
	LUT3 #(
		.INIT('h80)
	) name6954 (
		_w486_,
		_w487_,
		_w6987_,
		_w6988_
	);
	LUT2 #(
		.INIT('h8)
	) name6955 (
		_w330_,
		_w6988_,
		_w6989_
	);
	LUT2 #(
		.INIT('h6)
	) name6956 (
		_w330_,
		_w6988_,
		_w6990_
	);
	LUT4 #(
		.INIT('h00d4)
	) name6957 (
		_w157_,
		_w330_,
		_w2362_,
		_w6990_,
		_w6991_
	);
	LUT4 #(
		.INIT('h2b00)
	) name6958 (
		_w157_,
		_w330_,
		_w2362_,
		_w6990_,
		_w6992_
	);
	LUT4 #(
		.INIT('hba45)
	) name6959 (
		_w331_,
		_w332_,
		_w2362_,
		_w6990_,
		_w6993_
	);
	LUT3 #(
		.INIT('h1e)
	) name6960 (
		_w2411_,
		_w6983_,
		_w6993_,
		_w6994_
	);
	LUT4 #(
		.INIT('h4504)
	) name6961 (
		_w2412_,
		_w2541_,
		_w2543_,
		_w6981_,
		_w6995_
	);
	LUT4 #(
		.INIT('h6665)
	) name6962 (
		_w2412_,
		_w2544_,
		_w2545_,
		_w6981_,
		_w6996_
	);
	LUT4 #(
		.INIT('h4182)
	) name6963 (
		_w2411_,
		_w2412_,
		_w6982_,
		_w6993_,
		_w6997_
	);
	LUT4 #(
		.INIT('h8218)
	) name6964 (
		_w2412_,
		_w2541_,
		_w2543_,
		_w6981_,
		_w6998_
	);
	LUT3 #(
		.INIT('h1e)
	) name6965 (
		_w2622_,
		_w6978_,
		_w6980_,
		_w6999_
	);
	LUT3 #(
		.INIT('h90)
	) name6966 (
		_w2546_,
		_w6981_,
		_w6999_,
		_w7000_
	);
	LUT4 #(
		.INIT('h00b2)
	) name6967 (
		_w2867_,
		_w2869_,
		_w6975_,
		_w6977_,
		_w7001_
	);
	LUT4 #(
		.INIT('h54ab)
	) name6968 (
		_w2870_,
		_w2871_,
		_w6975_,
		_w6977_,
		_w7002_
	);
	LUT4 #(
		.INIT('h4182)
	) name6969 (
		_w2622_,
		_w6976_,
		_w6977_,
		_w6980_,
		_w7003_
	);
	LUT4 #(
		.INIT('h9204)
	) name6970 (
		_w2867_,
		_w2869_,
		_w6975_,
		_w6977_,
		_w7004_
	);
	LUT3 #(
		.INIT('h1e)
	) name6971 (
		_w2983_,
		_w6972_,
		_w6974_,
		_w7005_
	);
	LUT3 #(
		.INIT('h90)
	) name6972 (
		_w2872_,
		_w6975_,
		_w7005_,
		_w7006_
	);
	LUT4 #(
		.INIT('h00b2)
	) name6973 (
		_w3005_,
		_w3006_,
		_w6967_,
		_w6971_,
		_w7007_
	);
	LUT4 #(
		.INIT('h54ab)
	) name6974 (
		_w3007_,
		_w6967_,
		_w6968_,
		_w6971_,
		_w7008_
	);
	LUT4 #(
		.INIT('h9204)
	) name6975 (
		_w2981_,
		_w2982_,
		_w6970_,
		_w6974_,
		_w7009_
	);
	LUT4 #(
		.INIT('h9204)
	) name6976 (
		_w3005_,
		_w3006_,
		_w6967_,
		_w6971_,
		_w7010_
	);
	LUT3 #(
		.INIT('h1e)
	) name6977 (
		_w3257_,
		_w6964_,
		_w6966_,
		_w7011_
	);
	LUT3 #(
		.INIT('h90)
	) name6978 (
		_w6967_,
		_w6969_,
		_w7011_,
		_w7012_
	);
	LUT4 #(
		.INIT('h5110)
	) name6979 (
		_w3258_,
		_w3259_,
		_w3307_,
		_w6960_,
		_w7013_
	);
	LUT4 #(
		.INIT('h6665)
	) name6980 (
		_w3258_,
		_w3308_,
		_w6960_,
		_w6961_,
		_w7014_
	);
	LUT4 #(
		.INIT('h9204)
	) name6981 (
		_w3255_,
		_w3256_,
		_w6963_,
		_w6966_,
		_w7015_
	);
	LUT4 #(
		.INIT('h8224)
	) name6982 (
		_w3258_,
		_w3259_,
		_w3307_,
		_w6960_,
		_w7016_
	);
	LUT3 #(
		.INIT('h56)
	) name6983 (
		_w3409_,
		_w3650_,
		_w6959_,
		_w7017_
	);
	LUT3 #(
		.INIT('h90)
	) name6984 (
		_w6960_,
		_w6962_,
		_w7017_,
		_w7018_
	);
	LUT4 #(
		.INIT('h4504)
	) name6985 (
		_w3651_,
		_w3701_,
		_w3703_,
		_w6957_,
		_w7019_
	);
	LUT4 #(
		.INIT('h6665)
	) name6986 (
		_w3651_,
		_w3704_,
		_w3705_,
		_w6957_,
		_w7020_
	);
	LUT4 #(
		.INIT('h8224)
	) name6987 (
		_w3409_,
		_w3410_,
		_w3649_,
		_w6958_,
		_w7021_
	);
	LUT4 #(
		.INIT('h8218)
	) name6988 (
		_w3651_,
		_w3701_,
		_w3703_,
		_w6957_,
		_w7022_
	);
	LUT3 #(
		.INIT('h1e)
	) name6989 (
		_w3882_,
		_w6954_,
		_w6956_,
		_w7023_
	);
	LUT3 #(
		.INIT('h90)
	) name6990 (
		_w3706_,
		_w6957_,
		_w7023_,
		_w7024_
	);
	LUT4 #(
		.INIT('h5440)
	) name6991 (
		_w3883_,
		_w4025_,
		_w4027_,
		_w6952_,
		_w7025_
	);
	LUT4 #(
		.INIT('h6665)
	) name6992 (
		_w3883_,
		_w4028_,
		_w4029_,
		_w6952_,
		_w7026_
	);
	LUT4 #(
		.INIT('h9402)
	) name6993 (
		_w3772_,
		_w3881_,
		_w6953_,
		_w6956_,
		_w7027_
	);
	LUT4 #(
		.INIT('h2881)
	) name6994 (
		_w3883_,
		_w4025_,
		_w4027_,
		_w6952_,
		_w7028_
	);
	LUT3 #(
		.INIT('h56)
	) name6995 (
		_w4099_,
		_w4378_,
		_w6951_,
		_w7029_
	);
	LUT3 #(
		.INIT('h90)
	) name6996 (
		_w4030_,
		_w6952_,
		_w7029_,
		_w7030_
	);
	LUT4 #(
		.INIT('h4504)
	) name6997 (
		_w4379_,
		_w4453_,
		_w4454_,
		_w6947_,
		_w7031_
	);
	LUT4 #(
		.INIT('h6665)
	) name6998 (
		_w4379_,
		_w4455_,
		_w6947_,
		_w6948_,
		_w7032_
	);
	LUT4 #(
		.INIT('h8218)
	) name6999 (
		_w4099_,
		_w4376_,
		_w4377_,
		_w6950_,
		_w7033_
	);
	LUT4 #(
		.INIT('h8218)
	) name7000 (
		_w4379_,
		_w4453_,
		_w4454_,
		_w6947_,
		_w7034_
	);
	LUT3 #(
		.INIT('h1e)
	) name7001 (
		_w4695_,
		_w6944_,
		_w6946_,
		_w7035_
	);
	LUT3 #(
		.INIT('h90)
	) name7002 (
		_w6947_,
		_w6949_,
		_w7035_,
		_w7036_
	);
	LUT4 #(
		.INIT('h5110)
	) name7003 (
		_w4696_,
		_w4697_,
		_w4871_,
		_w6940_,
		_w7037_
	);
	LUT4 #(
		.INIT('h6665)
	) name7004 (
		_w4696_,
		_w4872_,
		_w6940_,
		_w6941_,
		_w7038_
	);
	LUT4 #(
		.INIT('h9204)
	) name7005 (
		_w4693_,
		_w4694_,
		_w6943_,
		_w6946_,
		_w7039_
	);
	LUT4 #(
		.INIT('h8224)
	) name7006 (
		_w4696_,
		_w4697_,
		_w4871_,
		_w6940_,
		_w7040_
	);
	LUT3 #(
		.INIT('h56)
	) name7007 (
		_w5067_,
		_w5282_,
		_w6939_,
		_w7041_
	);
	LUT3 #(
		.INIT('h90)
	) name7008 (
		_w6940_,
		_w6942_,
		_w7041_,
		_w7042_
	);
	LUT4 #(
		.INIT('h4504)
	) name7009 (
		_w5283_,
		_w5519_,
		_w5520_,
		_w6935_,
		_w7043_
	);
	LUT4 #(
		.INIT('h6665)
	) name7010 (
		_w5283_,
		_w5521_,
		_w6935_,
		_w6936_,
		_w7044_
	);
	LUT4 #(
		.INIT('h8218)
	) name7011 (
		_w5067_,
		_w5280_,
		_w5281_,
		_w6938_,
		_w7045_
	);
	LUT4 #(
		.INIT('h8218)
	) name7012 (
		_w5283_,
		_w5519_,
		_w5520_,
		_w6935_,
		_w7046_
	);
	LUT3 #(
		.INIT('h1e)
	) name7013 (
		_w6043_,
		_w6933_,
		_w6934_,
		_w7047_
	);
	LUT3 #(
		.INIT('h90)
	) name7014 (
		_w6935_,
		_w6937_,
		_w7047_,
		_w7048_
	);
	LUT4 #(
		.INIT('h4504)
	) name7015 (
		_w6044_,
		_w6328_,
		_w6329_,
		_w6929_,
		_w7049_
	);
	LUT4 #(
		.INIT('h6665)
	) name7016 (
		_w6044_,
		_w6330_,
		_w6929_,
		_w6930_,
		_w7050_
	);
	LUT4 #(
		.INIT('h9204)
	) name7017 (
		_w6040_,
		_w6042_,
		_w6932_,
		_w6934_,
		_w7051_
	);
	LUT4 #(
		.INIT('h8218)
	) name7018 (
		_w6044_,
		_w6328_,
		_w6329_,
		_w6929_,
		_w7052_
	);
	LUT3 #(
		.INIT('h1e)
	) name7019 (
		_w6645_,
		_w6926_,
		_w6928_,
		_w7053_
	);
	LUT3 #(
		.INIT('h90)
	) name7020 (
		_w6929_,
		_w6931_,
		_w7053_,
		_w7054_
	);
	LUT4 #(
		.INIT('h5110)
	) name7021 (
		_w6646_,
		_w6647_,
		_w6653_,
		_w6922_,
		_w7055_
	);
	LUT4 #(
		.INIT('h6665)
	) name7022 (
		_w6646_,
		_w6654_,
		_w6922_,
		_w6923_,
		_w7056_
	);
	LUT4 #(
		.INIT('h4182)
	) name7023 (
		_w6645_,
		_w6646_,
		_w6925_,
		_w6928_,
		_w7057_
	);
	LUT4 #(
		.INIT('h8224)
	) name7024 (
		_w6646_,
		_w6647_,
		_w6653_,
		_w6922_,
		_w7058_
	);
	LUT3 #(
		.INIT('h1e)
	) name7025 (
		_w6669_,
		_w6919_,
		_w6921_,
		_w7059_
	);
	LUT3 #(
		.INIT('h90)
	) name7026 (
		_w6922_,
		_w6924_,
		_w7059_,
		_w7060_
	);
	LUT4 #(
		.INIT('h00d4)
	) name7027 (
		_w6670_,
		_w6675_,
		_w6914_,
		_w6918_,
		_w7061_
	);
	LUT4 #(
		.INIT('h54ab)
	) name7028 (
		_w6676_,
		_w6914_,
		_w6915_,
		_w6918_,
		_w7062_
	);
	LUT4 #(
		.INIT('h9402)
	) name7029 (
		_w6662_,
		_w6668_,
		_w6917_,
		_w6921_,
		_w7063_
	);
	LUT4 #(
		.INIT('h2940)
	) name7030 (
		_w6662_,
		_w6668_,
		_w6917_,
		_w6921_,
		_w7064_
	);
	LUT4 #(
		.INIT('h1e2d)
	) name7031 (
		_w6669_,
		_w6919_,
		_w6921_,
		_w7061_,
		_w7065_
	);
	LUT2 #(
		.INIT('h9)
	) name7032 (
		_w6914_,
		_w6916_,
		_w7066_
	);
	LUT3 #(
		.INIT('he1)
	) name7033 (
		_w6689_,
		_w6911_,
		_w6913_,
		_w7067_
	);
	LUT3 #(
		.INIT('hc8)
	) name7034 (
		_w7062_,
		_w7066_,
		_w7067_,
		_w7068_
	);
	LUT3 #(
		.INIT('h45)
	) name7035 (
		_w7063_,
		_w7064_,
		_w7068_,
		_w7069_
	);
	LUT3 #(
		.INIT('h06)
	) name7036 (
		_w6922_,
		_w6924_,
		_w7059_,
		_w7070_
	);
	LUT3 #(
		.INIT('h69)
	) name7037 (
		_w6922_,
		_w6924_,
		_w7059_,
		_w7071_
	);
	LUT4 #(
		.INIT('h6959)
	) name7038 (
		_w6646_,
		_w6654_,
		_w6922_,
		_w6923_,
		_w7072_
	);
	LUT4 #(
		.INIT('hba00)
	) name7039 (
		_w7060_,
		_w7069_,
		_w7071_,
		_w7072_,
		_w7073_
	);
	LUT4 #(
		.INIT('h1e2d)
	) name7040 (
		_w6645_,
		_w6926_,
		_w6928_,
		_w7055_,
		_w7074_
	);
	LUT4 #(
		.INIT('h0155)
	) name7041 (
		_w7057_,
		_w7058_,
		_w7073_,
		_w7074_,
		_w7075_
	);
	LUT3 #(
		.INIT('h06)
	) name7042 (
		_w6929_,
		_w6931_,
		_w7053_,
		_w7076_
	);
	LUT3 #(
		.INIT('h69)
	) name7043 (
		_w6929_,
		_w6931_,
		_w7053_,
		_w7077_
	);
	LUT4 #(
		.INIT('h6959)
	) name7044 (
		_w6044_,
		_w6330_,
		_w6929_,
		_w6930_,
		_w7078_
	);
	LUT4 #(
		.INIT('hba00)
	) name7045 (
		_w7054_,
		_w7075_,
		_w7077_,
		_w7078_,
		_w7079_
	);
	LUT4 #(
		.INIT('h1e2d)
	) name7046 (
		_w6043_,
		_w6933_,
		_w6934_,
		_w7049_,
		_w7080_
	);
	LUT4 #(
		.INIT('h0155)
	) name7047 (
		_w7051_,
		_w7052_,
		_w7079_,
		_w7080_,
		_w7081_
	);
	LUT3 #(
		.INIT('h06)
	) name7048 (
		_w6935_,
		_w6937_,
		_w7047_,
		_w7082_
	);
	LUT3 #(
		.INIT('h69)
	) name7049 (
		_w6935_,
		_w6937_,
		_w7047_,
		_w7083_
	);
	LUT4 #(
		.INIT('h6959)
	) name7050 (
		_w5283_,
		_w5521_,
		_w6935_,
		_w6936_,
		_w7084_
	);
	LUT4 #(
		.INIT('hba00)
	) name7051 (
		_w7048_,
		_w7081_,
		_w7083_,
		_w7084_,
		_w7085_
	);
	LUT4 #(
		.INIT('h5659)
	) name7052 (
		_w5067_,
		_w5282_,
		_w6939_,
		_w7043_,
		_w7086_
	);
	LUT4 #(
		.INIT('h0155)
	) name7053 (
		_w7045_,
		_w7046_,
		_w7085_,
		_w7086_,
		_w7087_
	);
	LUT3 #(
		.INIT('h06)
	) name7054 (
		_w6940_,
		_w6942_,
		_w7041_,
		_w7088_
	);
	LUT3 #(
		.INIT('h69)
	) name7055 (
		_w6940_,
		_w6942_,
		_w7041_,
		_w7089_
	);
	LUT4 #(
		.INIT('h6959)
	) name7056 (
		_w4696_,
		_w4872_,
		_w6940_,
		_w6941_,
		_w7090_
	);
	LUT4 #(
		.INIT('hba00)
	) name7057 (
		_w7042_,
		_w7087_,
		_w7089_,
		_w7090_,
		_w7091_
	);
	LUT4 #(
		.INIT('h1e2d)
	) name7058 (
		_w4695_,
		_w6944_,
		_w6946_,
		_w7037_,
		_w7092_
	);
	LUT4 #(
		.INIT('h0155)
	) name7059 (
		_w7039_,
		_w7040_,
		_w7091_,
		_w7092_,
		_w7093_
	);
	LUT3 #(
		.INIT('h06)
	) name7060 (
		_w6947_,
		_w6949_,
		_w7035_,
		_w7094_
	);
	LUT3 #(
		.INIT('h69)
	) name7061 (
		_w6947_,
		_w6949_,
		_w7035_,
		_w7095_
	);
	LUT4 #(
		.INIT('h6959)
	) name7062 (
		_w4379_,
		_w4455_,
		_w6947_,
		_w6948_,
		_w7096_
	);
	LUT4 #(
		.INIT('hba00)
	) name7063 (
		_w7036_,
		_w7093_,
		_w7095_,
		_w7096_,
		_w7097_
	);
	LUT4 #(
		.INIT('h5659)
	) name7064 (
		_w4099_,
		_w4378_,
		_w6951_,
		_w7031_,
		_w7098_
	);
	LUT4 #(
		.INIT('h0155)
	) name7065 (
		_w7033_,
		_w7034_,
		_w7097_,
		_w7098_,
		_w7099_
	);
	LUT3 #(
		.INIT('h06)
	) name7066 (
		_w4030_,
		_w6952_,
		_w7029_,
		_w7100_
	);
	LUT3 #(
		.INIT('h69)
	) name7067 (
		_w4030_,
		_w6952_,
		_w7029_,
		_w7101_
	);
	LUT4 #(
		.INIT('h6599)
	) name7068 (
		_w3883_,
		_w4028_,
		_w4029_,
		_w6952_,
		_w7102_
	);
	LUT4 #(
		.INIT('hba00)
	) name7069 (
		_w7030_,
		_w7099_,
		_w7101_,
		_w7102_,
		_w7103_
	);
	LUT4 #(
		.INIT('h1e2d)
	) name7070 (
		_w3882_,
		_w6954_,
		_w6956_,
		_w7025_,
		_w7104_
	);
	LUT4 #(
		.INIT('h0155)
	) name7071 (
		_w7027_,
		_w7028_,
		_w7103_,
		_w7104_,
		_w7105_
	);
	LUT3 #(
		.INIT('h06)
	) name7072 (
		_w3706_,
		_w6957_,
		_w7023_,
		_w7106_
	);
	LUT3 #(
		.INIT('h69)
	) name7073 (
		_w3706_,
		_w6957_,
		_w7023_,
		_w7107_
	);
	LUT4 #(
		.INIT('h6599)
	) name7074 (
		_w3651_,
		_w3704_,
		_w3705_,
		_w6957_,
		_w7108_
	);
	LUT4 #(
		.INIT('hba00)
	) name7075 (
		_w7024_,
		_w7105_,
		_w7107_,
		_w7108_,
		_w7109_
	);
	LUT4 #(
		.INIT('h5659)
	) name7076 (
		_w3409_,
		_w3650_,
		_w6959_,
		_w7019_,
		_w7110_
	);
	LUT4 #(
		.INIT('h0155)
	) name7077 (
		_w7021_,
		_w7022_,
		_w7109_,
		_w7110_,
		_w7111_
	);
	LUT3 #(
		.INIT('h06)
	) name7078 (
		_w6960_,
		_w6962_,
		_w7017_,
		_w7112_
	);
	LUT3 #(
		.INIT('h69)
	) name7079 (
		_w6960_,
		_w6962_,
		_w7017_,
		_w7113_
	);
	LUT4 #(
		.INIT('h6959)
	) name7080 (
		_w3258_,
		_w3308_,
		_w6960_,
		_w6961_,
		_w7114_
	);
	LUT4 #(
		.INIT('hba00)
	) name7081 (
		_w7018_,
		_w7111_,
		_w7113_,
		_w7114_,
		_w7115_
	);
	LUT4 #(
		.INIT('h1e2d)
	) name7082 (
		_w3257_,
		_w6964_,
		_w6966_,
		_w7013_,
		_w7116_
	);
	LUT4 #(
		.INIT('h0155)
	) name7083 (
		_w7015_,
		_w7016_,
		_w7115_,
		_w7116_,
		_w7117_
	);
	LUT3 #(
		.INIT('h06)
	) name7084 (
		_w6967_,
		_w6969_,
		_w7011_,
		_w7118_
	);
	LUT3 #(
		.INIT('h69)
	) name7085 (
		_w6967_,
		_w6969_,
		_w7011_,
		_w7119_
	);
	LUT4 #(
		.INIT('h629d)
	) name7086 (
		_w3007_,
		_w6967_,
		_w6968_,
		_w6971_,
		_w7120_
	);
	LUT4 #(
		.INIT('hba00)
	) name7087 (
		_w7012_,
		_w7117_,
		_w7119_,
		_w7120_,
		_w7121_
	);
	LUT4 #(
		.INIT('h1e2d)
	) name7088 (
		_w2983_,
		_w6972_,
		_w6974_,
		_w7007_,
		_w7122_
	);
	LUT4 #(
		.INIT('h0155)
	) name7089 (
		_w7009_,
		_w7010_,
		_w7121_,
		_w7122_,
		_w7123_
	);
	LUT3 #(
		.INIT('h06)
	) name7090 (
		_w2872_,
		_w6975_,
		_w7005_,
		_w7124_
	);
	LUT3 #(
		.INIT('h69)
	) name7091 (
		_w2872_,
		_w6975_,
		_w7005_,
		_w7125_
	);
	LUT4 #(
		.INIT('h4ab5)
	) name7092 (
		_w2870_,
		_w2871_,
		_w6975_,
		_w6977_,
		_w7126_
	);
	LUT4 #(
		.INIT('hba00)
	) name7093 (
		_w7006_,
		_w7123_,
		_w7125_,
		_w7126_,
		_w7127_
	);
	LUT4 #(
		.INIT('h1e2d)
	) name7094 (
		_w2622_,
		_w6978_,
		_w6980_,
		_w7001_,
		_w7128_
	);
	LUT4 #(
		.INIT('h0155)
	) name7095 (
		_w7003_,
		_w7004_,
		_w7127_,
		_w7128_,
		_w7129_
	);
	LUT3 #(
		.INIT('h06)
	) name7096 (
		_w2546_,
		_w6981_,
		_w6999_,
		_w7130_
	);
	LUT3 #(
		.INIT('h69)
	) name7097 (
		_w2546_,
		_w6981_,
		_w6999_,
		_w7131_
	);
	LUT4 #(
		.INIT('h6599)
	) name7098 (
		_w2412_,
		_w2544_,
		_w2545_,
		_w6981_,
		_w7132_
	);
	LUT4 #(
		.INIT('hba00)
	) name7099 (
		_w7000_,
		_w7129_,
		_w7131_,
		_w7132_,
		_w7133_
	);
	LUT4 #(
		.INIT('h1e2d)
	) name7100 (
		_w2411_,
		_w6983_,
		_w6993_,
		_w6995_,
		_w7134_
	);
	LUT4 #(
		.INIT('h0155)
	) name7101 (
		_w6997_,
		_w6998_,
		_w7133_,
		_w7134_,
		_w7135_
	);
	LUT4 #(
		.INIT('h5501)
	) name7102 (
		_w6991_,
		_w2411_,
		_w6983_,
		_w6992_,
		_w7136_
	);
	LUT4 #(
		.INIT('h135f)
	) name7103 (
		_w65_,
		_w46_,
		_w158_,
		_w378_,
		_w7137_
	);
	LUT4 #(
		.INIT('h153f)
	) name7104 (
		_w52_,
		_w67_,
		_w419_,
		_w430_,
		_w7138_
	);
	LUT4 #(
		.INIT('h135f)
	) name7105 (
		_w52_,
		_w78_,
		_w39_,
		_w46_,
		_w7139_
	);
	LUT4 #(
		.INIT('h8000)
	) name7106 (
		_w198_,
		_w7139_,
		_w7137_,
		_w7138_,
		_w7140_
	);
	LUT4 #(
		.INIT('h153f)
	) name7107 (
		_w85_,
		_w67_,
		_w78_,
		_w201_,
		_w7141_
	);
	LUT4 #(
		.INIT('h1000)
	) name7108 (
		_w304_,
		_w264_,
		_w1169_,
		_w7141_,
		_w7142_
	);
	LUT4 #(
		.INIT('h135f)
	) name7109 (
		_w56_,
		_w41_,
		_w72_,
		_w236_,
		_w7143_
	);
	LUT3 #(
		.INIT('h40)
	) name7110 (
		_w180_,
		_w975_,
		_w7143_,
		_w7144_
	);
	LUT3 #(
		.INIT('h80)
	) name7111 (
		_w1673_,
		_w1726_,
		_w2116_,
		_w7145_
	);
	LUT4 #(
		.INIT('h8000)
	) name7112 (
		_w7144_,
		_w7145_,
		_w7140_,
		_w7142_,
		_w7146_
	);
	LUT2 #(
		.INIT('h8)
	) name7113 (
		_w2216_,
		_w7146_,
		_w7147_
	);
	LUT3 #(
		.INIT('h80)
	) name7114 (
		_w1569_,
		_w2566_,
		_w7147_,
		_w7148_
	);
	LUT4 #(
		.INIT('h135f)
	) name7115 (
		_w78_,
		_w56_,
		_w93_,
		_w158_,
		_w7149_
	);
	LUT3 #(
		.INIT('h80)
	) name7116 (
		_w1191_,
		_w2810_,
		_w7149_,
		_w7150_
	);
	LUT4 #(
		.INIT('h135f)
	) name7117 (
		_w110_,
		_w50_,
		_w184_,
		_w201_,
		_w7151_
	);
	LUT4 #(
		.INIT('h135f)
	) name7118 (
		_w56_,
		_w72_,
		_w39_,
		_w46_,
		_w7152_
	);
	LUT4 #(
		.INIT('h4000)
	) name7119 (
		_w468_,
		_w890_,
		_w7152_,
		_w7151_,
		_w7153_
	);
	LUT3 #(
		.INIT('h80)
	) name7120 (
		_w3046_,
		_w7150_,
		_w7153_,
		_w7154_
	);
	LUT3 #(
		.INIT('h80)
	) name7121 (
		_w944_,
		_w1154_,
		_w1362_,
		_w7155_
	);
	LUT4 #(
		.INIT('h153f)
	) name7122 (
		_w41_,
		_w39_,
		_w50_,
		_w419_,
		_w7156_
	);
	LUT4 #(
		.INIT('h8000)
	) name7123 (
		_w802_,
		_w772_,
		_w902_,
		_w7156_,
		_w7157_
	);
	LUT3 #(
		.INIT('h80)
	) name7124 (
		_w4205_,
		_w7155_,
		_w7157_,
		_w7158_
	);
	LUT4 #(
		.INIT('h4000)
	) name7125 (
		_w439_,
		_w832_,
		_w1852_,
		_w1853_,
		_w7159_
	);
	LUT4 #(
		.INIT('h8000)
	) name7126 (
		_w1597_,
		_w1599_,
		_w4229_,
		_w7159_,
		_w7160_
	);
	LUT3 #(
		.INIT('h80)
	) name7127 (
		_w7154_,
		_w7158_,
		_w7160_,
		_w7161_
	);
	LUT2 #(
		.INIT('h8)
	) name7128 (
		_w2588_,
		_w7161_,
		_w7162_
	);
	LUT2 #(
		.INIT('h8)
	) name7129 (
		_w7148_,
		_w7162_,
		_w7163_
	);
	LUT3 #(
		.INIT('h40)
	) name7130 (
		_w369_,
		_w357_,
		_w368_,
		_w7164_
	);
	LUT3 #(
		.INIT('h80)
	) name7131 (
		_w7148_,
		_w7162_,
		_w7164_,
		_w7165_
	);
	LUT2 #(
		.INIT('h1)
	) name7132 (
		_w6989_,
		_w7165_,
		_w7166_
	);
	LUT2 #(
		.INIT('h8)
	) name7133 (
		_w6989_,
		_w7165_,
		_w7167_
	);
	LUT2 #(
		.INIT('h6)
	) name7134 (
		_w6989_,
		_w7165_,
		_w7168_
	);
	LUT2 #(
		.INIT('h9)
	) name7135 (
		_w7136_,
		_w7168_,
		_w7169_
	);
	LUT3 #(
		.INIT('h48)
	) name7136 (
		_w7136_,
		_w6994_,
		_w7168_,
		_w7170_
	);
	LUT3 #(
		.INIT('h21)
	) name7137 (
		_w7136_,
		_w6994_,
		_w7168_,
		_w7171_
	);
	LUT3 #(
		.INIT('h96)
	) name7138 (
		_w7136_,
		_w6994_,
		_w7168_,
		_w7172_
	);
	LUT3 #(
		.INIT('h82)
	) name7139 (
		_w37_,
		_w7135_,
		_w7172_,
		_w7173_
	);
	LUT3 #(
		.INIT('h28)
	) name7140 (
		_w3262_,
		_w7136_,
		_w7168_,
		_w7174_
	);
	LUT2 #(
		.INIT('h8)
	) name7141 (
		_w3214_,
		_w6996_,
		_w7175_
	);
	LUT4 #(
		.INIT('h04c8)
	) name7142 (
		_w2411_,
		_w3249_,
		_w6983_,
		_w6993_,
		_w7176_
	);
	LUT2 #(
		.INIT('h1)
	) name7143 (
		_w7175_,
		_w7176_,
		_w7177_
	);
	LUT2 #(
		.INIT('h4)
	) name7144 (
		_w7174_,
		_w7177_,
		_w7178_
	);
	LUT3 #(
		.INIT('h9a)
	) name7145 (
		\a[23] ,
		_w7173_,
		_w7178_,
		_w7179_
	);
	LUT3 #(
		.INIT('h82)
	) name7146 (
		_w2875_,
		_w7129_,
		_w7131_,
		_w7180_
	);
	LUT3 #(
		.INIT('h84)
	) name7147 (
		_w2546_,
		_w2986_,
		_w6981_,
		_w7181_
	);
	LUT2 #(
		.INIT('h8)
	) name7148 (
		_w2874_,
		_w7002_,
		_w7182_
	);
	LUT4 #(
		.INIT('h04c8)
	) name7149 (
		_w2622_,
		_w2975_,
		_w6978_,
		_w6980_,
		_w7183_
	);
	LUT2 #(
		.INIT('h1)
	) name7150 (
		_w7182_,
		_w7183_,
		_w7184_
	);
	LUT2 #(
		.INIT('h4)
	) name7151 (
		_w7181_,
		_w7184_,
		_w7185_
	);
	LUT3 #(
		.INIT('h9a)
	) name7152 (
		\a[26] ,
		_w7180_,
		_w7185_,
		_w7186_
	);
	LUT3 #(
		.INIT('h80)
	) name7153 (
		_w1754_,
		_w1844_,
		_w3037_,
		_w7187_
	);
	LUT4 #(
		.INIT('h135f)
	) name7154 (
		_w52_,
		_w46_,
		_w236_,
		_w166_,
		_w7188_
	);
	LUT4 #(
		.INIT('h8000)
	) name7155 (
		_w472_,
		_w1537_,
		_w4133_,
		_w7188_,
		_w7189_
	);
	LUT2 #(
		.INIT('h8)
	) name7156 (
		_w7187_,
		_w7189_,
		_w7190_
	);
	LUT3 #(
		.INIT('h40)
	) name7157 (
		_w454_,
		_w566_,
		_w696_,
		_w7191_
	);
	LUT4 #(
		.INIT('h0777)
	) name7158 (
		_w78_,
		_w56_,
		_w41_,
		_w201_,
		_w7192_
	);
	LUT4 #(
		.INIT('h4000)
	) name7159 (
		_w159_,
		_w1878_,
		_w2397_,
		_w7192_,
		_w7193_
	);
	LUT4 #(
		.INIT('h8000)
	) name7160 (
		_w2087_,
		_w3429_,
		_w7193_,
		_w7191_,
		_w7194_
	);
	LUT2 #(
		.INIT('h8)
	) name7161 (
		_w7190_,
		_w7194_,
		_w7195_
	);
	LUT4 #(
		.INIT('h0777)
	) name7162 (
		_w38_,
		_w106_,
		_w59_,
		_w72_,
		_w7196_
	);
	LUT4 #(
		.INIT('h153f)
	) name7163 (
		_w38_,
		_w110_,
		_w43_,
		_w184_,
		_w7197_
	);
	LUT3 #(
		.INIT('h40)
	) name7164 (
		_w406_,
		_w7196_,
		_w7197_,
		_w7198_
	);
	LUT2 #(
		.INIT('h4)
	) name7165 (
		_w227_,
		_w1635_,
		_w7199_
	);
	LUT4 #(
		.INIT('h4000)
	) name7166 (
		_w429_,
		_w976_,
		_w2654_,
		_w3125_,
		_w7200_
	);
	LUT3 #(
		.INIT('h80)
	) name7167 (
		_w7199_,
		_w7198_,
		_w7200_,
		_w7201_
	);
	LUT4 #(
		.INIT('h135f)
	) name7168 (
		_w67_,
		_w90_,
		_w236_,
		_w378_,
		_w7202_
	);
	LUT2 #(
		.INIT('h4)
	) name7169 (
		_w478_,
		_w7202_,
		_w7203_
	);
	LUT3 #(
		.INIT('h40)
	) name7170 (
		_w141_,
		_w1472_,
		_w2209_,
		_w7204_
	);
	LUT2 #(
		.INIT('h8)
	) name7171 (
		_w7203_,
		_w7204_,
		_w7205_
	);
	LUT4 #(
		.INIT('h135f)
	) name7172 (
		_w47_,
		_w65_,
		_w184_,
		_w158_,
		_w7206_
	);
	LUT4 #(
		.INIT('h135f)
	) name7173 (
		_w55_,
		_w52_,
		_w236_,
		_w419_,
		_w7207_
	);
	LUT4 #(
		.INIT('h8000)
	) name7174 (
		_w867_,
		_w1080_,
		_w7206_,
		_w7207_,
		_w7208_
	);
	LUT4 #(
		.INIT('h0777)
	) name7175 (
		_w38_,
		_w122_,
		_w59_,
		_w184_,
		_w7209_
	);
	LUT4 #(
		.INIT('h135f)
	) name7176 (
		_w110_,
		_w47_,
		_w236_,
		_w430_,
		_w7210_
	);
	LUT4 #(
		.INIT('h153f)
	) name7177 (
		_w47_,
		_w46_,
		_w236_,
		_w176_,
		_w7211_
	);
	LUT3 #(
		.INIT('h37)
	) name7178 (
		_w122_,
		_w44_,
		_w166_,
		_w7212_
	);
	LUT4 #(
		.INIT('h8000)
	) name7179 (
		_w7211_,
		_w7212_,
		_w7209_,
		_w7210_,
		_w7213_
	);
	LUT3 #(
		.INIT('h80)
	) name7180 (
		_w1360_,
		_w1423_,
		_w2126_,
		_w7214_
	);
	LUT4 #(
		.INIT('h8000)
	) name7181 (
		_w3110_,
		_w7213_,
		_w7214_,
		_w7208_,
		_w7215_
	);
	LUT3 #(
		.INIT('h80)
	) name7182 (
		_w7201_,
		_w7205_,
		_w7215_,
		_w7216_
	);
	LUT3 #(
		.INIT('h80)
	) name7183 (
		_w2183_,
		_w7195_,
		_w7216_,
		_w7217_
	);
	LUT4 #(
		.INIT('h135f)
	) name7184 (
		_w55_,
		_w110_,
		_w78_,
		_w201_,
		_w7218_
	);
	LUT4 #(
		.INIT('h8000)
	) name7185 (
		_w873_,
		_w2170_,
		_w2256_,
		_w7218_,
		_w7219_
	);
	LUT4 #(
		.INIT('h135f)
	) name7186 (
		_w55_,
		_w110_,
		_w236_,
		_w166_,
		_w7220_
	);
	LUT4 #(
		.INIT('h153f)
	) name7187 (
		_w55_,
		_w41_,
		_w72_,
		_w166_,
		_w7221_
	);
	LUT4 #(
		.INIT('h8000)
	) name7188 (
		_w1165_,
		_w2468_,
		_w7220_,
		_w7221_,
		_w7222_
	);
	LUT4 #(
		.INIT('h8000)
	) name7189 (
		_w521_,
		_w767_,
		_w856_,
		_w1043_,
		_w7223_
	);
	LUT3 #(
		.INIT('h80)
	) name7190 (
		_w7219_,
		_w7222_,
		_w7223_,
		_w7224_
	);
	LUT3 #(
		.INIT('h1f)
	) name7191 (
		_w55_,
		_w50_,
		_w43_,
		_w7225_
	);
	LUT4 #(
		.INIT('h2000)
	) name7192 (
		_w292_,
		_w160_,
		_w1490_,
		_w7225_,
		_w7226_
	);
	LUT4 #(
		.INIT('h8000)
	) name7193 (
		_w2108_,
		_w3564_,
		_w3569_,
		_w7226_,
		_w7227_
	);
	LUT4 #(
		.INIT('h8000)
	) name7194 (
		_w2043_,
		_w2054_,
		_w7224_,
		_w7227_,
		_w7228_
	);
	LUT2 #(
		.INIT('h8)
	) name7195 (
		_w2775_,
		_w7228_,
		_w7229_
	);
	LUT4 #(
		.INIT('h153f)
	) name7196 (
		_w52_,
		_w59_,
		_w78_,
		_w72_,
		_w7230_
	);
	LUT2 #(
		.INIT('h8)
	) name7197 (
		_w2234_,
		_w7230_,
		_w7231_
	);
	LUT4 #(
		.INIT('h153f)
	) name7198 (
		_w50_,
		_w43_,
		_w93_,
		_w158_,
		_w7232_
	);
	LUT2 #(
		.INIT('h8)
	) name7199 (
		_w252_,
		_w7232_,
		_w7233_
	);
	LUT4 #(
		.INIT('h8000)
	) name7200 (
		_w252_,
		_w265_,
		_w4225_,
		_w7232_,
		_w7234_
	);
	LUT4 #(
		.INIT('h8000)
	) name7201 (
		_w54_,
		_w1514_,
		_w2517_,
		_w3561_,
		_w7235_
	);
	LUT4 #(
		.INIT('h153f)
	) name7202 (
		_w41_,
		_w46_,
		_w166_,
		_w176_,
		_w7236_
	);
	LUT4 #(
		.INIT('h0777)
	) name7203 (
		_w106_,
		_w90_,
		_w50_,
		_w430_,
		_w7237_
	);
	LUT4 #(
		.INIT('h4000)
	) name7204 (
		_w224_,
		_w555_,
		_w7236_,
		_w7237_,
		_w7238_
	);
	LUT4 #(
		.INIT('h8000)
	) name7205 (
		_w7231_,
		_w7235_,
		_w7238_,
		_w7234_,
		_w7239_
	);
	LUT3 #(
		.INIT('h80)
	) name7206 (
		_w2165_,
		_w7201_,
		_w7239_,
		_w7240_
	);
	LUT3 #(
		.INIT('h80)
	) name7207 (
		_w2389_,
		_w3354_,
		_w3356_,
		_w7241_
	);
	LUT2 #(
		.INIT('h8)
	) name7208 (
		_w7240_,
		_w7241_,
		_w7242_
	);
	LUT4 #(
		.INIT('h0777)
	) name7209 (
		_w2775_,
		_w7228_,
		_w7240_,
		_w7241_,
		_w7243_
	);
	LUT2 #(
		.INIT('h4)
	) name7210 (
		_w7136_,
		_w7166_,
		_w7244_
	);
	LUT4 #(
		.INIT('h8001)
	) name7211 (
		\a[14] ,
		\a[15] ,
		\a[16] ,
		\a[17] ,
		_w7245_
	);
	LUT4 #(
		.INIT('h559a)
	) name7212 (
		\a[17] ,
		_w7136_,
		_w7166_,
		_w7245_,
		_w7246_
	);
	LUT4 #(
		.INIT('h8000)
	) name7213 (
		_w2775_,
		_w7228_,
		_w7240_,
		_w7241_,
		_w7247_
	);
	LUT4 #(
		.INIT('h7888)
	) name7214 (
		_w2775_,
		_w7228_,
		_w7240_,
		_w7241_,
		_w7248_
	);
	LUT3 #(
		.INIT('h51)
	) name7215 (
		_w7243_,
		_w7246_,
		_w7247_,
		_w7249_
	);
	LUT4 #(
		.INIT('h2a02)
	) name7216 (
		_w7217_,
		_w7229_,
		_w7242_,
		_w7246_,
		_w7250_
	);
	LUT4 #(
		.INIT('h4054)
	) name7217 (
		_w7217_,
		_w7229_,
		_w7242_,
		_w7246_,
		_w7251_
	);
	LUT4 #(
		.INIT('h6656)
	) name7218 (
		_w7217_,
		_w7243_,
		_w7246_,
		_w7247_,
		_w7252_
	);
	LUT4 #(
		.INIT('h02a8)
	) name7219 (
		_w377_,
		_w7016_,
		_w7115_,
		_w7116_,
		_w7253_
	);
	LUT4 #(
		.INIT('h02a8)
	) name7220 (
		_w2527_,
		_w3257_,
		_w6964_,
		_w6966_,
		_w7254_
	);
	LUT3 #(
		.INIT('h82)
	) name7221 (
		_w376_,
		_w6960_,
		_w6962_,
		_w7255_
	);
	LUT3 #(
		.INIT('h07)
	) name7222 (
		_w2407_,
		_w7014_,
		_w7255_,
		_w7256_
	);
	LUT2 #(
		.INIT('h4)
	) name7223 (
		_w7254_,
		_w7256_,
		_w7257_
	);
	LUT2 #(
		.INIT('h4)
	) name7224 (
		_w7253_,
		_w7257_,
		_w7258_
	);
	LUT4 #(
		.INIT('h153f)
	) name7225 (
		_w52_,
		_w59_,
		_w39_,
		_w236_,
		_w7259_
	);
	LUT4 #(
		.INIT('h2000)
	) name7226 (
		_w219_,
		_w347_,
		_w512_,
		_w7259_,
		_w7260_
	);
	LUT4 #(
		.INIT('h4000)
	) name7227 (
		_w359_,
		_w863_,
		_w1401_,
		_w3132_,
		_w7261_
	);
	LUT2 #(
		.INIT('h8)
	) name7228 (
		_w7260_,
		_w7261_,
		_w7262_
	);
	LUT4 #(
		.INIT('h135f)
	) name7229 (
		_w106_,
		_w85_,
		_w56_,
		_w378_,
		_w7263_
	);
	LUT3 #(
		.INIT('h40)
	) name7230 (
		_w435_,
		_w1800_,
		_w7263_,
		_w7264_
	);
	LUT4 #(
		.INIT('h153f)
	) name7231 (
		_w59_,
		_w41_,
		_w166_,
		_w176_,
		_w7265_
	);
	LUT4 #(
		.INIT('h8000)
	) name7232 (
		_w788_,
		_w1576_,
		_w2431_,
		_w7265_,
		_w7266_
	);
	LUT3 #(
		.INIT('h80)
	) name7233 (
		_w1389_,
		_w7264_,
		_w7266_,
		_w7267_
	);
	LUT3 #(
		.INIT('h80)
	) name7234 (
		_w1823_,
		_w7262_,
		_w7267_,
		_w7268_
	);
	LUT4 #(
		.INIT('h8000)
	) name7235 (
		_w676_,
		_w1173_,
		_w1318_,
		_w1726_,
		_w7269_
	);
	LUT3 #(
		.INIT('h57)
	) name7236 (
		_w93_,
		_w166_,
		_w176_,
		_w7270_
	);
	LUT4 #(
		.INIT('h153f)
	) name7237 (
		_w56_,
		_w65_,
		_w236_,
		_w259_,
		_w7271_
	);
	LUT4 #(
		.INIT('h0777)
	) name7238 (
		_w90_,
		_w39_,
		_w43_,
		_w65_,
		_w7272_
	);
	LUT3 #(
		.INIT('h1f)
	) name7239 (
		_w38_,
		_w93_,
		_w201_,
		_w7273_
	);
	LUT4 #(
		.INIT('h8000)
	) name7240 (
		_w7272_,
		_w7273_,
		_w7270_,
		_w7271_,
		_w7274_
	);
	LUT4 #(
		.INIT('h4000)
	) name7241 (
		_w437_,
		_w828_,
		_w829_,
		_w2267_,
		_w7275_
	);
	LUT3 #(
		.INIT('h80)
	) name7242 (
		_w7269_,
		_w7274_,
		_w7275_,
		_w7276_
	);
	LUT4 #(
		.INIT('h8000)
	) name7243 (
		_w1830_,
		_w3537_,
		_w3548_,
		_w7276_,
		_w7277_
	);
	LUT2 #(
		.INIT('h8)
	) name7244 (
		_w7268_,
		_w7277_,
		_w7278_
	);
	LUT2 #(
		.INIT('h2)
	) name7245 (
		_w7217_,
		_w7278_,
		_w7279_
	);
	LUT2 #(
		.INIT('h4)
	) name7246 (
		_w7217_,
		_w7278_,
		_w7280_
	);
	LUT2 #(
		.INIT('h9)
	) name7247 (
		_w7217_,
		_w7278_,
		_w7281_
	);
	LUT3 #(
		.INIT('h82)
	) name7248 (
		_w377_,
		_w7117_,
		_w7119_,
		_w7282_
	);
	LUT3 #(
		.INIT('h82)
	) name7249 (
		_w2527_,
		_w6967_,
		_w6969_,
		_w7283_
	);
	LUT2 #(
		.INIT('h8)
	) name7250 (
		_w376_,
		_w7014_,
		_w7284_
	);
	LUT4 #(
		.INIT('h02a8)
	) name7251 (
		_w2407_,
		_w3257_,
		_w6964_,
		_w6966_,
		_w7285_
	);
	LUT2 #(
		.INIT('h1)
	) name7252 (
		_w7284_,
		_w7285_,
		_w7286_
	);
	LUT2 #(
		.INIT('h4)
	) name7253 (
		_w7283_,
		_w7286_,
		_w7287_
	);
	LUT3 #(
		.INIT('h65)
	) name7254 (
		_w7281_,
		_w7282_,
		_w7287_,
		_w7288_
	);
	LUT4 #(
		.INIT('h2b00)
	) name7255 (
		_w7217_,
		_w7249_,
		_w7258_,
		_w7288_,
		_w7289_
	);
	LUT4 #(
		.INIT('h54ab)
	) name7256 (
		_w7250_,
		_w7251_,
		_w7258_,
		_w7288_,
		_w7290_
	);
	LUT4 #(
		.INIT('h54ab)
	) name7257 (
		_w7018_,
		_w7111_,
		_w7112_,
		_w7114_,
		_w7291_
	);
	LUT4 #(
		.INIT('h2228)
	) name7258 (
		_w376_,
		_w3409_,
		_w3650_,
		_w6959_,
		_w7292_
	);
	LUT4 #(
		.INIT('h007d)
	) name7259 (
		_w2407_,
		_w6960_,
		_w6962_,
		_w7292_,
		_w7293_
	);
	LUT3 #(
		.INIT('h70)
	) name7260 (
		_w2527_,
		_w7014_,
		_w7293_,
		_w7294_
	);
	LUT3 #(
		.INIT('h70)
	) name7261 (
		_w377_,
		_w7291_,
		_w7294_,
		_w7295_
	);
	LUT3 #(
		.INIT('h06)
	) name7262 (
		_w7246_,
		_w7248_,
		_w7295_,
		_w7296_
	);
	LUT4 #(
		.INIT('h135f)
	) name7263 (
		_w110_,
		_w67_,
		_w78_,
		_w176_,
		_w7297_
	);
	LUT3 #(
		.INIT('h80)
	) name7264 (
		_w2809_,
		_w3335_,
		_w7297_,
		_w7298_
	);
	LUT4 #(
		.INIT('h153f)
	) name7265 (
		_w90_,
		_w47_,
		_w43_,
		_w201_,
		_w7299_
	);
	LUT4 #(
		.INIT('h153f)
	) name7266 (
		_w50_,
		_w46_,
		_w184_,
		_w378_,
		_w7300_
	);
	LUT4 #(
		.INIT('h8000)
	) name7267 (
		_w1519_,
		_w2280_,
		_w7299_,
		_w7300_,
		_w7301_
	);
	LUT4 #(
		.INIT('h153f)
	) name7268 (
		_w47_,
		_w93_,
		_w236_,
		_w259_,
		_w7302_
	);
	LUT4 #(
		.INIT('h153f)
	) name7269 (
		_w59_,
		_w46_,
		_w419_,
		_w430_,
		_w7303_
	);
	LUT3 #(
		.INIT('h80)
	) name7270 (
		_w535_,
		_w7302_,
		_w7303_,
		_w7304_
	);
	LUT4 #(
		.INIT('h8000)
	) name7271 (
		_w3919_,
		_w7304_,
		_w7298_,
		_w7301_,
		_w7305_
	);
	LUT2 #(
		.INIT('h8)
	) name7272 (
		_w3124_,
		_w7305_,
		_w7306_
	);
	LUT2 #(
		.INIT('h4)
	) name7273 (
		_w432_,
		_w2267_,
		_w7307_
	);
	LUT3 #(
		.INIT('h80)
	) name7274 (
		_w3124_,
		_w7305_,
		_w7307_,
		_w7308_
	);
	LUT4 #(
		.INIT('h8000)
	) name7275 (
		_w942_,
		_w975_,
		_w2112_,
		_w7221_,
		_w7309_
	);
	LUT4 #(
		.INIT('h0777)
	) name7276 (
		_w122_,
		_w67_,
		_w41_,
		_w201_,
		_w7310_
	);
	LUT4 #(
		.INIT('h135f)
	) name7277 (
		_w38_,
		_w44_,
		_w419_,
		_w430_,
		_w7311_
	);
	LUT4 #(
		.INIT('h4000)
	) name7278 (
		_w107_,
		_w876_,
		_w7310_,
		_w7311_,
		_w7312_
	);
	LUT2 #(
		.INIT('h8)
	) name7279 (
		_w7309_,
		_w7312_,
		_w7313_
	);
	LUT4 #(
		.INIT('h0777)
	) name7280 (
		_w122_,
		_w90_,
		_w39_,
		_w65_,
		_w7314_
	);
	LUT4 #(
		.INIT('h1000)
	) name7281 (
		_w160_,
		_w385_,
		_w1442_,
		_w7314_,
		_w7315_
	);
	LUT2 #(
		.INIT('h8)
	) name7282 (
		_w2117_,
		_w3561_,
		_w7316_
	);
	LUT4 #(
		.INIT('h4000)
	) name7283 (
		_w455_,
		_w1806_,
		_w2117_,
		_w3561_,
		_w7317_
	);
	LUT3 #(
		.INIT('h57)
	) name7284 (
		_w59_,
		_w43_,
		_w236_,
		_w7318_
	);
	LUT4 #(
		.INIT('h8000)
	) name7285 (
		_w496_,
		_w1318_,
		_w3087_,
		_w7318_,
		_w7319_
	);
	LUT4 #(
		.INIT('h8000)
	) name7286 (
		_w2462_,
		_w7319_,
		_w7315_,
		_w7317_,
		_w7320_
	);
	LUT4 #(
		.INIT('h8000)
	) name7287 (
		_w2216_,
		_w2227_,
		_w7313_,
		_w7320_,
		_w7321_
	);
	LUT2 #(
		.INIT('h8)
	) name7288 (
		_w7308_,
		_w7321_,
		_w7322_
	);
	LUT4 #(
		.INIT('h135f)
	) name7289 (
		_w56_,
		_w50_,
		_w201_,
		_w430_,
		_w7323_
	);
	LUT3 #(
		.INIT('h80)
	) name7290 (
		_w3462_,
		_w3471_,
		_w7323_,
		_w7324_
	);
	LUT4 #(
		.INIT('h0777)
	) name7291 (
		_w72_,
		_w93_,
		_w46_,
		_w419_,
		_w7325_
	);
	LUT4 #(
		.INIT('h153f)
	) name7292 (
		_w85_,
		_w78_,
		_w90_,
		_w236_,
		_w7326_
	);
	LUT4 #(
		.INIT('h8000)
	) name7293 (
		_w560_,
		_w2510_,
		_w7325_,
		_w7326_,
		_w7327_
	);
	LUT4 #(
		.INIT('h0777)
	) name7294 (
		_w59_,
		_w39_,
		_w50_,
		_w184_,
		_w7328_
	);
	LUT4 #(
		.INIT('h8000)
	) name7295 (
		_w54_,
		_w518_,
		_w3573_,
		_w7328_,
		_w7329_
	);
	LUT4 #(
		.INIT('h8000)
	) name7296 (
		_w1338_,
		_w1343_,
		_w7327_,
		_w7329_,
		_w7330_
	);
	LUT4 #(
		.INIT('h8000)
	) name7297 (
		_w813_,
		_w827_,
		_w2287_,
		_w7330_,
		_w7331_
	);
	LUT2 #(
		.INIT('h8)
	) name7298 (
		_w7324_,
		_w7331_,
		_w7332_
	);
	LUT3 #(
		.INIT('h1f)
	) name7299 (
		_w110_,
		_w93_,
		_w158_,
		_w7333_
	);
	LUT4 #(
		.INIT('h153f)
	) name7300 (
		_w38_,
		_w122_,
		_w52_,
		_w201_,
		_w7334_
	);
	LUT4 #(
		.INIT('h4000)
	) name7301 (
		_w389_,
		_w1556_,
		_w7334_,
		_w7333_,
		_w7335_
	);
	LUT3 #(
		.INIT('h37)
	) name7302 (
		_w122_,
		_w110_,
		_w419_,
		_w7336_
	);
	LUT4 #(
		.INIT('h135f)
	) name7303 (
		_w106_,
		_w59_,
		_w41_,
		_w176_,
		_w7337_
	);
	LUT4 #(
		.INIT('h8000)
	) name7304 (
		_w997_,
		_w1519_,
		_w7337_,
		_w7336_,
		_w7338_
	);
	LUT4 #(
		.INIT('h8000)
	) name7305 (
		_w987_,
		_w2738_,
		_w7338_,
		_w7335_,
		_w7339_
	);
	LUT2 #(
		.INIT('h8)
	) name7306 (
		_w650_,
		_w1184_,
		_w7340_
	);
	LUT4 #(
		.INIT('h8000)
	) name7307 (
		_w1180_,
		_w1434_,
		_w1475_,
		_w3107_,
		_w7341_
	);
	LUT4 #(
		.INIT('h8000)
	) name7308 (
		_w1727_,
		_w1730_,
		_w7340_,
		_w7341_,
		_w7342_
	);
	LUT4 #(
		.INIT('h8000)
	) name7309 (
		_w1261_,
		_w1750_,
		_w7339_,
		_w7342_,
		_w7343_
	);
	LUT2 #(
		.INIT('h8)
	) name7310 (
		_w4148_,
		_w7343_,
		_w7344_
	);
	LUT4 #(
		.INIT('h153f)
	) name7311 (
		_w4148_,
		_w7324_,
		_w7331_,
		_w7343_,
		_w7345_
	);
	LUT4 #(
		.INIT('h8001)
	) name7312 (
		\a[11] ,
		\a[12] ,
		\a[13] ,
		\a[14] ,
		_w7346_
	);
	LUT4 #(
		.INIT('h559a)
	) name7313 (
		\a[14] ,
		_w7136_,
		_w7166_,
		_w7346_,
		_w7347_
	);
	LUT4 #(
		.INIT('h8000)
	) name7314 (
		_w4148_,
		_w7324_,
		_w7331_,
		_w7343_,
		_w7348_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name7315 (
		_w4148_,
		_w7324_,
		_w7331_,
		_w7343_,
		_w7349_
	);
	LUT3 #(
		.INIT('h51)
	) name7316 (
		_w7345_,
		_w7347_,
		_w7348_,
		_w7350_
	);
	LUT4 #(
		.INIT('h2a02)
	) name7317 (
		_w7322_,
		_w7332_,
		_w7344_,
		_w7347_,
		_w7351_
	);
	LUT4 #(
		.INIT('h4054)
	) name7318 (
		_w7322_,
		_w7332_,
		_w7344_,
		_w7347_,
		_w7352_
	);
	LUT4 #(
		.INIT('h6656)
	) name7319 (
		_w7322_,
		_w7345_,
		_w7347_,
		_w7348_,
		_w7353_
	);
	LUT4 #(
		.INIT('h02a8)
	) name7320 (
		_w377_,
		_w7022_,
		_w7109_,
		_w7110_,
		_w7354_
	);
	LUT4 #(
		.INIT('h2228)
	) name7321 (
		_w2527_,
		_w3409_,
		_w3650_,
		_w6959_,
		_w7355_
	);
	LUT3 #(
		.INIT('h82)
	) name7322 (
		_w376_,
		_w3706_,
		_w6957_,
		_w7356_
	);
	LUT3 #(
		.INIT('h07)
	) name7323 (
		_w2407_,
		_w7020_,
		_w7356_,
		_w7357_
	);
	LUT2 #(
		.INIT('h4)
	) name7324 (
		_w7355_,
		_w7357_,
		_w7358_
	);
	LUT2 #(
		.INIT('h4)
	) name7325 (
		_w7354_,
		_w7358_,
		_w7359_
	);
	LUT4 #(
		.INIT('h8777)
	) name7326 (
		_w2775_,
		_w7228_,
		_w7308_,
		_w7321_,
		_w7360_
	);
	LUT4 #(
		.INIT('hd554)
	) name7327 (
		_w7229_,
		_w7322_,
		_w7350_,
		_w7359_,
		_w7361_
	);
	LUT3 #(
		.INIT('h90)
	) name7328 (
		_w7246_,
		_w7248_,
		_w7295_,
		_w7362_
	);
	LUT3 #(
		.INIT('h69)
	) name7329 (
		_w7246_,
		_w7248_,
		_w7295_,
		_w7363_
	);
	LUT3 #(
		.INIT('h54)
	) name7330 (
		_w7296_,
		_w7361_,
		_w7362_,
		_w7364_
	);
	LUT2 #(
		.INIT('h9)
	) name7331 (
		_w7252_,
		_w7258_,
		_w7365_
	);
	LUT4 #(
		.INIT('hba00)
	) name7332 (
		_w7296_,
		_w7361_,
		_w7363_,
		_w7365_,
		_w7366_
	);
	LUT4 #(
		.INIT('h0045)
	) name7333 (
		_w7296_,
		_w7361_,
		_w7363_,
		_w7365_,
		_w7367_
	);
	LUT4 #(
		.INIT('h54ab)
	) name7334 (
		_w7296_,
		_w7361_,
		_w7362_,
		_w7365_,
		_w7368_
	);
	LUT4 #(
		.INIT('h02a8)
	) name7335 (
		_w2550_,
		_w7010_,
		_w7121_,
		_w7122_,
		_w7369_
	);
	LUT4 #(
		.INIT('h02a8)
	) name7336 (
		_w2854_,
		_w2983_,
		_w6972_,
		_w6974_,
		_w7370_
	);
	LUT3 #(
		.INIT('h82)
	) name7337 (
		_w2549_,
		_w6967_,
		_w6969_,
		_w7371_
	);
	LUT3 #(
		.INIT('h07)
	) name7338 (
		_w2617_,
		_w7008_,
		_w7371_,
		_w7372_
	);
	LUT2 #(
		.INIT('h4)
	) name7339 (
		_w7370_,
		_w7372_,
		_w7373_
	);
	LUT3 #(
		.INIT('h9a)
	) name7340 (
		\a[29] ,
		_w7369_,
		_w7373_,
		_w7374_
	);
	LUT4 #(
		.INIT('h20a2)
	) name7341 (
		_w7290_,
		_w7364_,
		_w7365_,
		_w7374_,
		_w7375_
	);
	LUT4 #(
		.INIT('h6665)
	) name7342 (
		_w7290_,
		_w7366_,
		_w7367_,
		_w7374_,
		_w7376_
	);
	LUT3 #(
		.INIT('h82)
	) name7343 (
		_w2550_,
		_w7123_,
		_w7125_,
		_w7377_
	);
	LUT3 #(
		.INIT('h82)
	) name7344 (
		_w2854_,
		_w2872_,
		_w6975_,
		_w7378_
	);
	LUT2 #(
		.INIT('h8)
	) name7345 (
		_w2549_,
		_w7008_,
		_w7379_
	);
	LUT4 #(
		.INIT('h02a8)
	) name7346 (
		_w2617_,
		_w2983_,
		_w6972_,
		_w6974_,
		_w7380_
	);
	LUT2 #(
		.INIT('h1)
	) name7347 (
		_w7379_,
		_w7380_,
		_w7381_
	);
	LUT2 #(
		.INIT('h4)
	) name7348 (
		_w7378_,
		_w7381_,
		_w7382_
	);
	LUT3 #(
		.INIT('h9a)
	) name7349 (
		\a[29] ,
		_w7377_,
		_w7382_,
		_w7383_
	);
	LUT3 #(
		.INIT('h96)
	) name7350 (
		_w7376_,
		_w7383_,
		_w7186_,
		_w7384_
	);
	LUT2 #(
		.INIT('h9)
	) name7351 (
		_w7368_,
		_w7374_,
		_w7385_
	);
	LUT4 #(
		.INIT('h54ab)
	) name7352 (
		_w7351_,
		_w7352_,
		_w7359_,
		_w7360_,
		_w7386_
	);
	LUT3 #(
		.INIT('h82)
	) name7353 (
		_w377_,
		_w7111_,
		_w7113_,
		_w7387_
	);
	LUT3 #(
		.INIT('h82)
	) name7354 (
		_w2527_,
		_w6960_,
		_w6962_,
		_w7388_
	);
	LUT2 #(
		.INIT('h8)
	) name7355 (
		_w376_,
		_w7020_,
		_w7389_
	);
	LUT4 #(
		.INIT('h2228)
	) name7356 (
		_w2407_,
		_w3409_,
		_w3650_,
		_w6959_,
		_w7390_
	);
	LUT2 #(
		.INIT('h1)
	) name7357 (
		_w7389_,
		_w7390_,
		_w7391_
	);
	LUT2 #(
		.INIT('h4)
	) name7358 (
		_w7388_,
		_w7391_,
		_w7392_
	);
	LUT2 #(
		.INIT('h4)
	) name7359 (
		_w7387_,
		_w7392_,
		_w7393_
	);
	LUT3 #(
		.INIT('h82)
	) name7360 (
		_w2550_,
		_w7117_,
		_w7119_,
		_w7394_
	);
	LUT3 #(
		.INIT('h82)
	) name7361 (
		_w2854_,
		_w6967_,
		_w6969_,
		_w7395_
	);
	LUT2 #(
		.INIT('h8)
	) name7362 (
		_w2549_,
		_w7014_,
		_w7396_
	);
	LUT4 #(
		.INIT('h02a8)
	) name7363 (
		_w2617_,
		_w3257_,
		_w6964_,
		_w6966_,
		_w7397_
	);
	LUT2 #(
		.INIT('h1)
	) name7364 (
		_w7396_,
		_w7397_,
		_w7398_
	);
	LUT2 #(
		.INIT('h4)
	) name7365 (
		_w7395_,
		_w7398_,
		_w7399_
	);
	LUT3 #(
		.INIT('h9a)
	) name7366 (
		\a[29] ,
		_w7394_,
		_w7399_,
		_w7400_
	);
	LUT3 #(
		.INIT('hd4)
	) name7367 (
		_w7386_,
		_w7393_,
		_w7400_,
		_w7401_
	);
	LUT2 #(
		.INIT('h9)
	) name7368 (
		_w7361_,
		_w7363_,
		_w7402_
	);
	LUT4 #(
		.INIT('h54ab)
	) name7369 (
		_w7012_,
		_w7117_,
		_w7118_,
		_w7120_,
		_w7403_
	);
	LUT4 #(
		.INIT('h02a8)
	) name7370 (
		_w2549_,
		_w3257_,
		_w6964_,
		_w6966_,
		_w7404_
	);
	LUT4 #(
		.INIT('h007d)
	) name7371 (
		_w2617_,
		_w6967_,
		_w6969_,
		_w7404_,
		_w7405_
	);
	LUT3 #(
		.INIT('h70)
	) name7372 (
		_w2854_,
		_w7008_,
		_w7405_,
		_w7406_
	);
	LUT4 #(
		.INIT('h95aa)
	) name7373 (
		\a[29] ,
		_w2550_,
		_w7403_,
		_w7406_,
		_w7407_
	);
	LUT3 #(
		.INIT('hb2)
	) name7374 (
		_w7401_,
		_w7402_,
		_w7407_,
		_w7408_
	);
	LUT4 #(
		.INIT('h02a8)
	) name7375 (
		_w2875_,
		_w7004_,
		_w7127_,
		_w7128_,
		_w7409_
	);
	LUT4 #(
		.INIT('h04c8)
	) name7376 (
		_w2622_,
		_w2986_,
		_w6978_,
		_w6980_,
		_w7410_
	);
	LUT3 #(
		.INIT('h84)
	) name7377 (
		_w2872_,
		_w2874_,
		_w6975_,
		_w7411_
	);
	LUT3 #(
		.INIT('h07)
	) name7378 (
		_w2975_,
		_w7002_,
		_w7411_,
		_w7412_
	);
	LUT2 #(
		.INIT('h4)
	) name7379 (
		_w7410_,
		_w7412_,
		_w7413_
	);
	LUT3 #(
		.INIT('h9a)
	) name7380 (
		\a[26] ,
		_w7409_,
		_w7413_,
		_w7414_
	);
	LUT3 #(
		.INIT('hd4)
	) name7381 (
		_w7385_,
		_w7408_,
		_w7414_,
		_w7415_
	);
	LUT3 #(
		.INIT('h69)
	) name7382 (
		_w7384_,
		_w7415_,
		_w7179_,
		_w7416_
	);
	LUT2 #(
		.INIT('h8)
	) name7383 (
		_w7136_,
		_w7167_,
		_w7417_
	);
	LUT3 #(
		.INIT('h7e)
	) name7384 (
		_w6989_,
		_w7136_,
		_w7165_,
		_w7418_
	);
	LUT4 #(
		.INIT('h8a88)
	) name7385 (
		_w7417_,
		_w7170_,
		_w7135_,
		_w7172_,
		_w7419_
	);
	LUT4 #(
		.INIT('h028a)
	) name7386 (
		_w3311_,
		_w7136_,
		_w7166_,
		_w7167_,
		_w7420_
	);
	LUT4 #(
		.INIT('h781e)
	) name7387 (
		\a[17] ,
		\a[18] ,
		\a[19] ,
		\a[20] ,
		_w7421_
	);
	LUT3 #(
		.INIT('hb0)
	) name7388 (
		_w7136_,
		_w7166_,
		_w7421_,
		_w7422_
	);
	LUT2 #(
		.INIT('h1)
	) name7389 (
		_w7420_,
		_w7422_,
		_w7423_
	);
	LUT4 #(
		.INIT('h5700)
	) name7390 (
		_w3312_,
		_w7418_,
		_w7419_,
		_w7423_,
		_w7424_
	);
	LUT2 #(
		.INIT('h6)
	) name7391 (
		\a[20] ,
		_w7424_,
		_w7425_
	);
	LUT4 #(
		.INIT('h54ab)
	) name7392 (
		_w7006_,
		_w7123_,
		_w7124_,
		_w7126_,
		_w7426_
	);
	LUT4 #(
		.INIT('h02a8)
	) name7393 (
		_w2874_,
		_w2983_,
		_w6972_,
		_w6974_,
		_w7427_
	);
	LUT4 #(
		.INIT('h007b)
	) name7394 (
		_w2872_,
		_w2975_,
		_w6975_,
		_w7427_,
		_w7428_
	);
	LUT3 #(
		.INIT('h70)
	) name7395 (
		_w2986_,
		_w7002_,
		_w7428_,
		_w7429_
	);
	LUT4 #(
		.INIT('h95aa)
	) name7396 (
		\a[26] ,
		_w2875_,
		_w7426_,
		_w7429_,
		_w7430_
	);
	LUT4 #(
		.INIT('h0096)
	) name7397 (
		_w7401_,
		_w7402_,
		_w7407_,
		_w7430_,
		_w7431_
	);
	LUT4 #(
		.INIT('h6900)
	) name7398 (
		_w7401_,
		_w7402_,
		_w7407_,
		_w7430_,
		_w7432_
	);
	LUT4 #(
		.INIT('h9669)
	) name7399 (
		_w7401_,
		_w7402_,
		_w7407_,
		_w7430_,
		_w7433_
	);
	LUT4 #(
		.INIT('h1000)
	) name7400 (
		_w60_,
		_w244_,
		_w830_,
		_w1303_,
		_w7434_
	);
	LUT4 #(
		.INIT('h4000)
	) name7401 (
		_w393_,
		_w403_,
		_w1084_,
		_w2453_,
		_w7435_
	);
	LUT2 #(
		.INIT('h8)
	) name7402 (
		_w7434_,
		_w7435_,
		_w7436_
	);
	LUT4 #(
		.INIT('h153f)
	) name7403 (
		_w85_,
		_w90_,
		_w39_,
		_w166_,
		_w7437_
	);
	LUT3 #(
		.INIT('h80)
	) name7404 (
		_w356_,
		_w497_,
		_w7437_,
		_w7438_
	);
	LUT3 #(
		.INIT('h80)
	) name7405 (
		_w1180_,
		_w1222_,
		_w2582_,
		_w7439_
	);
	LUT4 #(
		.INIT('h0777)
	) name7406 (
		_w106_,
		_w67_,
		_w44_,
		_w184_,
		_w7440_
	);
	LUT4 #(
		.INIT('h8000)
	) name7407 (
		_w597_,
		_w598_,
		_w793_,
		_w7440_,
		_w7441_
	);
	LUT3 #(
		.INIT('h80)
	) name7408 (
		_w7438_,
		_w7439_,
		_w7441_,
		_w7442_
	);
	LUT2 #(
		.INIT('h8)
	) name7409 (
		_w7436_,
		_w7442_,
		_w7443_
	);
	LUT4 #(
		.INIT('h135f)
	) name7410 (
		_w67_,
		_w72_,
		_w43_,
		_w44_,
		_w7444_
	);
	LUT4 #(
		.INIT('h135f)
	) name7411 (
		_w47_,
		_w44_,
		_w166_,
		_w259_,
		_w7445_
	);
	LUT4 #(
		.INIT('h8000)
	) name7412 (
		_w611_,
		_w1003_,
		_w7445_,
		_w7444_,
		_w7446_
	);
	LUT4 #(
		.INIT('h0777)
	) name7413 (
		_w50_,
		_w43_,
		_w93_,
		_w158_,
		_w7447_
	);
	LUT4 #(
		.INIT('h4000)
	) name7414 (
		_w454_,
		_w1575_,
		_w3022_,
		_w7447_,
		_w7448_
	);
	LUT4 #(
		.INIT('h8000)
	) name7415 (
		_w1870_,
		_w2028_,
		_w7446_,
		_w7448_,
		_w7449_
	);
	LUT4 #(
		.INIT('h8000)
	) name7416 (
		_w604_,
		_w1248_,
		_w1754_,
		_w3811_,
		_w7450_
	);
	LUT4 #(
		.INIT('h135f)
	) name7417 (
		_w67_,
		_w47_,
		_w236_,
		_w176_,
		_w7451_
	);
	LUT4 #(
		.INIT('h8000)
	) name7418 (
		_w513_,
		_w2706_,
		_w2803_,
		_w7451_,
		_w7452_
	);
	LUT4 #(
		.INIT('h8000)
	) name7419 (
		_w2660_,
		_w2663_,
		_w7450_,
		_w7452_,
		_w7453_
	);
	LUT4 #(
		.INIT('h8000)
	) name7420 (
		_w1903_,
		_w1914_,
		_w7449_,
		_w7453_,
		_w7454_
	);
	LUT4 #(
		.INIT('h0888)
	) name7421 (
		_w7324_,
		_w7331_,
		_w7443_,
		_w7454_,
		_w7455_
	);
	LUT4 #(
		.INIT('h7000)
	) name7422 (
		_w7324_,
		_w7331_,
		_w7443_,
		_w7454_,
		_w7456_
	);
	LUT4 #(
		.INIT('h8777)
	) name7423 (
		_w7324_,
		_w7331_,
		_w7443_,
		_w7454_,
		_w7457_
	);
	LUT3 #(
		.INIT('h82)
	) name7424 (
		_w377_,
		_w7105_,
		_w7107_,
		_w7458_
	);
	LUT3 #(
		.INIT('h82)
	) name7425 (
		_w2527_,
		_w3706_,
		_w6957_,
		_w7459_
	);
	LUT2 #(
		.INIT('h8)
	) name7426 (
		_w376_,
		_w7026_,
		_w7460_
	);
	LUT4 #(
		.INIT('h02a8)
	) name7427 (
		_w2407_,
		_w3882_,
		_w6954_,
		_w6956_,
		_w7461_
	);
	LUT2 #(
		.INIT('h1)
	) name7428 (
		_w7460_,
		_w7461_,
		_w7462_
	);
	LUT2 #(
		.INIT('h4)
	) name7429 (
		_w7459_,
		_w7462_,
		_w7463_
	);
	LUT4 #(
		.INIT('h4544)
	) name7430 (
		_w7455_,
		_w7456_,
		_w7458_,
		_w7463_,
		_w7464_
	);
	LUT4 #(
		.INIT('h54ab)
	) name7431 (
		_w7024_,
		_w7105_,
		_w7106_,
		_w7108_,
		_w7465_
	);
	LUT4 #(
		.INIT('h02a8)
	) name7432 (
		_w376_,
		_w3882_,
		_w6954_,
		_w6956_,
		_w7466_
	);
	LUT4 #(
		.INIT('h007d)
	) name7433 (
		_w2407_,
		_w3706_,
		_w6957_,
		_w7466_,
		_w7467_
	);
	LUT3 #(
		.INIT('h70)
	) name7434 (
		_w2527_,
		_w7020_,
		_w7467_,
		_w7468_
	);
	LUT3 #(
		.INIT('h70)
	) name7435 (
		_w377_,
		_w7465_,
		_w7468_,
		_w7469_
	);
	LUT4 #(
		.INIT('hf990)
	) name7436 (
		_w7347_,
		_w7349_,
		_w7464_,
		_w7469_,
		_w7470_
	);
	LUT4 #(
		.INIT('h02a8)
	) name7437 (
		_w2550_,
		_w7016_,
		_w7115_,
		_w7116_,
		_w7471_
	);
	LUT4 #(
		.INIT('h02a8)
	) name7438 (
		_w2854_,
		_w3257_,
		_w6964_,
		_w6966_,
		_w7472_
	);
	LUT3 #(
		.INIT('h82)
	) name7439 (
		_w2549_,
		_w6960_,
		_w6962_,
		_w7473_
	);
	LUT3 #(
		.INIT('h07)
	) name7440 (
		_w2617_,
		_w7014_,
		_w7473_,
		_w7474_
	);
	LUT2 #(
		.INIT('h4)
	) name7441 (
		_w7472_,
		_w7474_,
		_w7475_
	);
	LUT3 #(
		.INIT('h9a)
	) name7442 (
		\a[29] ,
		_w7471_,
		_w7475_,
		_w7476_
	);
	LUT4 #(
		.INIT('hf660)
	) name7443 (
		_w7353_,
		_w7359_,
		_w7470_,
		_w7476_,
		_w7477_
	);
	LUT4 #(
		.INIT('h0096)
	) name7444 (
		_w7386_,
		_w7393_,
		_w7400_,
		_w7477_,
		_w7478_
	);
	LUT4 #(
		.INIT('h6900)
	) name7445 (
		_w7386_,
		_w7393_,
		_w7400_,
		_w7477_,
		_w7479_
	);
	LUT3 #(
		.INIT('h82)
	) name7446 (
		_w2875_,
		_w7123_,
		_w7125_,
		_w7480_
	);
	LUT3 #(
		.INIT('h84)
	) name7447 (
		_w2872_,
		_w2986_,
		_w6975_,
		_w7481_
	);
	LUT2 #(
		.INIT('h8)
	) name7448 (
		_w2874_,
		_w7008_,
		_w7482_
	);
	LUT4 #(
		.INIT('h02a8)
	) name7449 (
		_w2975_,
		_w2983_,
		_w6972_,
		_w6974_,
		_w7483_
	);
	LUT2 #(
		.INIT('h1)
	) name7450 (
		_w7482_,
		_w7483_,
		_w7484_
	);
	LUT2 #(
		.INIT('h4)
	) name7451 (
		_w7481_,
		_w7484_,
		_w7485_
	);
	LUT3 #(
		.INIT('h9a)
	) name7452 (
		\a[26] ,
		_w7480_,
		_w7485_,
		_w7486_
	);
	LUT3 #(
		.INIT('h54)
	) name7453 (
		_w7478_,
		_w7479_,
		_w7486_,
		_w7487_
	);
	LUT3 #(
		.INIT('h54)
	) name7454 (
		_w7431_,
		_w7432_,
		_w7487_,
		_w7488_
	);
	LUT3 #(
		.INIT('h69)
	) name7455 (
		_w7385_,
		_w7408_,
		_w7414_,
		_w7489_
	);
	LUT4 #(
		.INIT('h02a8)
	) name7456 (
		_w37_,
		_w6998_,
		_w7133_,
		_w7134_,
		_w7490_
	);
	LUT4 #(
		.INIT('h04c8)
	) name7457 (
		_w2411_,
		_w3262_,
		_w6983_,
		_w6993_,
		_w7491_
	);
	LUT3 #(
		.INIT('h82)
	) name7458 (
		_w3214_,
		_w2546_,
		_w6981_,
		_w7492_
	);
	LUT3 #(
		.INIT('h07)
	) name7459 (
		_w3249_,
		_w6996_,
		_w7492_,
		_w7493_
	);
	LUT2 #(
		.INIT('h4)
	) name7460 (
		_w7491_,
		_w7493_,
		_w7494_
	);
	LUT3 #(
		.INIT('h9a)
	) name7461 (
		\a[23] ,
		_w7490_,
		_w7494_,
		_w7495_
	);
	LUT4 #(
		.INIT('h0115)
	) name7462 (
		_w7425_,
		_w7488_,
		_w7489_,
		_w7495_,
		_w7496_
	);
	LUT4 #(
		.INIT('ha880)
	) name7463 (
		_w7425_,
		_w7488_,
		_w7489_,
		_w7495_,
		_w7497_
	);
	LUT4 #(
		.INIT('h566a)
	) name7464 (
		_w7425_,
		_w7488_,
		_w7489_,
		_w7495_,
		_w7498_
	);
	LUT2 #(
		.INIT('h9)
	) name7465 (
		_w7416_,
		_w7498_,
		_w7499_
	);
	LUT4 #(
		.INIT('h54ab)
	) name7466 (
		_w7000_,
		_w7129_,
		_w7130_,
		_w7132_,
		_w7500_
	);
	LUT4 #(
		.INIT('h02a8)
	) name7467 (
		_w3214_,
		_w2622_,
		_w6978_,
		_w6980_,
		_w7501_
	);
	LUT4 #(
		.INIT('h007b)
	) name7468 (
		_w2546_,
		_w3249_,
		_w6981_,
		_w7501_,
		_w7502_
	);
	LUT3 #(
		.INIT('h70)
	) name7469 (
		_w3262_,
		_w6996_,
		_w7502_,
		_w7503_
	);
	LUT4 #(
		.INIT('h95aa)
	) name7470 (
		\a[23] ,
		_w37_,
		_w7500_,
		_w7503_,
		_w7504_
	);
	LUT3 #(
		.INIT('h09)
	) name7471 (
		_w7433_,
		_w7487_,
		_w7504_,
		_w7505_
	);
	LUT3 #(
		.INIT('h96)
	) name7472 (
		_w7433_,
		_w7487_,
		_w7504_,
		_w7506_
	);
	LUT4 #(
		.INIT('h9669)
	) name7473 (
		_w7386_,
		_w7393_,
		_w7400_,
		_w7477_,
		_w7507_
	);
	LUT2 #(
		.INIT('h9)
	) name7474 (
		_w7486_,
		_w7507_,
		_w7508_
	);
	LUT4 #(
		.INIT('h2228)
	) name7475 (
		_w2549_,
		_w3409_,
		_w3650_,
		_w6959_,
		_w7509_
	);
	LUT4 #(
		.INIT('h007d)
	) name7476 (
		_w2617_,
		_w6960_,
		_w6962_,
		_w7509_,
		_w7510_
	);
	LUT3 #(
		.INIT('h70)
	) name7477 (
		_w2854_,
		_w7014_,
		_w7510_,
		_w7511_
	);
	LUT4 #(
		.INIT('h95aa)
	) name7478 (
		\a[29] ,
		_w2550_,
		_w7291_,
		_w7511_,
		_w7512_
	);
	LUT4 #(
		.INIT('h6996)
	) name7479 (
		_w7347_,
		_w7349_,
		_w7464_,
		_w7469_,
		_w7513_
	);
	LUT2 #(
		.INIT('h4)
	) name7480 (
		_w7512_,
		_w7513_,
		_w7514_
	);
	LUT4 #(
		.INIT('h0777)
	) name7481 (
		_w85_,
		_w43_,
		_w44_,
		_w184_,
		_w7515_
	);
	LUT4 #(
		.INIT('h0777)
	) name7482 (
		_w43_,
		_w65_,
		_w46_,
		_w378_,
		_w7516_
	);
	LUT4 #(
		.INIT('h4000)
	) name7483 (
		_w363_,
		_w1074_,
		_w7516_,
		_w7515_,
		_w7517_
	);
	LUT4 #(
		.INIT('h135f)
	) name7484 (
		_w56_,
		_w47_,
		_w39_,
		_w43_,
		_w7518_
	);
	LUT4 #(
		.INIT('h8000)
	) name7485 (
		_w292_,
		_w287_,
		_w3109_,
		_w7518_,
		_w7519_
	);
	LUT3 #(
		.INIT('h80)
	) name7486 (
		_w3034_,
		_w7517_,
		_w7519_,
		_w7520_
	);
	LUT3 #(
		.INIT('h37)
	) name7487 (
		_w122_,
		_w65_,
		_w166_,
		_w7521_
	);
	LUT4 #(
		.INIT('h8000)
	) name7488 (
		_w657_,
		_w1628_,
		_w2274_,
		_w7521_,
		_w7522_
	);
	LUT3 #(
		.INIT('h1f)
	) name7489 (
		_w56_,
		_w93_,
		_w158_,
		_w7523_
	);
	LUT4 #(
		.INIT('h153f)
	) name7490 (
		_w110_,
		_w65_,
		_w378_,
		_w430_,
		_w7524_
	);
	LUT4 #(
		.INIT('h8000)
	) name7491 (
		_w777_,
		_w1410_,
		_w7523_,
		_w7524_,
		_w7525_
	);
	LUT4 #(
		.INIT('h153f)
	) name7492 (
		_w56_,
		_w41_,
		_w39_,
		_w236_,
		_w7526_
	);
	LUT4 #(
		.INIT('h153f)
	) name7493 (
		_w85_,
		_w41_,
		_w176_,
		_w378_,
		_w7527_
	);
	LUT4 #(
		.INIT('h4000)
	) name7494 (
		_w432_,
		_w1847_,
		_w7526_,
		_w7527_,
		_w7528_
	);
	LUT4 #(
		.INIT('h4000)
	) name7495 (
		_w452_,
		_w793_,
		_w902_,
		_w2372_,
		_w7529_
	);
	LUT4 #(
		.INIT('h8000)
	) name7496 (
		_w7522_,
		_w7525_,
		_w7528_,
		_w7529_,
		_w7530_
	);
	LUT4 #(
		.INIT('h8000)
	) name7497 (
		_w2233_,
		_w2245_,
		_w7520_,
		_w7530_,
		_w7531_
	);
	LUT2 #(
		.INIT('h8)
	) name7498 (
		_w3951_,
		_w7531_,
		_w7532_
	);
	LUT3 #(
		.INIT('h80)
	) name7499 (
		_w982_,
		_w1307_,
		_w3804_,
		_w7533_
	);
	LUT3 #(
		.INIT('h40)
	) name7500 (
		_w94_,
		_w1993_,
		_w2136_,
		_w7534_
	);
	LUT2 #(
		.INIT('h8)
	) name7501 (
		_w1363_,
		_w7534_,
		_w7535_
	);
	LUT4 #(
		.INIT('h4000)
	) name7502 (
		_w355_,
		_w824_,
		_w825_,
		_w2008_,
		_w7536_
	);
	LUT4 #(
		.INIT('h135f)
	) name7503 (
		_w65_,
		_w44_,
		_w184_,
		_w158_,
		_w7537_
	);
	LUT3 #(
		.INIT('h80)
	) name7504 (
		_w1668_,
		_w2137_,
		_w7537_,
		_w7538_
	);
	LUT4 #(
		.INIT('h0777)
	) name7505 (
		_w59_,
		_w78_,
		_w50_,
		_w419_,
		_w7539_
	);
	LUT4 #(
		.INIT('h4000)
	) name7506 (
		_w337_,
		_w560_,
		_w1333_,
		_w7539_,
		_w7540_
	);
	LUT4 #(
		.INIT('h8000)
	) name7507 (
		_w3110_,
		_w7538_,
		_w7540_,
		_w7536_,
		_w7541_
	);
	LUT4 #(
		.INIT('h8000)
	) name7508 (
		_w633_,
		_w647_,
		_w7535_,
		_w7541_,
		_w7542_
	);
	LUT2 #(
		.INIT('h8)
	) name7509 (
		_w7533_,
		_w7542_,
		_w7543_
	);
	LUT4 #(
		.INIT('h0777)
	) name7510 (
		_w3951_,
		_w7531_,
		_w7533_,
		_w7542_,
		_w7544_
	);
	LUT4 #(
		.INIT('h8001)
	) name7511 (
		\a[8] ,
		\a[9] ,
		\a[10] ,
		\a[11] ,
		_w7545_
	);
	LUT4 #(
		.INIT('h559a)
	) name7512 (
		\a[11] ,
		_w7136_,
		_w7166_,
		_w7545_,
		_w7546_
	);
	LUT4 #(
		.INIT('h8000)
	) name7513 (
		_w3951_,
		_w7531_,
		_w7533_,
		_w7542_,
		_w7547_
	);
	LUT4 #(
		.INIT('h7888)
	) name7514 (
		_w3951_,
		_w7531_,
		_w7533_,
		_w7542_,
		_w7548_
	);
	LUT3 #(
		.INIT('h51)
	) name7515 (
		_w7544_,
		_w7546_,
		_w7547_,
		_w7549_
	);
	LUT4 #(
		.INIT('h2a02)
	) name7516 (
		_w7332_,
		_w7532_,
		_w7543_,
		_w7546_,
		_w7550_
	);
	LUT4 #(
		.INIT('h4054)
	) name7517 (
		_w7332_,
		_w7532_,
		_w7543_,
		_w7546_,
		_w7551_
	);
	LUT4 #(
		.INIT('h6656)
	) name7518 (
		_w7332_,
		_w7544_,
		_w7546_,
		_w7547_,
		_w7552_
	);
	LUT4 #(
		.INIT('h02a8)
	) name7519 (
		_w377_,
		_w7028_,
		_w7103_,
		_w7104_,
		_w7553_
	);
	LUT4 #(
		.INIT('h02a8)
	) name7520 (
		_w2527_,
		_w3882_,
		_w6954_,
		_w6956_,
		_w7554_
	);
	LUT3 #(
		.INIT('h82)
	) name7521 (
		_w376_,
		_w4030_,
		_w6952_,
		_w7555_
	);
	LUT3 #(
		.INIT('h07)
	) name7522 (
		_w2407_,
		_w7026_,
		_w7555_,
		_w7556_
	);
	LUT2 #(
		.INIT('h4)
	) name7523 (
		_w7554_,
		_w7556_,
		_w7557_
	);
	LUT2 #(
		.INIT('h4)
	) name7524 (
		_w7553_,
		_w7557_,
		_w7558_
	);
	LUT3 #(
		.INIT('h65)
	) name7525 (
		_w7457_,
		_w7458_,
		_w7463_,
		_w7559_
	);
	LUT4 #(
		.INIT('h2b00)
	) name7526 (
		_w7332_,
		_w7549_,
		_w7558_,
		_w7559_,
		_w7560_
	);
	LUT4 #(
		.INIT('h54ab)
	) name7527 (
		_w7550_,
		_w7551_,
		_w7558_,
		_w7559_,
		_w7561_
	);
	LUT4 #(
		.INIT('h54ab)
	) name7528 (
		_w7030_,
		_w7099_,
		_w7100_,
		_w7102_,
		_w7562_
	);
	LUT4 #(
		.INIT('h2228)
	) name7529 (
		_w376_,
		_w4099_,
		_w4378_,
		_w6951_,
		_w7563_
	);
	LUT4 #(
		.INIT('h007d)
	) name7530 (
		_w2407_,
		_w4030_,
		_w6952_,
		_w7563_,
		_w7564_
	);
	LUT3 #(
		.INIT('h70)
	) name7531 (
		_w2527_,
		_w7026_,
		_w7564_,
		_w7565_
	);
	LUT3 #(
		.INIT('h70)
	) name7532 (
		_w377_,
		_w7562_,
		_w7565_,
		_w7566_
	);
	LUT3 #(
		.INIT('h06)
	) name7533 (
		_w7546_,
		_w7548_,
		_w7566_,
		_w7567_
	);
	LUT4 #(
		.INIT('h135f)
	) name7534 (
		_w38_,
		_w67_,
		_w78_,
		_w166_,
		_w7568_
	);
	LUT3 #(
		.INIT('h40)
	) name7535 (
		_w362_,
		_w1014_,
		_w7568_,
		_w7569_
	);
	LUT3 #(
		.INIT('h80)
	) name7536 (
		_w2208_,
		_w3160_,
		_w7569_,
		_w7570_
	);
	LUT4 #(
		.INIT('h0777)
	) name7537 (
		_w78_,
		_w56_,
		_w47_,
		_w72_,
		_w7571_
	);
	LUT4 #(
		.INIT('h0777)
	) name7538 (
		_w106_,
		_w90_,
		_w44_,
		_w166_,
		_w7572_
	);
	LUT2 #(
		.INIT('h8)
	) name7539 (
		_w7571_,
		_w7572_,
		_w7573_
	);
	LUT4 #(
		.INIT('h135f)
	) name7540 (
		_w90_,
		_w46_,
		_w236_,
		_w378_,
		_w7574_
	);
	LUT3 #(
		.INIT('h37)
	) name7541 (
		_w55_,
		_w72_,
		_w93_,
		_w7575_
	);
	LUT4 #(
		.INIT('h4000)
	) name7542 (
		_w450_,
		_w739_,
		_w7575_,
		_w7574_,
		_w7576_
	);
	LUT4 #(
		.INIT('h8000)
	) name7543 (
		_w777_,
		_w1470_,
		_w1481_,
		_w1514_,
		_w7577_
	);
	LUT4 #(
		.INIT('h8000)
	) name7544 (
		_w756_,
		_w7573_,
		_w7577_,
		_w7576_,
		_w7578_
	);
	LUT3 #(
		.INIT('h80)
	) name7545 (
		_w1805_,
		_w7570_,
		_w7578_,
		_w7579_
	);
	LUT3 #(
		.INIT('h80)
	) name7546 (
		_w3444_,
		_w3469_,
		_w7211_,
		_w7580_
	);
	LUT4 #(
		.INIT('h2000)
	) name7547 (
		_w148_,
		_w325_,
		_w495_,
		_w1931_,
		_w7581_
	);
	LUT2 #(
		.INIT('h8)
	) name7548 (
		_w7580_,
		_w7581_,
		_w7582_
	);
	LUT4 #(
		.INIT('h8000)
	) name7549 (
		_w219_,
		_w196_,
		_w681_,
		_w2661_,
		_w7583_
	);
	LUT4 #(
		.INIT('h0777)
	) name7550 (
		_w56_,
		_w72_,
		_w43_,
		_w44_,
		_w7584_
	);
	LUT4 #(
		.INIT('h153f)
	) name7551 (
		_w47_,
		_w46_,
		_w184_,
		_w378_,
		_w7585_
	);
	LUT4 #(
		.INIT('h8000)
	) name7552 (
		_w496_,
		_w750_,
		_w7584_,
		_w7585_,
		_w7586_
	);
	LUT4 #(
		.INIT('h8000)
	) name7553 (
		_w403_,
		_w829_,
		_w1084_,
		_w1658_,
		_w7587_
	);
	LUT3 #(
		.INIT('h80)
	) name7554 (
		_w7583_,
		_w7586_,
		_w7587_,
		_w7588_
	);
	LUT3 #(
		.INIT('h80)
	) name7555 (
		_w3090_,
		_w7582_,
		_w7588_,
		_w7589_
	);
	LUT2 #(
		.INIT('h8)
	) name7556 (
		_w7579_,
		_w7589_,
		_w7590_
	);
	LUT4 #(
		.INIT('h135f)
	) name7557 (
		_w52_,
		_w90_,
		_w166_,
		_w378_,
		_w7591_
	);
	LUT4 #(
		.INIT('h135f)
	) name7558 (
		_w67_,
		_w72_,
		_w43_,
		_w93_,
		_w7592_
	);
	LUT4 #(
		.INIT('h4000)
	) name7559 (
		_w468_,
		_w1871_,
		_w7592_,
		_w7591_,
		_w7593_
	);
	LUT3 #(
		.INIT('h80)
	) name7560 (
		_w898_,
		_w2783_,
		_w7593_,
		_w7594_
	);
	LUT3 #(
		.INIT('h80)
	) name7561 (
		_w311_,
		_w803_,
		_w1549_,
		_w7595_
	);
	LUT4 #(
		.INIT('h153f)
	) name7562 (
		_w55_,
		_w78_,
		_w93_,
		_w201_,
		_w7596_
	);
	LUT4 #(
		.INIT('h135f)
	) name7563 (
		_w50_,
		_w65_,
		_w201_,
		_w166_,
		_w7597_
	);
	LUT4 #(
		.INIT('h2000)
	) name7564 (
		_w370_,
		_w412_,
		_w7596_,
		_w7597_,
		_w7598_
	);
	LUT4 #(
		.INIT('h1000)
	) name7565 (
		_w358_,
		_w429_,
		_w798_,
		_w2086_,
		_w7599_
	);
	LUT4 #(
		.INIT('h0200)
	) name7566 (
		_w81_,
		_w402_,
		_w379_,
		_w512_,
		_w7600_
	);
	LUT4 #(
		.INIT('h8000)
	) name7567 (
		_w7595_,
		_w7598_,
		_w7599_,
		_w7600_,
		_w7601_
	);
	LUT3 #(
		.INIT('h80)
	) name7568 (
		_w446_,
		_w1342_,
		_w1752_,
		_w7602_
	);
	LUT4 #(
		.INIT('h153f)
	) name7569 (
		_w38_,
		_w78_,
		_w90_,
		_w39_,
		_w7603_
	);
	LUT3 #(
		.INIT('h1f)
	) name7570 (
		_w67_,
		_w47_,
		_w166_,
		_w7604_
	);
	LUT4 #(
		.INIT('h8000)
	) name7571 (
		_w312_,
		_w944_,
		_w7603_,
		_w7604_,
		_w7605_
	);
	LUT3 #(
		.INIT('h80)
	) name7572 (
		_w7233_,
		_w7602_,
		_w7605_,
		_w7606_
	);
	LUT3 #(
		.INIT('h80)
	) name7573 (
		_w1003_,
		_w1045_,
		_w1978_,
		_w7607_
	);
	LUT4 #(
		.INIT('h153f)
	) name7574 (
		_w90_,
		_w41_,
		_w184_,
		_w176_,
		_w7608_
	);
	LUT4 #(
		.INIT('h153f)
	) name7575 (
		_w90_,
		_w43_,
		_w44_,
		_w201_,
		_w7609_
	);
	LUT4 #(
		.INIT('h4000)
	) name7576 (
		_w439_,
		_w978_,
		_w7609_,
		_w7608_,
		_w7610_
	);
	LUT4 #(
		.INIT('h4000)
	) name7577 (
		_w104_,
		_w643_,
		_w1450_,
		_w3029_,
		_w7611_
	);
	LUT3 #(
		.INIT('h80)
	) name7578 (
		_w7607_,
		_w7610_,
		_w7611_,
		_w7612_
	);
	LUT4 #(
		.INIT('h8000)
	) name7579 (
		_w7606_,
		_w7612_,
		_w7594_,
		_w7601_,
		_w7613_
	);
	LUT2 #(
		.INIT('h8)
	) name7580 (
		_w2036_,
		_w7613_,
		_w7614_
	);
	LUT4 #(
		.INIT('h153f)
	) name7581 (
		_w59_,
		_w47_,
		_w43_,
		_w259_,
		_w7615_
	);
	LUT4 #(
		.INIT('h8000)
	) name7582 (
		_w678_,
		_w1628_,
		_w1647_,
		_w7615_,
		_w7616_
	);
	LUT3 #(
		.INIT('h80)
	) name7583 (
		_w1675_,
		_w1860_,
		_w7616_,
		_w7617_
	);
	LUT4 #(
		.INIT('h153f)
	) name7584 (
		_w52_,
		_w44_,
		_w158_,
		_w176_,
		_w7618_
	);
	LUT3 #(
		.INIT('h1f)
	) name7585 (
		_w56_,
		_w44_,
		_w430_,
		_w7619_
	);
	LUT4 #(
		.INIT('h8000)
	) name7586 (
		_w621_,
		_w783_,
		_w7618_,
		_w7619_,
		_w7620_
	);
	LUT4 #(
		.INIT('h1000)
	) name7587 (
		_w190_,
		_w310_,
		_w1097_,
		_w3432_,
		_w7621_
	);
	LUT2 #(
		.INIT('h8)
	) name7588 (
		_w7620_,
		_w7621_,
		_w7622_
	);
	LUT2 #(
		.INIT('h4)
	) name7589 (
		_w206_,
		_w4265_,
		_w7623_
	);
	LUT4 #(
		.INIT('h153f)
	) name7590 (
		_w55_,
		_w50_,
		_w43_,
		_w378_,
		_w7624_
	);
	LUT4 #(
		.INIT('h135f)
	) name7591 (
		_w110_,
		_w90_,
		_w184_,
		_w236_,
		_w7625_
	);
	LUT4 #(
		.INIT('h4000)
	) name7592 (
		_w206_,
		_w4265_,
		_w7624_,
		_w7625_,
		_w7626_
	);
	LUT3 #(
		.INIT('h80)
	) name7593 (
		_w937_,
		_w1682_,
		_w2764_,
		_w7627_
	);
	LUT3 #(
		.INIT('h80)
	) name7594 (
		_w1775_,
		_w7626_,
		_w7627_,
		_w7628_
	);
	LUT3 #(
		.INIT('h80)
	) name7595 (
		_w7617_,
		_w7622_,
		_w7628_,
		_w7629_
	);
	LUT4 #(
		.INIT('h8000)
	) name7596 (
		_w1336_,
		_w1349_,
		_w2488_,
		_w2498_,
		_w7630_
	);
	LUT2 #(
		.INIT('h8)
	) name7597 (
		_w7629_,
		_w7630_,
		_w7631_
	);
	LUT4 #(
		.INIT('h0777)
	) name7598 (
		_w2036_,
		_w7613_,
		_w7629_,
		_w7630_,
		_w7632_
	);
	LUT4 #(
		.INIT('h8001)
	) name7599 (
		\a[5] ,
		\a[6] ,
		\a[7] ,
		\a[8] ,
		_w7633_
	);
	LUT4 #(
		.INIT('h559a)
	) name7600 (
		\a[8] ,
		_w7136_,
		_w7166_,
		_w7633_,
		_w7634_
	);
	LUT4 #(
		.INIT('h8000)
	) name7601 (
		_w2036_,
		_w7613_,
		_w7629_,
		_w7630_,
		_w7635_
	);
	LUT4 #(
		.INIT('h7888)
	) name7602 (
		_w2036_,
		_w7613_,
		_w7629_,
		_w7630_,
		_w7636_
	);
	LUT3 #(
		.INIT('h51)
	) name7603 (
		_w7632_,
		_w7634_,
		_w7635_,
		_w7637_
	);
	LUT4 #(
		.INIT('h2a02)
	) name7604 (
		_w7532_,
		_w7614_,
		_w7631_,
		_w7634_,
		_w7638_
	);
	LUT4 #(
		.INIT('h4054)
	) name7605 (
		_w7532_,
		_w7614_,
		_w7631_,
		_w7634_,
		_w7639_
	);
	LUT4 #(
		.INIT('h6656)
	) name7606 (
		_w7532_,
		_w7632_,
		_w7634_,
		_w7635_,
		_w7640_
	);
	LUT4 #(
		.INIT('h02a8)
	) name7607 (
		_w377_,
		_w7034_,
		_w7097_,
		_w7098_,
		_w7641_
	);
	LUT4 #(
		.INIT('h2228)
	) name7608 (
		_w2527_,
		_w4099_,
		_w4378_,
		_w6951_,
		_w7642_
	);
	LUT3 #(
		.INIT('h82)
	) name7609 (
		_w376_,
		_w6947_,
		_w6949_,
		_w7643_
	);
	LUT3 #(
		.INIT('h07)
	) name7610 (
		_w2407_,
		_w7032_,
		_w7643_,
		_w7644_
	);
	LUT2 #(
		.INIT('h4)
	) name7611 (
		_w7642_,
		_w7644_,
		_w7645_
	);
	LUT2 #(
		.INIT('h4)
	) name7612 (
		_w7641_,
		_w7645_,
		_w7646_
	);
	LUT4 #(
		.INIT('h8777)
	) name7613 (
		_w3951_,
		_w7531_,
		_w7579_,
		_w7589_,
		_w7647_
	);
	LUT4 #(
		.INIT('hd554)
	) name7614 (
		_w7532_,
		_w7590_,
		_w7637_,
		_w7646_,
		_w7648_
	);
	LUT3 #(
		.INIT('h90)
	) name7615 (
		_w7546_,
		_w7548_,
		_w7566_,
		_w7649_
	);
	LUT3 #(
		.INIT('h69)
	) name7616 (
		_w7546_,
		_w7548_,
		_w7566_,
		_w7650_
	);
	LUT3 #(
		.INIT('h54)
	) name7617 (
		_w7567_,
		_w7648_,
		_w7649_,
		_w7651_
	);
	LUT2 #(
		.INIT('h9)
	) name7618 (
		_w7552_,
		_w7558_,
		_w7652_
	);
	LUT4 #(
		.INIT('hba00)
	) name7619 (
		_w7567_,
		_w7648_,
		_w7650_,
		_w7652_,
		_w7653_
	);
	LUT4 #(
		.INIT('h0045)
	) name7620 (
		_w7567_,
		_w7648_,
		_w7650_,
		_w7652_,
		_w7654_
	);
	LUT4 #(
		.INIT('h54ab)
	) name7621 (
		_w7567_,
		_w7648_,
		_w7649_,
		_w7652_,
		_w7655_
	);
	LUT4 #(
		.INIT('h02a8)
	) name7622 (
		_w2550_,
		_w7022_,
		_w7109_,
		_w7110_,
		_w7656_
	);
	LUT4 #(
		.INIT('h2228)
	) name7623 (
		_w2854_,
		_w3409_,
		_w3650_,
		_w6959_,
		_w7657_
	);
	LUT3 #(
		.INIT('h82)
	) name7624 (
		_w2549_,
		_w3706_,
		_w6957_,
		_w7658_
	);
	LUT3 #(
		.INIT('h07)
	) name7625 (
		_w2617_,
		_w7020_,
		_w7658_,
		_w7659_
	);
	LUT2 #(
		.INIT('h4)
	) name7626 (
		_w7657_,
		_w7659_,
		_w7660_
	);
	LUT3 #(
		.INIT('h9a)
	) name7627 (
		\a[29] ,
		_w7656_,
		_w7660_,
		_w7661_
	);
	LUT4 #(
		.INIT('h20a2)
	) name7628 (
		_w7561_,
		_w7651_,
		_w7652_,
		_w7661_,
		_w7662_
	);
	LUT2 #(
		.INIT('h2)
	) name7629 (
		_w7512_,
		_w7513_,
		_w7663_
	);
	LUT2 #(
		.INIT('h9)
	) name7630 (
		_w7512_,
		_w7513_,
		_w7664_
	);
	LUT4 #(
		.INIT('h5501)
	) name7631 (
		_w7514_,
		_w7560_,
		_w7662_,
		_w7663_,
		_w7665_
	);
	LUT4 #(
		.INIT('h9669)
	) name7632 (
		_w7353_,
		_w7359_,
		_w7470_,
		_w7476_,
		_w7666_
	);
	LUT4 #(
		.INIT('h02a8)
	) name7633 (
		_w2875_,
		_w7010_,
		_w7121_,
		_w7122_,
		_w7667_
	);
	LUT4 #(
		.INIT('h04c8)
	) name7634 (
		_w2983_,
		_w2986_,
		_w6972_,
		_w6974_,
		_w7668_
	);
	LUT3 #(
		.INIT('h82)
	) name7635 (
		_w2874_,
		_w6967_,
		_w6969_,
		_w7669_
	);
	LUT3 #(
		.INIT('h07)
	) name7636 (
		_w2975_,
		_w7008_,
		_w7669_,
		_w7670_
	);
	LUT2 #(
		.INIT('h4)
	) name7637 (
		_w7668_,
		_w7670_,
		_w7671_
	);
	LUT3 #(
		.INIT('h9a)
	) name7638 (
		\a[26] ,
		_w7667_,
		_w7671_,
		_w7672_
	);
	LUT3 #(
		.INIT('hb2)
	) name7639 (
		_w7665_,
		_w7666_,
		_w7672_,
		_w7673_
	);
	LUT4 #(
		.INIT('h20a2)
	) name7640 (
		_w7508_,
		_w7665_,
		_w7666_,
		_w7672_,
		_w7674_
	);
	LUT4 #(
		.INIT('h4504)
	) name7641 (
		_w7508_,
		_w7665_,
		_w7666_,
		_w7672_,
		_w7675_
	);
	LUT3 #(
		.INIT('h82)
	) name7642 (
		_w37_,
		_w7129_,
		_w7131_,
		_w7676_
	);
	LUT3 #(
		.INIT('h84)
	) name7643 (
		_w2546_,
		_w3262_,
		_w6981_,
		_w7677_
	);
	LUT2 #(
		.INIT('h8)
	) name7644 (
		_w3214_,
		_w7002_,
		_w7678_
	);
	LUT4 #(
		.INIT('h04c8)
	) name7645 (
		_w2622_,
		_w3249_,
		_w6978_,
		_w6980_,
		_w7679_
	);
	LUT2 #(
		.INIT('h1)
	) name7646 (
		_w7678_,
		_w7679_,
		_w7680_
	);
	LUT2 #(
		.INIT('h4)
	) name7647 (
		_w7677_,
		_w7680_,
		_w7681_
	);
	LUT3 #(
		.INIT('h9a)
	) name7648 (
		\a[23] ,
		_w7676_,
		_w7681_,
		_w7682_
	);
	LUT4 #(
		.INIT('h088a)
	) name7649 (
		_w7506_,
		_w7508_,
		_w7673_,
		_w7682_,
		_w7683_
	);
	LUT3 #(
		.INIT('h69)
	) name7650 (
		_w7488_,
		_w7489_,
		_w7495_,
		_w7684_
	);
	LUT3 #(
		.INIT('h32)
	) name7651 (
		_w7136_,
		_w7166_,
		_w7167_,
		_w7685_
	);
	LUT4 #(
		.INIT('hba00)
	) name7652 (
		_w7170_,
		_w7135_,
		_w7172_,
		_w7685_,
		_w7686_
	);
	LUT4 #(
		.INIT('h0a02)
	) name7653 (
		_w3312_,
		_w7169_,
		_w7419_,
		_w7686_,
		_w7687_
	);
	LUT3 #(
		.INIT('h28)
	) name7654 (
		_w3311_,
		_w7136_,
		_w7168_,
		_w7688_
	);
	LUT3 #(
		.INIT('h40)
	) name7655 (
		_w3654_,
		_w7136_,
		_w7167_,
		_w7689_
	);
	LUT3 #(
		.INIT('h31)
	) name7656 (
		_w7422_,
		_w7688_,
		_w7689_,
		_w7690_
	);
	LUT3 #(
		.INIT('h9a)
	) name7657 (
		\a[20] ,
		_w7687_,
		_w7690_,
		_w7691_
	);
	LUT4 #(
		.INIT('h1f01)
	) name7658 (
		_w7505_,
		_w7683_,
		_w7684_,
		_w7691_,
		_w7692_
	);
	LUT2 #(
		.INIT('h2)
	) name7659 (
		_w7499_,
		_w7692_,
		_w7693_
	);
	LUT2 #(
		.INIT('h4)
	) name7660 (
		_w7499_,
		_w7692_,
		_w7694_
	);
	LUT2 #(
		.INIT('h9)
	) name7661 (
		_w7499_,
		_w7692_,
		_w7695_
	);
	LUT4 #(
		.INIT('h54ab)
	) name7662 (
		_w7170_,
		_w7135_,
		_w7171_,
		_w7685_,
		_w7696_
	);
	LUT3 #(
		.INIT('h28)
	) name7663 (
		_w3645_,
		_w7136_,
		_w7168_,
		_w7697_
	);
	LUT4 #(
		.INIT('h028a)
	) name7664 (
		_w3654_,
		_w7136_,
		_w7166_,
		_w7167_,
		_w7698_
	);
	LUT4 #(
		.INIT('h04c8)
	) name7665 (
		_w2411_,
		_w3311_,
		_w6983_,
		_w6993_,
		_w7699_
	);
	LUT3 #(
		.INIT('h01)
	) name7666 (
		_w7698_,
		_w7699_,
		_w7697_,
		_w7700_
	);
	LUT4 #(
		.INIT('h95aa)
	) name7667 (
		\a[20] ,
		_w3312_,
		_w7696_,
		_w7700_,
		_w7701_
	);
	LUT4 #(
		.INIT('h9a59)
	) name7668 (
		_w7508_,
		_w7665_,
		_w7666_,
		_w7672_,
		_w7702_
	);
	LUT2 #(
		.INIT('h9)
	) name7669 (
		_w7682_,
		_w7702_,
		_w7703_
	);
	LUT4 #(
		.INIT('h02a8)
	) name7670 (
		_w2874_,
		_w3257_,
		_w6964_,
		_w6966_,
		_w7704_
	);
	LUT4 #(
		.INIT('h007d)
	) name7671 (
		_w2975_,
		_w6967_,
		_w6969_,
		_w7704_,
		_w7705_
	);
	LUT3 #(
		.INIT('h70)
	) name7672 (
		_w2986_,
		_w7008_,
		_w7705_,
		_w7706_
	);
	LUT4 #(
		.INIT('h95aa)
	) name7673 (
		\a[26] ,
		_w2875_,
		_w7403_,
		_w7706_,
		_w7707_
	);
	LUT4 #(
		.INIT('h001e)
	) name7674 (
		_w7560_,
		_w7662_,
		_w7664_,
		_w7707_,
		_w7708_
	);
	LUT4 #(
		.INIT('h6665)
	) name7675 (
		_w7561_,
		_w7653_,
		_w7654_,
		_w7661_,
		_w7709_
	);
	LUT3 #(
		.INIT('h82)
	) name7676 (
		_w2550_,
		_w7111_,
		_w7113_,
		_w7710_
	);
	LUT3 #(
		.INIT('h82)
	) name7677 (
		_w2854_,
		_w6960_,
		_w6962_,
		_w7711_
	);
	LUT2 #(
		.INIT('h8)
	) name7678 (
		_w2549_,
		_w7020_,
		_w7712_
	);
	LUT4 #(
		.INIT('h2228)
	) name7679 (
		_w2617_,
		_w3409_,
		_w3650_,
		_w6959_,
		_w7713_
	);
	LUT2 #(
		.INIT('h1)
	) name7680 (
		_w7712_,
		_w7713_,
		_w7714_
	);
	LUT2 #(
		.INIT('h4)
	) name7681 (
		_w7711_,
		_w7714_,
		_w7715_
	);
	LUT3 #(
		.INIT('h9a)
	) name7682 (
		\a[29] ,
		_w7710_,
		_w7715_,
		_w7716_
	);
	LUT3 #(
		.INIT('h82)
	) name7683 (
		_w2875_,
		_w7117_,
		_w7119_,
		_w7717_
	);
	LUT3 #(
		.INIT('h82)
	) name7684 (
		_w2986_,
		_w6967_,
		_w6969_,
		_w7718_
	);
	LUT2 #(
		.INIT('h8)
	) name7685 (
		_w2874_,
		_w7014_,
		_w7719_
	);
	LUT4 #(
		.INIT('h02a8)
	) name7686 (
		_w2975_,
		_w3257_,
		_w6964_,
		_w6966_,
		_w7720_
	);
	LUT2 #(
		.INIT('h1)
	) name7687 (
		_w7719_,
		_w7720_,
		_w7721_
	);
	LUT2 #(
		.INIT('h4)
	) name7688 (
		_w7718_,
		_w7721_,
		_w7722_
	);
	LUT3 #(
		.INIT('h9a)
	) name7689 (
		\a[26] ,
		_w7717_,
		_w7722_,
		_w7723_
	);
	LUT3 #(
		.INIT('hd4)
	) name7690 (
		_w7709_,
		_w7716_,
		_w7723_,
		_w7724_
	);
	LUT4 #(
		.INIT('he100)
	) name7691 (
		_w7560_,
		_w7662_,
		_w7664_,
		_w7707_,
		_w7725_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name7692 (
		_w7560_,
		_w7662_,
		_w7664_,
		_w7707_,
		_w7726_
	);
	LUT3 #(
		.INIT('h54)
	) name7693 (
		_w7708_,
		_w7724_,
		_w7725_,
		_w7727_
	);
	LUT3 #(
		.INIT('h96)
	) name7694 (
		_w7665_,
		_w7666_,
		_w7672_,
		_w7728_
	);
	LUT4 #(
		.INIT('h02a8)
	) name7695 (
		_w37_,
		_w7004_,
		_w7127_,
		_w7128_,
		_w7729_
	);
	LUT4 #(
		.INIT('h04c8)
	) name7696 (
		_w2622_,
		_w3262_,
		_w6978_,
		_w6980_,
		_w7730_
	);
	LUT3 #(
		.INIT('h82)
	) name7697 (
		_w3214_,
		_w2872_,
		_w6975_,
		_w7731_
	);
	LUT3 #(
		.INIT('h07)
	) name7698 (
		_w3249_,
		_w7002_,
		_w7731_,
		_w7732_
	);
	LUT2 #(
		.INIT('h4)
	) name7699 (
		_w7730_,
		_w7732_,
		_w7733_
	);
	LUT3 #(
		.INIT('h9a)
	) name7700 (
		\a[23] ,
		_w7729_,
		_w7733_,
		_w7734_
	);
	LUT3 #(
		.INIT('hb2)
	) name7701 (
		_w7727_,
		_w7728_,
		_w7734_,
		_w7735_
	);
	LUT3 #(
		.INIT('h82)
	) name7702 (
		_w3312_,
		_w7135_,
		_w7172_,
		_w7736_
	);
	LUT3 #(
		.INIT('h28)
	) name7703 (
		_w3654_,
		_w7136_,
		_w7168_,
		_w7737_
	);
	LUT2 #(
		.INIT('h8)
	) name7704 (
		_w3311_,
		_w6996_,
		_w7738_
	);
	LUT4 #(
		.INIT('h04c8)
	) name7705 (
		_w2411_,
		_w3645_,
		_w6983_,
		_w6993_,
		_w7739_
	);
	LUT2 #(
		.INIT('h1)
	) name7706 (
		_w7738_,
		_w7739_,
		_w7740_
	);
	LUT2 #(
		.INIT('h4)
	) name7707 (
		_w7737_,
		_w7740_,
		_w7741_
	);
	LUT3 #(
		.INIT('h9a)
	) name7708 (
		\a[20] ,
		_w7736_,
		_w7741_,
		_w7742_
	);
	LUT3 #(
		.INIT('hd4)
	) name7709 (
		_w7703_,
		_w7735_,
		_w7742_,
		_w7743_
	);
	LUT4 #(
		.INIT('h0445)
	) name7710 (
		_w7701_,
		_w7703_,
		_w7735_,
		_w7742_,
		_w7744_
	);
	LUT4 #(
		.INIT('h6665)
	) name7711 (
		_w7506_,
		_w7674_,
		_w7675_,
		_w7682_,
		_w7745_
	);
	LUT4 #(
		.INIT('ha220)
	) name7712 (
		_w7701_,
		_w7703_,
		_w7735_,
		_w7742_,
		_w7746_
	);
	LUT4 #(
		.INIT('h599a)
	) name7713 (
		_w7701_,
		_w7703_,
		_w7735_,
		_w7742_,
		_w7747_
	);
	LUT3 #(
		.INIT('h51)
	) name7714 (
		_w7744_,
		_w7745_,
		_w7746_,
		_w7748_
	);
	LUT4 #(
		.INIT('he11e)
	) name7715 (
		_w7505_,
		_w7683_,
		_w7684_,
		_w7691_,
		_w7749_
	);
	LUT4 #(
		.INIT('h0071)
	) name7716 (
		_w7701_,
		_w7743_,
		_w7745_,
		_w7749_,
		_w7750_
	);
	LUT2 #(
		.INIT('h6)
	) name7717 (
		_w7745_,
		_w7747_,
		_w7751_
	);
	LUT4 #(
		.INIT('h028a)
	) name7718 (
		_w3709_,
		_w7136_,
		_w7166_,
		_w7167_,
		_w7752_
	);
	LUT4 #(
		.INIT('h87e1)
	) name7719 (
		\a[14] ,
		\a[15] ,
		\a[16] ,
		\a[17] ,
		_w7753_
	);
	LUT3 #(
		.INIT('h0b)
	) name7720 (
		_w7136_,
		_w7166_,
		_w7753_,
		_w7754_
	);
	LUT2 #(
		.INIT('h1)
	) name7721 (
		_w7752_,
		_w7754_,
		_w7755_
	);
	LUT4 #(
		.INIT('h5700)
	) name7722 (
		_w3710_,
		_w7418_,
		_w7419_,
		_w7755_,
		_w7756_
	);
	LUT2 #(
		.INIT('h6)
	) name7723 (
		\a[17] ,
		_w7756_,
		_w7757_
	);
	LUT4 #(
		.INIT('h02a8)
	) name7724 (
		_w3214_,
		_w2983_,
		_w6972_,
		_w6974_,
		_w7758_
	);
	LUT4 #(
		.INIT('h007b)
	) name7725 (
		_w2872_,
		_w3249_,
		_w6975_,
		_w7758_,
		_w7759_
	);
	LUT3 #(
		.INIT('h70)
	) name7726 (
		_w3262_,
		_w7002_,
		_w7759_,
		_w7760_
	);
	LUT4 #(
		.INIT('h95aa)
	) name7727 (
		\a[23] ,
		_w37_,
		_w7426_,
		_w7760_,
		_w7761_
	);
	LUT3 #(
		.INIT('h09)
	) name7728 (
		_w7724_,
		_w7726_,
		_w7761_,
		_w7762_
	);
	LUT3 #(
		.INIT('h60)
	) name7729 (
		_w7724_,
		_w7726_,
		_w7761_,
		_w7763_
	);
	LUT3 #(
		.INIT('h96)
	) name7730 (
		_w7724_,
		_w7726_,
		_w7761_,
		_w7764_
	);
	LUT3 #(
		.INIT('h96)
	) name7731 (
		_w7709_,
		_w7716_,
		_w7723_,
		_w7765_
	);
	LUT2 #(
		.INIT('h9)
	) name7732 (
		_w7655_,
		_w7661_,
		_w7766_
	);
	LUT4 #(
		.INIT('h54ab)
	) name7733 (
		_w7638_,
		_w7639_,
		_w7646_,
		_w7647_,
		_w7767_
	);
	LUT3 #(
		.INIT('h82)
	) name7734 (
		_w377_,
		_w7099_,
		_w7101_,
		_w7768_
	);
	LUT3 #(
		.INIT('h82)
	) name7735 (
		_w2527_,
		_w4030_,
		_w6952_,
		_w7769_
	);
	LUT2 #(
		.INIT('h8)
	) name7736 (
		_w376_,
		_w7032_,
		_w7770_
	);
	LUT4 #(
		.INIT('h2228)
	) name7737 (
		_w2407_,
		_w4099_,
		_w4378_,
		_w6951_,
		_w7771_
	);
	LUT2 #(
		.INIT('h1)
	) name7738 (
		_w7770_,
		_w7771_,
		_w7772_
	);
	LUT2 #(
		.INIT('h4)
	) name7739 (
		_w7769_,
		_w7772_,
		_w7773_
	);
	LUT2 #(
		.INIT('h4)
	) name7740 (
		_w7768_,
		_w7773_,
		_w7774_
	);
	LUT3 #(
		.INIT('h82)
	) name7741 (
		_w2550_,
		_w7105_,
		_w7107_,
		_w7775_
	);
	LUT3 #(
		.INIT('h82)
	) name7742 (
		_w2854_,
		_w3706_,
		_w6957_,
		_w7776_
	);
	LUT2 #(
		.INIT('h8)
	) name7743 (
		_w2549_,
		_w7026_,
		_w7777_
	);
	LUT4 #(
		.INIT('h02a8)
	) name7744 (
		_w2617_,
		_w3882_,
		_w6954_,
		_w6956_,
		_w7778_
	);
	LUT2 #(
		.INIT('h1)
	) name7745 (
		_w7777_,
		_w7778_,
		_w7779_
	);
	LUT2 #(
		.INIT('h4)
	) name7746 (
		_w7776_,
		_w7779_,
		_w7780_
	);
	LUT3 #(
		.INIT('h9a)
	) name7747 (
		\a[29] ,
		_w7775_,
		_w7780_,
		_w7781_
	);
	LUT3 #(
		.INIT('hd4)
	) name7748 (
		_w7767_,
		_w7774_,
		_w7781_,
		_w7782_
	);
	LUT2 #(
		.INIT('h9)
	) name7749 (
		_w7648_,
		_w7650_,
		_w7783_
	);
	LUT4 #(
		.INIT('h02a8)
	) name7750 (
		_w2549_,
		_w3882_,
		_w6954_,
		_w6956_,
		_w7784_
	);
	LUT4 #(
		.INIT('h007d)
	) name7751 (
		_w2617_,
		_w3706_,
		_w6957_,
		_w7784_,
		_w7785_
	);
	LUT3 #(
		.INIT('h70)
	) name7752 (
		_w2854_,
		_w7020_,
		_w7785_,
		_w7786_
	);
	LUT4 #(
		.INIT('h95aa)
	) name7753 (
		\a[29] ,
		_w2550_,
		_w7465_,
		_w7786_,
		_w7787_
	);
	LUT3 #(
		.INIT('hb2)
	) name7754 (
		_w7782_,
		_w7783_,
		_w7787_,
		_w7788_
	);
	LUT4 #(
		.INIT('h02a8)
	) name7755 (
		_w2875_,
		_w7016_,
		_w7115_,
		_w7116_,
		_w7789_
	);
	LUT4 #(
		.INIT('h02a8)
	) name7756 (
		_w2986_,
		_w3257_,
		_w6964_,
		_w6966_,
		_w7790_
	);
	LUT3 #(
		.INIT('h82)
	) name7757 (
		_w2874_,
		_w6960_,
		_w6962_,
		_w7791_
	);
	LUT3 #(
		.INIT('h07)
	) name7758 (
		_w2975_,
		_w7014_,
		_w7791_,
		_w7792_
	);
	LUT2 #(
		.INIT('h4)
	) name7759 (
		_w7790_,
		_w7792_,
		_w7793_
	);
	LUT3 #(
		.INIT('h9a)
	) name7760 (
		\a[26] ,
		_w7789_,
		_w7793_,
		_w7794_
	);
	LUT3 #(
		.INIT('hd4)
	) name7761 (
		_w7766_,
		_w7788_,
		_w7794_,
		_w7795_
	);
	LUT3 #(
		.INIT('h82)
	) name7762 (
		_w37_,
		_w7123_,
		_w7125_,
		_w7796_
	);
	LUT3 #(
		.INIT('h84)
	) name7763 (
		_w2872_,
		_w3262_,
		_w6975_,
		_w7797_
	);
	LUT2 #(
		.INIT('h8)
	) name7764 (
		_w3214_,
		_w7008_,
		_w7798_
	);
	LUT4 #(
		.INIT('h04c8)
	) name7765 (
		_w2983_,
		_w3249_,
		_w6972_,
		_w6974_,
		_w7799_
	);
	LUT2 #(
		.INIT('h1)
	) name7766 (
		_w7798_,
		_w7799_,
		_w7800_
	);
	LUT2 #(
		.INIT('h4)
	) name7767 (
		_w7797_,
		_w7800_,
		_w7801_
	);
	LUT3 #(
		.INIT('h9a)
	) name7768 (
		\a[23] ,
		_w7796_,
		_w7801_,
		_w7802_
	);
	LUT3 #(
		.INIT('hd4)
	) name7769 (
		_w7765_,
		_w7795_,
		_w7802_,
		_w7803_
	);
	LUT3 #(
		.INIT('h54)
	) name7770 (
		_w7762_,
		_w7763_,
		_w7803_,
		_w7804_
	);
	LUT3 #(
		.INIT('h69)
	) name7771 (
		_w7727_,
		_w7728_,
		_w7734_,
		_w7805_
	);
	LUT4 #(
		.INIT('h02a8)
	) name7772 (
		_w3312_,
		_w6998_,
		_w7133_,
		_w7134_,
		_w7806_
	);
	LUT4 #(
		.INIT('h04c8)
	) name7773 (
		_w2411_,
		_w3654_,
		_w6983_,
		_w6993_,
		_w7807_
	);
	LUT3 #(
		.INIT('h84)
	) name7774 (
		_w2546_,
		_w3311_,
		_w6981_,
		_w7808_
	);
	LUT3 #(
		.INIT('h07)
	) name7775 (
		_w3645_,
		_w6996_,
		_w7808_,
		_w7809_
	);
	LUT2 #(
		.INIT('h4)
	) name7776 (
		_w7807_,
		_w7809_,
		_w7810_
	);
	LUT3 #(
		.INIT('h9a)
	) name7777 (
		\a[20] ,
		_w7806_,
		_w7810_,
		_w7811_
	);
	LUT4 #(
		.INIT('h0115)
	) name7778 (
		_w7757_,
		_w7804_,
		_w7805_,
		_w7811_,
		_w7812_
	);
	LUT4 #(
		.INIT('ha880)
	) name7779 (
		_w7757_,
		_w7804_,
		_w7805_,
		_w7811_,
		_w7813_
	);
	LUT3 #(
		.INIT('h96)
	) name7780 (
		_w7703_,
		_w7735_,
		_w7742_,
		_w7814_
	);
	LUT3 #(
		.INIT('h45)
	) name7781 (
		_w7812_,
		_w7813_,
		_w7814_,
		_w7815_
	);
	LUT2 #(
		.INIT('h2)
	) name7782 (
		_w7751_,
		_w7815_,
		_w7816_
	);
	LUT4 #(
		.INIT('h566a)
	) name7783 (
		_w7757_,
		_w7804_,
		_w7805_,
		_w7811_,
		_w7817_
	);
	LUT2 #(
		.INIT('h6)
	) name7784 (
		_w7814_,
		_w7817_,
		_w7818_
	);
	LUT4 #(
		.INIT('h04c8)
	) name7785 (
		_w2622_,
		_w3311_,
		_w6978_,
		_w6980_,
		_w7819_
	);
	LUT4 #(
		.INIT('h007b)
	) name7786 (
		_w2546_,
		_w3645_,
		_w6981_,
		_w7819_,
		_w7820_
	);
	LUT3 #(
		.INIT('h70)
	) name7787 (
		_w3654_,
		_w6996_,
		_w7820_,
		_w7821_
	);
	LUT4 #(
		.INIT('h95aa)
	) name7788 (
		\a[20] ,
		_w3312_,
		_w7500_,
		_w7821_,
		_w7822_
	);
	LUT3 #(
		.INIT('h09)
	) name7789 (
		_w7764_,
		_w7803_,
		_w7822_,
		_w7823_
	);
	LUT3 #(
		.INIT('h60)
	) name7790 (
		_w7764_,
		_w7803_,
		_w7822_,
		_w7824_
	);
	LUT3 #(
		.INIT('h96)
	) name7791 (
		_w7764_,
		_w7803_,
		_w7822_,
		_w7825_
	);
	LUT3 #(
		.INIT('h96)
	) name7792 (
		_w7765_,
		_w7795_,
		_w7802_,
		_w7826_
	);
	LUT4 #(
		.INIT('h2228)
	) name7793 (
		_w2874_,
		_w3409_,
		_w3650_,
		_w6959_,
		_w7827_
	);
	LUT4 #(
		.INIT('h007d)
	) name7794 (
		_w2975_,
		_w6960_,
		_w6962_,
		_w7827_,
		_w7828_
	);
	LUT3 #(
		.INIT('h70)
	) name7795 (
		_w2986_,
		_w7014_,
		_w7828_,
		_w7829_
	);
	LUT4 #(
		.INIT('h95aa)
	) name7796 (
		\a[26] ,
		_w2875_,
		_w7291_,
		_w7829_,
		_w7830_
	);
	LUT4 #(
		.INIT('h0096)
	) name7797 (
		_w7782_,
		_w7783_,
		_w7787_,
		_w7830_,
		_w7831_
	);
	LUT4 #(
		.INIT('h9669)
	) name7798 (
		_w7782_,
		_w7783_,
		_w7787_,
		_w7830_,
		_w7832_
	);
	LUT2 #(
		.INIT('h9)
	) name7799 (
		_w7640_,
		_w7646_,
		_w7833_
	);
	LUT2 #(
		.INIT('h4)
	) name7800 (
		_w241_,
		_w1362_,
		_w7834_
	);
	LUT3 #(
		.INIT('h10)
	) name7801 (
		_w77_,
		_w241_,
		_w1362_,
		_w7835_
	);
	LUT3 #(
		.INIT('h80)
	) name7802 (
		_w260_,
		_w1991_,
		_w7624_,
		_w7836_
	);
	LUT3 #(
		.INIT('h80)
	) name7803 (
		_w703_,
		_w7835_,
		_w7836_,
		_w7837_
	);
	LUT4 #(
		.INIT('h0777)
	) name7804 (
		_w122_,
		_w85_,
		_w43_,
		_w44_,
		_w7838_
	);
	LUT4 #(
		.INIT('h0800)
	) name7805 (
		_w116_,
		_w296_,
		_w463_,
		_w7838_,
		_w7839_
	);
	LUT4 #(
		.INIT('h4000)
	) name7806 (
		_w202_,
		_w969_,
		_w1359_,
		_w3549_,
		_w7840_
	);
	LUT4 #(
		.INIT('h8000)
	) name7807 (
		_w745_,
		_w748_,
		_w7839_,
		_w7840_,
		_w7841_
	);
	LUT4 #(
		.INIT('h8000)
	) name7808 (
		_w1731_,
		_w1740_,
		_w7837_,
		_w7841_,
		_w7842_
	);
	LUT2 #(
		.INIT('h8)
	) name7809 (
		_w1817_,
		_w7842_,
		_w7843_
	);
	LUT3 #(
		.INIT('h01)
	) name7810 (
		\a[0] ,
		\a[1] ,
		\a[2] ,
		_w7844_
	);
	LUT4 #(
		.INIT('hdf9a)
	) name7811 (
		\a[2] ,
		_w7136_,
		_w7166_,
		_w7844_,
		_w7845_
	);
	LUT4 #(
		.INIT('h153f)
	) name7812 (
		_w38_,
		_w52_,
		_w72_,
		_w184_,
		_w7846_
	);
	LUT2 #(
		.INIT('h4)
	) name7813 (
		_w432_,
		_w7846_,
		_w7847_
	);
	LUT4 #(
		.INIT('h8000)
	) name7814 (
		_w795_,
		_w906_,
		_w990_,
		_w1342_,
		_w7848_
	);
	LUT3 #(
		.INIT('h80)
	) name7815 (
		_w1703_,
		_w2102_,
		_w2516_,
		_w7849_
	);
	LUT4 #(
		.INIT('h8000)
	) name7816 (
		_w736_,
		_w7847_,
		_w7849_,
		_w7848_,
		_w7850_
	);
	LUT4 #(
		.INIT('h153f)
	) name7817 (
		_w52_,
		_w59_,
		_w236_,
		_w430_,
		_w7851_
	);
	LUT4 #(
		.INIT('h8000)
	) name7818 (
		_w834_,
		_w7571_,
		_w7572_,
		_w7851_,
		_w7852_
	);
	LUT3 #(
		.INIT('h40)
	) name7819 (
		_w223_,
		_w953_,
		_w1761_,
		_w7853_
	);
	LUT3 #(
		.INIT('h80)
	) name7820 (
		_w2575_,
		_w7852_,
		_w7853_,
		_w7854_
	);
	LUT4 #(
		.INIT('h4000)
	) name7821 (
		_w247_,
		_w902_,
		_w964_,
		_w1961_,
		_w7855_
	);
	LUT4 #(
		.INIT('h4000)
	) name7822 (
		_w431_,
		_w650_,
		_w1184_,
		_w2790_,
		_w7856_
	);
	LUT4 #(
		.INIT('h8000)
	) name7823 (
		_w2168_,
		_w2171_,
		_w7855_,
		_w7856_,
		_w7857_
	);
	LUT3 #(
		.INIT('h80)
	) name7824 (
		_w7850_,
		_w7854_,
		_w7857_,
		_w7858_
	);
	LUT4 #(
		.INIT('h8000)
	) name7825 (
		_w931_,
		_w1576_,
		_w2177_,
		_w2625_,
		_w7859_
	);
	LUT4 #(
		.INIT('h153f)
	) name7826 (
		_w47_,
		_w39_,
		_w44_,
		_w378_,
		_w7860_
	);
	LUT4 #(
		.INIT('h4000)
	) name7827 (
		_w308_,
		_w675_,
		_w1012_,
		_w7860_,
		_w7861_
	);
	LUT4 #(
		.INIT('h8000)
	) name7828 (
		_w3955_,
		_w4231_,
		_w7859_,
		_w7861_,
		_w7862_
	);
	LUT4 #(
		.INIT('h8000)
	) name7829 (
		_w2695_,
		_w2697_,
		_w7522_,
		_w7525_,
		_w7863_
	);
	LUT2 #(
		.INIT('h8)
	) name7830 (
		_w7862_,
		_w7863_,
		_w7864_
	);
	LUT2 #(
		.INIT('h8)
	) name7831 (
		_w7858_,
		_w7864_,
		_w7865_
	);
	LUT4 #(
		.INIT('h87e1)
	) name7832 (
		\a[2] ,
		\a[3] ,
		\a[4] ,
		\a[5] ,
		_w7866_
	);
	LUT4 #(
		.INIT('h8001)
	) name7833 (
		\a[2] ,
		\a[3] ,
		\a[4] ,
		\a[5] ,
		_w7867_
	);
	LUT4 #(
		.INIT('h559a)
	) name7834 (
		\a[5] ,
		_w7136_,
		_w7166_,
		_w7867_,
		_w7868_
	);
	LUT3 #(
		.INIT('h4d)
	) name7835 (
		_w7845_,
		_w7865_,
		_w7868_,
		_w7869_
	);
	LUT4 #(
		.INIT('h8a08)
	) name7836 (
		_w7614_,
		_w7845_,
		_w7865_,
		_w7868_,
		_w7870_
	);
	LUT4 #(
		.INIT('h1051)
	) name7837 (
		_w7614_,
		_w7845_,
		_w7865_,
		_w7868_,
		_w7871_
	);
	LUT4 #(
		.INIT('h65a6)
	) name7838 (
		_w7614_,
		_w7845_,
		_w7865_,
		_w7868_,
		_w7872_
	);
	LUT4 #(
		.INIT('h02a8)
	) name7839 (
		_w377_,
		_w7040_,
		_w7091_,
		_w7092_,
		_w7873_
	);
	LUT4 #(
		.INIT('h02a8)
	) name7840 (
		_w2527_,
		_w4695_,
		_w6944_,
		_w6946_,
		_w7874_
	);
	LUT3 #(
		.INIT('h82)
	) name7841 (
		_w376_,
		_w6940_,
		_w6942_,
		_w7875_
	);
	LUT3 #(
		.INIT('h07)
	) name7842 (
		_w2407_,
		_w7038_,
		_w7875_,
		_w7876_
	);
	LUT2 #(
		.INIT('h4)
	) name7843 (
		_w7874_,
		_w7876_,
		_w7877_
	);
	LUT2 #(
		.INIT('h4)
	) name7844 (
		_w7873_,
		_w7877_,
		_w7878_
	);
	LUT4 #(
		.INIT('h953f)
	) name7845 (
		_w1817_,
		_w2036_,
		_w7613_,
		_w7842_,
		_w7879_
	);
	LUT4 #(
		.INIT('hd554)
	) name7846 (
		_w7614_,
		_w7843_,
		_w7869_,
		_w7878_,
		_w7880_
	);
	LUT2 #(
		.INIT('h6)
	) name7847 (
		_w7634_,
		_w7636_,
		_w7881_
	);
	LUT4 #(
		.INIT('h54ab)
	) name7848 (
		_w7036_,
		_w7093_,
		_w7094_,
		_w7096_,
		_w7882_
	);
	LUT4 #(
		.INIT('h02a8)
	) name7849 (
		_w376_,
		_w4695_,
		_w6944_,
		_w6946_,
		_w7883_
	);
	LUT4 #(
		.INIT('h007d)
	) name7850 (
		_w2407_,
		_w6947_,
		_w6949_,
		_w7883_,
		_w7884_
	);
	LUT3 #(
		.INIT('h70)
	) name7851 (
		_w2527_,
		_w7032_,
		_w7884_,
		_w7885_
	);
	LUT3 #(
		.INIT('h70)
	) name7852 (
		_w377_,
		_w7882_,
		_w7885_,
		_w7886_
	);
	LUT3 #(
		.INIT('hb2)
	) name7853 (
		_w7880_,
		_w7881_,
		_w7886_,
		_w7887_
	);
	LUT4 #(
		.INIT('h20a2)
	) name7854 (
		_w7833_,
		_w7880_,
		_w7881_,
		_w7886_,
		_w7888_
	);
	LUT4 #(
		.INIT('h4504)
	) name7855 (
		_w7833_,
		_w7880_,
		_w7881_,
		_w7886_,
		_w7889_
	);
	LUT4 #(
		.INIT('h9a59)
	) name7856 (
		_w7833_,
		_w7880_,
		_w7881_,
		_w7886_,
		_w7890_
	);
	LUT4 #(
		.INIT('h02a8)
	) name7857 (
		_w2550_,
		_w7028_,
		_w7103_,
		_w7104_,
		_w7891_
	);
	LUT4 #(
		.INIT('h02a8)
	) name7858 (
		_w2854_,
		_w3882_,
		_w6954_,
		_w6956_,
		_w7892_
	);
	LUT3 #(
		.INIT('h82)
	) name7859 (
		_w2549_,
		_w4030_,
		_w6952_,
		_w7893_
	);
	LUT3 #(
		.INIT('h07)
	) name7860 (
		_w2617_,
		_w7026_,
		_w7893_,
		_w7894_
	);
	LUT2 #(
		.INIT('h4)
	) name7861 (
		_w7892_,
		_w7894_,
		_w7895_
	);
	LUT3 #(
		.INIT('h9a)
	) name7862 (
		\a[29] ,
		_w7891_,
		_w7895_,
		_w7896_
	);
	LUT3 #(
		.INIT('h54)
	) name7863 (
		_w7888_,
		_w7889_,
		_w7896_,
		_w7897_
	);
	LUT3 #(
		.INIT('h96)
	) name7864 (
		_w7767_,
		_w7774_,
		_w7781_,
		_w7898_
	);
	LUT4 #(
		.INIT('h2b00)
	) name7865 (
		_w7833_,
		_w7887_,
		_w7896_,
		_w7898_,
		_w7899_
	);
	LUT4 #(
		.INIT('h00d4)
	) name7866 (
		_w7833_,
		_w7887_,
		_w7896_,
		_w7898_,
		_w7900_
	);
	LUT3 #(
		.INIT('h82)
	) name7867 (
		_w2875_,
		_w7111_,
		_w7113_,
		_w7901_
	);
	LUT3 #(
		.INIT('h82)
	) name7868 (
		_w2986_,
		_w6960_,
		_w6962_,
		_w7902_
	);
	LUT2 #(
		.INIT('h8)
	) name7869 (
		_w2874_,
		_w7020_,
		_w7903_
	);
	LUT4 #(
		.INIT('h2228)
	) name7870 (
		_w2975_,
		_w3409_,
		_w3650_,
		_w6959_,
		_w7904_
	);
	LUT2 #(
		.INIT('h1)
	) name7871 (
		_w7903_,
		_w7904_,
		_w7905_
	);
	LUT2 #(
		.INIT('h4)
	) name7872 (
		_w7902_,
		_w7905_,
		_w7906_
	);
	LUT3 #(
		.INIT('h9a)
	) name7873 (
		\a[26] ,
		_w7901_,
		_w7906_,
		_w7907_
	);
	LUT4 #(
		.INIT('h20a2)
	) name7874 (
		_w7832_,
		_w7897_,
		_w7898_,
		_w7907_,
		_w7908_
	);
	LUT3 #(
		.INIT('h96)
	) name7875 (
		_w7766_,
		_w7788_,
		_w7794_,
		_w7909_
	);
	LUT4 #(
		.INIT('h02a8)
	) name7876 (
		_w37_,
		_w7010_,
		_w7121_,
		_w7122_,
		_w7910_
	);
	LUT4 #(
		.INIT('h04c8)
	) name7877 (
		_w2983_,
		_w3262_,
		_w6972_,
		_w6974_,
		_w7911_
	);
	LUT3 #(
		.INIT('h82)
	) name7878 (
		_w3214_,
		_w6967_,
		_w6969_,
		_w7912_
	);
	LUT3 #(
		.INIT('h07)
	) name7879 (
		_w3249_,
		_w7008_,
		_w7912_,
		_w7913_
	);
	LUT2 #(
		.INIT('h4)
	) name7880 (
		_w7911_,
		_w7913_,
		_w7914_
	);
	LUT3 #(
		.INIT('h9a)
	) name7881 (
		\a[23] ,
		_w7910_,
		_w7914_,
		_w7915_
	);
	LUT4 #(
		.INIT('h1f01)
	) name7882 (
		_w7831_,
		_w7908_,
		_w7909_,
		_w7915_,
		_w7916_
	);
	LUT3 #(
		.INIT('h82)
	) name7883 (
		_w3312_,
		_w7129_,
		_w7131_,
		_w7917_
	);
	LUT3 #(
		.INIT('h84)
	) name7884 (
		_w2546_,
		_w3654_,
		_w6981_,
		_w7918_
	);
	LUT2 #(
		.INIT('h8)
	) name7885 (
		_w3311_,
		_w7002_,
		_w7919_
	);
	LUT4 #(
		.INIT('h04c8)
	) name7886 (
		_w2622_,
		_w3645_,
		_w6978_,
		_w6980_,
		_w7920_
	);
	LUT2 #(
		.INIT('h1)
	) name7887 (
		_w7919_,
		_w7920_,
		_w7921_
	);
	LUT2 #(
		.INIT('h4)
	) name7888 (
		_w7918_,
		_w7921_,
		_w7922_
	);
	LUT3 #(
		.INIT('h9a)
	) name7889 (
		\a[20] ,
		_w7917_,
		_w7922_,
		_w7923_
	);
	LUT3 #(
		.INIT('hd4)
	) name7890 (
		_w7826_,
		_w7916_,
		_w7923_,
		_w7924_
	);
	LUT3 #(
		.INIT('h54)
	) name7891 (
		_w7823_,
		_w7824_,
		_w7924_,
		_w7925_
	);
	LUT3 #(
		.INIT('h69)
	) name7892 (
		_w7804_,
		_w7805_,
		_w7811_,
		_w7926_
	);
	LUT4 #(
		.INIT('h0a02)
	) name7893 (
		_w3710_,
		_w7169_,
		_w7419_,
		_w7686_,
		_w7927_
	);
	LUT3 #(
		.INIT('h28)
	) name7894 (
		_w3709_,
		_w7136_,
		_w7168_,
		_w7928_
	);
	LUT3 #(
		.INIT('h40)
	) name7895 (
		_w3886_,
		_w7136_,
		_w7167_,
		_w7929_
	);
	LUT3 #(
		.INIT('h31)
	) name7896 (
		_w7754_,
		_w7928_,
		_w7929_,
		_w7930_
	);
	LUT3 #(
		.INIT('h9a)
	) name7897 (
		\a[17] ,
		_w7927_,
		_w7930_,
		_w7931_
	);
	LUT3 #(
		.INIT('hb2)
	) name7898 (
		_w7925_,
		_w7926_,
		_w7931_,
		_w7932_
	);
	LUT2 #(
		.INIT('h2)
	) name7899 (
		_w7818_,
		_w7932_,
		_w7933_
	);
	LUT2 #(
		.INIT('h4)
	) name7900 (
		_w7818_,
		_w7932_,
		_w7934_
	);
	LUT2 #(
		.INIT('h9)
	) name7901 (
		_w7818_,
		_w7932_,
		_w7935_
	);
	LUT3 #(
		.INIT('h28)
	) name7902 (
		_w3877_,
		_w7136_,
		_w7168_,
		_w7936_
	);
	LUT4 #(
		.INIT('h028a)
	) name7903 (
		_w3886_,
		_w7136_,
		_w7166_,
		_w7167_,
		_w7937_
	);
	LUT4 #(
		.INIT('h04c8)
	) name7904 (
		_w2411_,
		_w3709_,
		_w6983_,
		_w6993_,
		_w7938_
	);
	LUT3 #(
		.INIT('h01)
	) name7905 (
		_w7937_,
		_w7938_,
		_w7936_,
		_w7939_
	);
	LUT4 #(
		.INIT('h95aa)
	) name7906 (
		\a[17] ,
		_w3710_,
		_w7696_,
		_w7939_,
		_w7940_
	);
	LUT3 #(
		.INIT('h96)
	) name7907 (
		_w7826_,
		_w7916_,
		_w7923_,
		_w7941_
	);
	LUT4 #(
		.INIT('h6665)
	) name7908 (
		_w7832_,
		_w7899_,
		_w7900_,
		_w7907_,
		_w7942_
	);
	LUT4 #(
		.INIT('h02a8)
	) name7909 (
		_w3214_,
		_w3257_,
		_w6964_,
		_w6966_,
		_w7943_
	);
	LUT4 #(
		.INIT('h007d)
	) name7910 (
		_w3249_,
		_w6967_,
		_w6969_,
		_w7943_,
		_w7944_
	);
	LUT3 #(
		.INIT('h70)
	) name7911 (
		_w3262_,
		_w7008_,
		_w7944_,
		_w7945_
	);
	LUT4 #(
		.INIT('h95aa)
	) name7912 (
		\a[23] ,
		_w37_,
		_w7403_,
		_w7945_,
		_w7946_
	);
	LUT2 #(
		.INIT('h2)
	) name7913 (
		_w7942_,
		_w7946_,
		_w7947_
	);
	LUT2 #(
		.INIT('h9)
	) name7914 (
		_w7942_,
		_w7946_,
		_w7948_
	);
	LUT4 #(
		.INIT('h54ab)
	) name7915 (
		_w7888_,
		_w7889_,
		_w7896_,
		_w7898_,
		_w7949_
	);
	LUT2 #(
		.INIT('h9)
	) name7916 (
		_w7907_,
		_w7949_,
		_w7950_
	);
	LUT4 #(
		.INIT('h2228)
	) name7917 (
		_w2549_,
		_w4099_,
		_w4378_,
		_w6951_,
		_w7951_
	);
	LUT4 #(
		.INIT('h007d)
	) name7918 (
		_w2617_,
		_w4030_,
		_w6952_,
		_w7951_,
		_w7952_
	);
	LUT3 #(
		.INIT('h70)
	) name7919 (
		_w2854_,
		_w7026_,
		_w7952_,
		_w7953_
	);
	LUT4 #(
		.INIT('h95aa)
	) name7920 (
		\a[29] ,
		_w2550_,
		_w7562_,
		_w7953_,
		_w7954_
	);
	LUT4 #(
		.INIT('h0096)
	) name7921 (
		_w7880_,
		_w7881_,
		_w7886_,
		_w7954_,
		_w7955_
	);
	LUT4 #(
		.INIT('h54ab)
	) name7922 (
		_w7870_,
		_w7871_,
		_w7878_,
		_w7879_,
		_w7956_
	);
	LUT3 #(
		.INIT('h82)
	) name7923 (
		_w377_,
		_w7093_,
		_w7095_,
		_w7957_
	);
	LUT3 #(
		.INIT('h82)
	) name7924 (
		_w2527_,
		_w6947_,
		_w6949_,
		_w7958_
	);
	LUT2 #(
		.INIT('h8)
	) name7925 (
		_w376_,
		_w7038_,
		_w7959_
	);
	LUT4 #(
		.INIT('h02a8)
	) name7926 (
		_w2407_,
		_w4695_,
		_w6944_,
		_w6946_,
		_w7960_
	);
	LUT2 #(
		.INIT('h1)
	) name7927 (
		_w7959_,
		_w7960_,
		_w7961_
	);
	LUT2 #(
		.INIT('h4)
	) name7928 (
		_w7958_,
		_w7961_,
		_w7962_
	);
	LUT2 #(
		.INIT('h4)
	) name7929 (
		_w7957_,
		_w7962_,
		_w7963_
	);
	LUT2 #(
		.INIT('h2)
	) name7930 (
		_w7956_,
		_w7963_,
		_w7964_
	);
	LUT4 #(
		.INIT('h8000)
	) name7931 (
		_w1774_,
		_w1877_,
		_w2000_,
		_w2807_,
		_w7965_
	);
	LUT3 #(
		.INIT('h1f)
	) name7932 (
		_w39_,
		_w43_,
		_w93_,
		_w7966_
	);
	LUT3 #(
		.INIT('h57)
	) name7933 (
		_w55_,
		_w176_,
		_w430_,
		_w7967_
	);
	LUT4 #(
		.INIT('h8000)
	) name7934 (
		_w894_,
		_w1649_,
		_w7966_,
		_w7967_,
		_w7968_
	);
	LUT4 #(
		.INIT('h8000)
	) name7935 (
		_w1370_,
		_w2224_,
		_w7965_,
		_w7968_,
		_w7969_
	);
	LUT3 #(
		.INIT('h80)
	) name7936 (
		_w569_,
		_w2456_,
		_w7969_,
		_w7970_
	);
	LUT2 #(
		.INIT('h8)
	) name7937 (
		_w2648_,
		_w7970_,
		_w7971_
	);
	LUT2 #(
		.INIT('h1)
	) name7938 (
		_w7845_,
		_w7971_,
		_w7972_
	);
	LUT3 #(
		.INIT('h40)
	) name7939 (
		_w420_,
		_w908_,
		_w7297_,
		_w7973_
	);
	LUT4 #(
		.INIT('h8000)
	) name7940 (
		_w1687_,
		_w1837_,
		_w3022_,
		_w7196_,
		_w7974_
	);
	LUT3 #(
		.INIT('h80)
	) name7941 (
		_w7144_,
		_w7973_,
		_w7974_,
		_w7975_
	);
	LUT4 #(
		.INIT('h153f)
	) name7942 (
		_w38_,
		_w67_,
		_w72_,
		_w259_,
		_w7976_
	);
	LUT4 #(
		.INIT('h8000)
	) name7943 (
		_w54_,
		_w957_,
		_w1439_,
		_w7976_,
		_w7977_
	);
	LUT4 #(
		.INIT('h4000)
	) name7944 (
		_w128_,
		_w254_,
		_w1013_,
		_w1374_,
		_w7978_
	);
	LUT4 #(
		.INIT('h8000)
	) name7945 (
		_w1044_,
		_w1048_,
		_w7977_,
		_w7978_,
		_w7979_
	);
	LUT3 #(
		.INIT('h80)
	) name7946 (
		_w1129_,
		_w7975_,
		_w7979_,
		_w7980_
	);
	LUT2 #(
		.INIT('h8)
	) name7947 (
		_w7858_,
		_w7980_,
		_w7981_
	);
	LUT3 #(
		.INIT('h80)
	) name7948 (
		_w1437_,
		_w2126_,
		_w2662_,
		_w7982_
	);
	LUT4 #(
		.INIT('h135f)
	) name7949 (
		_w43_,
		_w65_,
		_w46_,
		_w259_,
		_w7983_
	);
	LUT4 #(
		.INIT('h2000)
	) name7950 (
		_w343_,
		_w473_,
		_w948_,
		_w7983_,
		_w7984_
	);
	LUT4 #(
		.INIT('h8000)
	) name7951 (
		_w283_,
		_w2379_,
		_w2702_,
		_w2703_,
		_w7985_
	);
	LUT3 #(
		.INIT('h80)
	) name7952 (
		_w7982_,
		_w7984_,
		_w7985_,
		_w7986_
	);
	LUT2 #(
		.INIT('h4)
	) name7953 (
		_w250_,
		_w1586_,
		_w7987_
	);
	LUT3 #(
		.INIT('h80)
	) name7954 (
		_w1894_,
		_w1992_,
		_w3585_,
		_w7988_
	);
	LUT4 #(
		.INIT('h8000)
	) name7955 (
		_w1708_,
		_w1710_,
		_w7987_,
		_w7988_,
		_w7989_
	);
	LUT4 #(
		.INIT('h135f)
	) name7956 (
		_w110_,
		_w39_,
		_w43_,
		_w44_,
		_w7990_
	);
	LUT4 #(
		.INIT('h4000)
	) name7957 (
		_w432_,
		_w1513_,
		_w1682_,
		_w7990_,
		_w7991_
	);
	LUT3 #(
		.INIT('h80)
	) name7958 (
		_w7986_,
		_w7989_,
		_w7991_,
		_w7992_
	);
	LUT4 #(
		.INIT('h153f)
	) name7959 (
		_w38_,
		_w122_,
		_w93_,
		_w430_,
		_w7993_
	);
	LUT4 #(
		.INIT('h4000)
	) name7960 (
		_w210_,
		_w627_,
		_w4200_,
		_w7993_,
		_w7994_
	);
	LUT2 #(
		.INIT('h8)
	) name7961 (
		_w3166_,
		_w7994_,
		_w7995_
	);
	LUT4 #(
		.INIT('h1000)
	) name7962 (
		_w40_,
		_w141_,
		_w1472_,
		_w1888_,
		_w7996_
	);
	LUT4 #(
		.INIT('h135f)
	) name7963 (
		_w56_,
		_w47_,
		_w184_,
		_w259_,
		_w7997_
	);
	LUT4 #(
		.INIT('h4000)
	) name7964 (
		_w426_,
		_w7571_,
		_w7572_,
		_w7997_,
		_w7998_
	);
	LUT4 #(
		.INIT('h153f)
	) name7965 (
		_w72_,
		_w43_,
		_w93_,
		_w46_,
		_w7999_
	);
	LUT4 #(
		.INIT('h153f)
	) name7966 (
		_w85_,
		_w65_,
		_w166_,
		_w430_,
		_w8000_
	);
	LUT4 #(
		.INIT('h8000)
	) name7967 (
		_w650_,
		_w1570_,
		_w7999_,
		_w8000_,
		_w8001_
	);
	LUT4 #(
		.INIT('h8000)
	) name7968 (
		_w1720_,
		_w8001_,
		_w7996_,
		_w7998_,
		_w8002_
	);
	LUT4 #(
		.INIT('h8000)
	) name7969 (
		_w1830_,
		_w7276_,
		_w7995_,
		_w8002_,
		_w8003_
	);
	LUT2 #(
		.INIT('h8)
	) name7970 (
		_w7992_,
		_w8003_,
		_w8004_
	);
	LUT4 #(
		.INIT('h54ab)
	) name7971 (
		_w7048_,
		_w7081_,
		_w7082_,
		_w7084_,
		_w8005_
	);
	LUT4 #(
		.INIT('h02a8)
	) name7972 (
		_w376_,
		_w6043_,
		_w6933_,
		_w6934_,
		_w8006_
	);
	LUT4 #(
		.INIT('h007d)
	) name7973 (
		_w2407_,
		_w6935_,
		_w6937_,
		_w8006_,
		_w8007_
	);
	LUT3 #(
		.INIT('h70)
	) name7974 (
		_w2527_,
		_w7044_,
		_w8007_,
		_w8008_
	);
	LUT3 #(
		.INIT('h70)
	) name7975 (
		_w377_,
		_w8005_,
		_w8008_,
		_w8009_
	);
	LUT4 #(
		.INIT('heaa8)
	) name7976 (
		_w7845_,
		_w7981_,
		_w8004_,
		_w8009_,
		_w8010_
	);
	LUT2 #(
		.INIT('h8)
	) name7977 (
		_w7845_,
		_w7971_,
		_w8011_
	);
	LUT2 #(
		.INIT('h6)
	) name7978 (
		_w7845_,
		_w7971_,
		_w8012_
	);
	LUT3 #(
		.INIT('h54)
	) name7979 (
		_w7972_,
		_w8010_,
		_w8011_,
		_w8013_
	);
	LUT3 #(
		.INIT('h69)
	) name7980 (
		_w7845_,
		_w7865_,
		_w7868_,
		_w8014_
	);
	LUT4 #(
		.INIT('h1700)
	) name7981 (
		_w7845_,
		_w7971_,
		_w8010_,
		_w8014_,
		_w8015_
	);
	LUT4 #(
		.INIT('h00e8)
	) name7982 (
		_w7845_,
		_w7971_,
		_w8010_,
		_w8014_,
		_w8016_
	);
	LUT4 #(
		.INIT('h54ab)
	) name7983 (
		_w7972_,
		_w8010_,
		_w8011_,
		_w8014_,
		_w8017_
	);
	LUT4 #(
		.INIT('h54ab)
	) name7984 (
		_w7042_,
		_w7087_,
		_w7088_,
		_w7090_,
		_w8018_
	);
	LUT4 #(
		.INIT('h2228)
	) name7985 (
		_w376_,
		_w5067_,
		_w5282_,
		_w6939_,
		_w8019_
	);
	LUT4 #(
		.INIT('h007d)
	) name7986 (
		_w2407_,
		_w6940_,
		_w6942_,
		_w8019_,
		_w8020_
	);
	LUT3 #(
		.INIT('h70)
	) name7987 (
		_w2527_,
		_w7038_,
		_w8020_,
		_w8021_
	);
	LUT3 #(
		.INIT('h70)
	) name7988 (
		_w377_,
		_w8018_,
		_w8021_,
		_w8022_
	);
	LUT3 #(
		.INIT('h54)
	) name7989 (
		_w8015_,
		_w8016_,
		_w8022_,
		_w8023_
	);
	LUT2 #(
		.INIT('h9)
	) name7990 (
		_w7872_,
		_w7878_,
		_w8024_
	);
	LUT4 #(
		.INIT('h4d00)
	) name7991 (
		_w8013_,
		_w8014_,
		_w8022_,
		_w8024_,
		_w8025_
	);
	LUT4 #(
		.INIT('h00b2)
	) name7992 (
		_w8013_,
		_w8014_,
		_w8022_,
		_w8024_,
		_w8026_
	);
	LUT4 #(
		.INIT('h54ab)
	) name7993 (
		_w8015_,
		_w8016_,
		_w8022_,
		_w8024_,
		_w8027_
	);
	LUT4 #(
		.INIT('h02a8)
	) name7994 (
		_w2550_,
		_w7034_,
		_w7097_,
		_w7098_,
		_w8028_
	);
	LUT4 #(
		.INIT('h2228)
	) name7995 (
		_w2854_,
		_w4099_,
		_w4378_,
		_w6951_,
		_w8029_
	);
	LUT3 #(
		.INIT('h82)
	) name7996 (
		_w2549_,
		_w6947_,
		_w6949_,
		_w8030_
	);
	LUT3 #(
		.INIT('h07)
	) name7997 (
		_w2617_,
		_w7032_,
		_w8030_,
		_w8031_
	);
	LUT2 #(
		.INIT('h4)
	) name7998 (
		_w8029_,
		_w8031_,
		_w8032_
	);
	LUT3 #(
		.INIT('h9a)
	) name7999 (
		\a[29] ,
		_w8028_,
		_w8032_,
		_w8033_
	);
	LUT2 #(
		.INIT('h9)
	) name8000 (
		_w7956_,
		_w7963_,
		_w8034_
	);
	LUT4 #(
		.INIT('h4d00)
	) name8001 (
		_w8023_,
		_w8024_,
		_w8033_,
		_w8034_,
		_w8035_
	);
	LUT4 #(
		.INIT('h9669)
	) name8002 (
		_w7880_,
		_w7881_,
		_w7886_,
		_w7954_,
		_w8036_
	);
	LUT4 #(
		.INIT('h0155)
	) name8003 (
		_w7955_,
		_w7964_,
		_w8035_,
		_w8036_,
		_w8037_
	);
	LUT2 #(
		.INIT('h9)
	) name8004 (
		_w7890_,
		_w7896_,
		_w8038_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8005 (
		_w2875_,
		_w7022_,
		_w7109_,
		_w7110_,
		_w8039_
	);
	LUT4 #(
		.INIT('h2228)
	) name8006 (
		_w2986_,
		_w3409_,
		_w3650_,
		_w6959_,
		_w8040_
	);
	LUT3 #(
		.INIT('h82)
	) name8007 (
		_w2874_,
		_w3706_,
		_w6957_,
		_w8041_
	);
	LUT3 #(
		.INIT('h07)
	) name8008 (
		_w2975_,
		_w7020_,
		_w8041_,
		_w8042_
	);
	LUT2 #(
		.INIT('h4)
	) name8009 (
		_w8040_,
		_w8042_,
		_w8043_
	);
	LUT3 #(
		.INIT('h9a)
	) name8010 (
		\a[26] ,
		_w8039_,
		_w8043_,
		_w8044_
	);
	LUT3 #(
		.INIT('hb2)
	) name8011 (
		_w8037_,
		_w8038_,
		_w8044_,
		_w8045_
	);
	LUT4 #(
		.INIT('h20a2)
	) name8012 (
		_w7950_,
		_w8037_,
		_w8038_,
		_w8044_,
		_w8046_
	);
	LUT4 #(
		.INIT('h4504)
	) name8013 (
		_w7950_,
		_w8037_,
		_w8038_,
		_w8044_,
		_w8047_
	);
	LUT3 #(
		.INIT('h82)
	) name8014 (
		_w37_,
		_w7117_,
		_w7119_,
		_w8048_
	);
	LUT3 #(
		.INIT('h82)
	) name8015 (
		_w3262_,
		_w6967_,
		_w6969_,
		_w8049_
	);
	LUT2 #(
		.INIT('h8)
	) name8016 (
		_w3214_,
		_w7014_,
		_w8050_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8017 (
		_w3249_,
		_w3257_,
		_w6964_,
		_w6966_,
		_w8051_
	);
	LUT2 #(
		.INIT('h1)
	) name8018 (
		_w8050_,
		_w8051_,
		_w8052_
	);
	LUT2 #(
		.INIT('h4)
	) name8019 (
		_w8049_,
		_w8052_,
		_w8053_
	);
	LUT3 #(
		.INIT('h9a)
	) name8020 (
		\a[23] ,
		_w8048_,
		_w8053_,
		_w8054_
	);
	LUT4 #(
		.INIT('h088a)
	) name8021 (
		_w7948_,
		_w7950_,
		_w8045_,
		_w8054_,
		_w8055_
	);
	LUT4 #(
		.INIT('he11e)
	) name8022 (
		_w7831_,
		_w7908_,
		_w7909_,
		_w7915_,
		_w8056_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8023 (
		_w3312_,
		_w7004_,
		_w7127_,
		_w7128_,
		_w8057_
	);
	LUT4 #(
		.INIT('h04c8)
	) name8024 (
		_w2622_,
		_w3654_,
		_w6978_,
		_w6980_,
		_w8058_
	);
	LUT3 #(
		.INIT('h84)
	) name8025 (
		_w2872_,
		_w3311_,
		_w6975_,
		_w8059_
	);
	LUT3 #(
		.INIT('h07)
	) name8026 (
		_w3645_,
		_w7002_,
		_w8059_,
		_w8060_
	);
	LUT2 #(
		.INIT('h4)
	) name8027 (
		_w8058_,
		_w8060_,
		_w8061_
	);
	LUT3 #(
		.INIT('h9a)
	) name8028 (
		\a[20] ,
		_w8057_,
		_w8061_,
		_w8062_
	);
	LUT4 #(
		.INIT('hf110)
	) name8029 (
		_w7947_,
		_w8055_,
		_w8056_,
		_w8062_,
		_w8063_
	);
	LUT3 #(
		.INIT('h82)
	) name8030 (
		_w3710_,
		_w7135_,
		_w7172_,
		_w8064_
	);
	LUT3 #(
		.INIT('h28)
	) name8031 (
		_w3886_,
		_w7136_,
		_w7168_,
		_w8065_
	);
	LUT2 #(
		.INIT('h8)
	) name8032 (
		_w3709_,
		_w6996_,
		_w8066_
	);
	LUT4 #(
		.INIT('h04c8)
	) name8033 (
		_w2411_,
		_w3877_,
		_w6983_,
		_w6993_,
		_w8067_
	);
	LUT2 #(
		.INIT('h1)
	) name8034 (
		_w8066_,
		_w8067_,
		_w8068_
	);
	LUT2 #(
		.INIT('h4)
	) name8035 (
		_w8065_,
		_w8068_,
		_w8069_
	);
	LUT3 #(
		.INIT('h9a)
	) name8036 (
		\a[17] ,
		_w8064_,
		_w8069_,
		_w8070_
	);
	LUT3 #(
		.INIT('hd4)
	) name8037 (
		_w7941_,
		_w8063_,
		_w8070_,
		_w8071_
	);
	LUT4 #(
		.INIT('h0445)
	) name8038 (
		_w7940_,
		_w7941_,
		_w8063_,
		_w8070_,
		_w8072_
	);
	LUT2 #(
		.INIT('h9)
	) name8039 (
		_w7825_,
		_w7924_,
		_w8073_
	);
	LUT4 #(
		.INIT('ha220)
	) name8040 (
		_w7940_,
		_w7941_,
		_w8063_,
		_w8070_,
		_w8074_
	);
	LUT4 #(
		.INIT('h599a)
	) name8041 (
		_w7940_,
		_w7941_,
		_w8063_,
		_w8070_,
		_w8075_
	);
	LUT3 #(
		.INIT('h69)
	) name8042 (
		_w7925_,
		_w7926_,
		_w7931_,
		_w8076_
	);
	LUT4 #(
		.INIT('h0071)
	) name8043 (
		_w7940_,
		_w8071_,
		_w8073_,
		_w8076_,
		_w8077_
	);
	LUT2 #(
		.INIT('h6)
	) name8044 (
		_w8073_,
		_w8075_,
		_w8078_
	);
	LUT4 #(
		.INIT('h028a)
	) name8045 (
		_w4033_,
		_w7136_,
		_w7166_,
		_w7167_,
		_w8079_
	);
	LUT4 #(
		.INIT('h87e1)
	) name8046 (
		\a[11] ,
		\a[12] ,
		\a[13] ,
		\a[14] ,
		_w8080_
	);
	LUT3 #(
		.INIT('h0b)
	) name8047 (
		_w7136_,
		_w7166_,
		_w8080_,
		_w8081_
	);
	LUT2 #(
		.INIT('h1)
	) name8048 (
		_w8079_,
		_w8081_,
		_w8082_
	);
	LUT4 #(
		.INIT('h5700)
	) name8049 (
		_w4034_,
		_w7418_,
		_w7419_,
		_w8082_,
		_w8083_
	);
	LUT2 #(
		.INIT('h6)
	) name8050 (
		\a[14] ,
		_w8083_,
		_w8084_
	);
	LUT4 #(
		.INIT('h6665)
	) name8051 (
		_w7948_,
		_w8046_,
		_w8047_,
		_w8054_,
		_w8085_
	);
	LUT4 #(
		.INIT('h04c8)
	) name8052 (
		_w2983_,
		_w3311_,
		_w6972_,
		_w6974_,
		_w8086_
	);
	LUT4 #(
		.INIT('h007b)
	) name8053 (
		_w2872_,
		_w3645_,
		_w6975_,
		_w8086_,
		_w8087_
	);
	LUT3 #(
		.INIT('h70)
	) name8054 (
		_w3654_,
		_w7002_,
		_w8087_,
		_w8088_
	);
	LUT4 #(
		.INIT('h95aa)
	) name8055 (
		\a[20] ,
		_w3312_,
		_w7426_,
		_w8088_,
		_w8089_
	);
	LUT2 #(
		.INIT('h2)
	) name8056 (
		_w8085_,
		_w8089_,
		_w8090_
	);
	LUT2 #(
		.INIT('h4)
	) name8057 (
		_w8085_,
		_w8089_,
		_w8091_
	);
	LUT2 #(
		.INIT('h9)
	) name8058 (
		_w8085_,
		_w8089_,
		_w8092_
	);
	LUT4 #(
		.INIT('h9a59)
	) name8059 (
		_w7950_,
		_w8037_,
		_w8038_,
		_w8044_,
		_w8093_
	);
	LUT2 #(
		.INIT('h9)
	) name8060 (
		_w8054_,
		_w8093_,
		_w8094_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8061 (
		_w2874_,
		_w3882_,
		_w6954_,
		_w6956_,
		_w8095_
	);
	LUT4 #(
		.INIT('h007d)
	) name8062 (
		_w2975_,
		_w3706_,
		_w6957_,
		_w8095_,
		_w8096_
	);
	LUT3 #(
		.INIT('h70)
	) name8063 (
		_w2986_,
		_w7020_,
		_w8096_,
		_w8097_
	);
	LUT4 #(
		.INIT('h95aa)
	) name8064 (
		\a[26] ,
		_w2875_,
		_w7465_,
		_w8097_,
		_w8098_
	);
	LUT4 #(
		.INIT('h001e)
	) name8065 (
		_w7964_,
		_w8035_,
		_w8036_,
		_w8098_,
		_w8099_
	);
	LUT4 #(
		.INIT('h54ab)
	) name8066 (
		_w8025_,
		_w8026_,
		_w8033_,
		_w8034_,
		_w8100_
	);
	LUT3 #(
		.INIT('h82)
	) name8067 (
		_w2550_,
		_w7099_,
		_w7101_,
		_w8101_
	);
	LUT3 #(
		.INIT('h82)
	) name8068 (
		_w2854_,
		_w4030_,
		_w6952_,
		_w8102_
	);
	LUT2 #(
		.INIT('h8)
	) name8069 (
		_w2549_,
		_w7032_,
		_w8103_
	);
	LUT4 #(
		.INIT('h2228)
	) name8070 (
		_w2617_,
		_w4099_,
		_w4378_,
		_w6951_,
		_w8104_
	);
	LUT2 #(
		.INIT('h1)
	) name8071 (
		_w8103_,
		_w8104_,
		_w8105_
	);
	LUT2 #(
		.INIT('h4)
	) name8072 (
		_w8102_,
		_w8105_,
		_w8106_
	);
	LUT3 #(
		.INIT('h9a)
	) name8073 (
		\a[29] ,
		_w8101_,
		_w8106_,
		_w8107_
	);
	LUT3 #(
		.INIT('h82)
	) name8074 (
		_w2875_,
		_w7105_,
		_w7107_,
		_w8108_
	);
	LUT3 #(
		.INIT('h82)
	) name8075 (
		_w2986_,
		_w3706_,
		_w6957_,
		_w8109_
	);
	LUT2 #(
		.INIT('h8)
	) name8076 (
		_w2874_,
		_w7026_,
		_w8110_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8077 (
		_w2975_,
		_w3882_,
		_w6954_,
		_w6956_,
		_w8111_
	);
	LUT2 #(
		.INIT('h1)
	) name8078 (
		_w8110_,
		_w8111_,
		_w8112_
	);
	LUT2 #(
		.INIT('h4)
	) name8079 (
		_w8109_,
		_w8112_,
		_w8113_
	);
	LUT3 #(
		.INIT('h9a)
	) name8080 (
		\a[26] ,
		_w8108_,
		_w8113_,
		_w8114_
	);
	LUT3 #(
		.INIT('hd4)
	) name8081 (
		_w8100_,
		_w8107_,
		_w8114_,
		_w8115_
	);
	LUT4 #(
		.INIT('he100)
	) name8082 (
		_w7964_,
		_w8035_,
		_w8036_,
		_w8098_,
		_w8116_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name8083 (
		_w7964_,
		_w8035_,
		_w8036_,
		_w8098_,
		_w8117_
	);
	LUT3 #(
		.INIT('h54)
	) name8084 (
		_w8099_,
		_w8115_,
		_w8116_,
		_w8118_
	);
	LUT3 #(
		.INIT('h96)
	) name8085 (
		_w8037_,
		_w8038_,
		_w8044_,
		_w8119_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8086 (
		_w37_,
		_w7016_,
		_w7115_,
		_w7116_,
		_w8120_
	);
	LUT4 #(
		.INIT('h04c8)
	) name8087 (
		_w3257_,
		_w3262_,
		_w6964_,
		_w6966_,
		_w8121_
	);
	LUT3 #(
		.INIT('h82)
	) name8088 (
		_w3214_,
		_w6960_,
		_w6962_,
		_w8122_
	);
	LUT3 #(
		.INIT('h07)
	) name8089 (
		_w3249_,
		_w7014_,
		_w8122_,
		_w8123_
	);
	LUT2 #(
		.INIT('h4)
	) name8090 (
		_w8121_,
		_w8123_,
		_w8124_
	);
	LUT3 #(
		.INIT('h9a)
	) name8091 (
		\a[23] ,
		_w8120_,
		_w8124_,
		_w8125_
	);
	LUT3 #(
		.INIT('hb2)
	) name8092 (
		_w8118_,
		_w8119_,
		_w8125_,
		_w8126_
	);
	LUT3 #(
		.INIT('h82)
	) name8093 (
		_w3312_,
		_w7123_,
		_w7125_,
		_w8127_
	);
	LUT3 #(
		.INIT('h84)
	) name8094 (
		_w2872_,
		_w3654_,
		_w6975_,
		_w8128_
	);
	LUT2 #(
		.INIT('h8)
	) name8095 (
		_w3311_,
		_w7008_,
		_w8129_
	);
	LUT4 #(
		.INIT('h04c8)
	) name8096 (
		_w2983_,
		_w3645_,
		_w6972_,
		_w6974_,
		_w8130_
	);
	LUT2 #(
		.INIT('h1)
	) name8097 (
		_w8129_,
		_w8130_,
		_w8131_
	);
	LUT2 #(
		.INIT('h4)
	) name8098 (
		_w8128_,
		_w8131_,
		_w8132_
	);
	LUT3 #(
		.INIT('h9a)
	) name8099 (
		\a[20] ,
		_w8127_,
		_w8132_,
		_w8133_
	);
	LUT3 #(
		.INIT('hd4)
	) name8100 (
		_w8094_,
		_w8126_,
		_w8133_,
		_w8134_
	);
	LUT3 #(
		.INIT('h54)
	) name8101 (
		_w8090_,
		_w8091_,
		_w8134_,
		_w8135_
	);
	LUT4 #(
		.INIT('he11e)
	) name8102 (
		_w7947_,
		_w8055_,
		_w8056_,
		_w8062_,
		_w8136_
	);
	LUT4 #(
		.INIT('h2b00)
	) name8103 (
		_w8085_,
		_w8089_,
		_w8134_,
		_w8136_,
		_w8137_
	);
	LUT4 #(
		.INIT('h00d4)
	) name8104 (
		_w8085_,
		_w8089_,
		_w8134_,
		_w8136_,
		_w8138_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8105 (
		_w3710_,
		_w6998_,
		_w7133_,
		_w7134_,
		_w8139_
	);
	LUT4 #(
		.INIT('h04c8)
	) name8106 (
		_w2411_,
		_w3886_,
		_w6983_,
		_w6993_,
		_w8140_
	);
	LUT3 #(
		.INIT('h84)
	) name8107 (
		_w2546_,
		_w3709_,
		_w6981_,
		_w8141_
	);
	LUT3 #(
		.INIT('h07)
	) name8108 (
		_w3877_,
		_w6996_,
		_w8141_,
		_w8142_
	);
	LUT2 #(
		.INIT('h4)
	) name8109 (
		_w8140_,
		_w8142_,
		_w8143_
	);
	LUT3 #(
		.INIT('h9a)
	) name8110 (
		\a[17] ,
		_w8139_,
		_w8143_,
		_w8144_
	);
	LUT3 #(
		.INIT('h54)
	) name8111 (
		_w8137_,
		_w8138_,
		_w8144_,
		_w8145_
	);
	LUT4 #(
		.INIT('h1051)
	) name8112 (
		_w8084_,
		_w8135_,
		_w8136_,
		_w8144_,
		_w8146_
	);
	LUT4 #(
		.INIT('h8a08)
	) name8113 (
		_w8084_,
		_w8135_,
		_w8136_,
		_w8144_,
		_w8147_
	);
	LUT3 #(
		.INIT('h96)
	) name8114 (
		_w7941_,
		_w8063_,
		_w8070_,
		_w8148_
	);
	LUT3 #(
		.INIT('h45)
	) name8115 (
		_w8146_,
		_w8147_,
		_w8148_,
		_w8149_
	);
	LUT4 #(
		.INIT('h2a02)
	) name8116 (
		_w8078_,
		_w8084_,
		_w8145_,
		_w8148_,
		_w8150_
	);
	LUT4 #(
		.INIT('h999a)
	) name8117 (
		_w8084_,
		_w8137_,
		_w8138_,
		_w8144_,
		_w8151_
	);
	LUT2 #(
		.INIT('h6)
	) name8118 (
		_w8148_,
		_w8151_,
		_w8152_
	);
	LUT4 #(
		.INIT('h04c8)
	) name8119 (
		_w2622_,
		_w3709_,
		_w6978_,
		_w6980_,
		_w8153_
	);
	LUT4 #(
		.INIT('h007b)
	) name8120 (
		_w2546_,
		_w3877_,
		_w6981_,
		_w8153_,
		_w8154_
	);
	LUT3 #(
		.INIT('h70)
	) name8121 (
		_w3886_,
		_w6996_,
		_w8154_,
		_w8155_
	);
	LUT4 #(
		.INIT('h95aa)
	) name8122 (
		\a[17] ,
		_w3710_,
		_w7500_,
		_w8155_,
		_w8156_
	);
	LUT3 #(
		.INIT('h09)
	) name8123 (
		_w8092_,
		_w8134_,
		_w8156_,
		_w8157_
	);
	LUT3 #(
		.INIT('h60)
	) name8124 (
		_w8092_,
		_w8134_,
		_w8156_,
		_w8158_
	);
	LUT3 #(
		.INIT('h96)
	) name8125 (
		_w8092_,
		_w8134_,
		_w8156_,
		_w8159_
	);
	LUT3 #(
		.INIT('h96)
	) name8126 (
		_w8094_,
		_w8126_,
		_w8133_,
		_w8160_
	);
	LUT4 #(
		.INIT('h2228)
	) name8127 (
		_w3214_,
		_w3409_,
		_w3650_,
		_w6959_,
		_w8161_
	);
	LUT4 #(
		.INIT('h007d)
	) name8128 (
		_w3249_,
		_w6960_,
		_w6962_,
		_w8161_,
		_w8162_
	);
	LUT3 #(
		.INIT('h70)
	) name8129 (
		_w3262_,
		_w7014_,
		_w8162_,
		_w8163_
	);
	LUT4 #(
		.INIT('h95aa)
	) name8130 (
		\a[23] ,
		_w37_,
		_w7291_,
		_w8163_,
		_w8164_
	);
	LUT3 #(
		.INIT('h09)
	) name8131 (
		_w8115_,
		_w8117_,
		_w8164_,
		_w8165_
	);
	LUT3 #(
		.INIT('h60)
	) name8132 (
		_w8115_,
		_w8117_,
		_w8164_,
		_w8166_
	);
	LUT3 #(
		.INIT('h96)
	) name8133 (
		_w8115_,
		_w8117_,
		_w8164_,
		_w8167_
	);
	LUT3 #(
		.INIT('h96)
	) name8134 (
		_w8100_,
		_w8107_,
		_w8114_,
		_w8168_
	);
	LUT2 #(
		.INIT('h9)
	) name8135 (
		_w8027_,
		_w8033_,
		_w8169_
	);
	LUT3 #(
		.INIT('h82)
	) name8136 (
		_w377_,
		_w7087_,
		_w7089_,
		_w8170_
	);
	LUT3 #(
		.INIT('h82)
	) name8137 (
		_w2527_,
		_w6940_,
		_w6942_,
		_w8171_
	);
	LUT2 #(
		.INIT('h8)
	) name8138 (
		_w376_,
		_w7044_,
		_w8172_
	);
	LUT4 #(
		.INIT('h2228)
	) name8139 (
		_w2407_,
		_w5067_,
		_w5282_,
		_w6939_,
		_w8173_
	);
	LUT2 #(
		.INIT('h1)
	) name8140 (
		_w8172_,
		_w8173_,
		_w8174_
	);
	LUT2 #(
		.INIT('h4)
	) name8141 (
		_w8171_,
		_w8174_,
		_w8175_
	);
	LUT2 #(
		.INIT('h4)
	) name8142 (
		_w8170_,
		_w8175_,
		_w8176_
	);
	LUT3 #(
		.INIT('h09)
	) name8143 (
		_w8010_,
		_w8012_,
		_w8176_,
		_w8177_
	);
	LUT4 #(
		.INIT('h6339)
	) name8144 (
		_w7845_,
		_w7981_,
		_w8004_,
		_w8009_,
		_w8178_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8145 (
		_w377_,
		_w7046_,
		_w7085_,
		_w7086_,
		_w8179_
	);
	LUT4 #(
		.INIT('h2228)
	) name8146 (
		_w2527_,
		_w5067_,
		_w5282_,
		_w6939_,
		_w8180_
	);
	LUT3 #(
		.INIT('h82)
	) name8147 (
		_w376_,
		_w6935_,
		_w6937_,
		_w8181_
	);
	LUT3 #(
		.INIT('h07)
	) name8148 (
		_w2407_,
		_w7044_,
		_w8181_,
		_w8182_
	);
	LUT2 #(
		.INIT('h4)
	) name8149 (
		_w8180_,
		_w8182_,
		_w8183_
	);
	LUT2 #(
		.INIT('h4)
	) name8150 (
		_w8179_,
		_w8183_,
		_w8184_
	);
	LUT2 #(
		.INIT('h2)
	) name8151 (
		_w8178_,
		_w8184_,
		_w8185_
	);
	LUT4 #(
		.INIT('h8000)
	) name8152 (
		_w817_,
		_w889_,
		_w857_,
		_w2257_,
		_w8186_
	);
	LUT3 #(
		.INIT('h80)
	) name8153 (
		_w1987_,
		_w7517_,
		_w8186_,
		_w8187_
	);
	LUT4 #(
		.INIT('h135f)
	) name8154 (
		_w106_,
		_w67_,
		_w90_,
		_w158_,
		_w8188_
	);
	LUT3 #(
		.INIT('h20)
	) name8155 (
		_w277_,
		_w396_,
		_w8188_,
		_w8189_
	);
	LUT2 #(
		.INIT('h8)
	) name8156 (
		_w2590_,
		_w8189_,
		_w8190_
	);
	LUT4 #(
		.INIT('h153f)
	) name8157 (
		_w59_,
		_w43_,
		_w44_,
		_w184_,
		_w8191_
	);
	LUT4 #(
		.INIT('h4000)
	) name8158 (
		_w346_,
		_w820_,
		_w2219_,
		_w8191_,
		_w8192_
	);
	LUT4 #(
		.INIT('h8000)
	) name8159 (
		_w302_,
		_w403_,
		_w663_,
		_w839_,
		_w8193_
	);
	LUT4 #(
		.INIT('h8000)
	) name8160 (
		_w2590_,
		_w8189_,
		_w8192_,
		_w8193_,
		_w8194_
	);
	LUT4 #(
		.INIT('h8000)
	) name8161 (
		_w1057_,
		_w1070_,
		_w8187_,
		_w8194_,
		_w8195_
	);
	LUT2 #(
		.INIT('h8)
	) name8162 (
		_w3357_,
		_w8195_,
		_w8196_
	);
	LUT3 #(
		.INIT('h82)
	) name8163 (
		_w377_,
		_w7081_,
		_w7083_,
		_w8197_
	);
	LUT3 #(
		.INIT('h82)
	) name8164 (
		_w2527_,
		_w6935_,
		_w6937_,
		_w8198_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8165 (
		_w2407_,
		_w6043_,
		_w6933_,
		_w6934_,
		_w8199_
	);
	LUT2 #(
		.INIT('h8)
	) name8166 (
		_w376_,
		_w7050_,
		_w8200_
	);
	LUT2 #(
		.INIT('h1)
	) name8167 (
		_w8199_,
		_w8200_,
		_w8201_
	);
	LUT2 #(
		.INIT('h4)
	) name8168 (
		_w8198_,
		_w8201_,
		_w8202_
	);
	LUT3 #(
		.INIT('h45)
	) name8169 (
		_w8196_,
		_w8197_,
		_w8202_,
		_w8203_
	);
	LUT4 #(
		.INIT('h153f)
	) name8170 (
		_w67_,
		_w44_,
		_w166_,
		_w259_,
		_w8204_
	);
	LUT4 #(
		.INIT('h135f)
	) name8171 (
		_w106_,
		_w52_,
		_w44_,
		_w430_,
		_w8205_
	);
	LUT2 #(
		.INIT('h8)
	) name8172 (
		_w8204_,
		_w8205_,
		_w8206_
	);
	LUT4 #(
		.INIT('h0777)
	) name8173 (
		_w122_,
		_w85_,
		_w41_,
		_w72_,
		_w8207_
	);
	LUT4 #(
		.INIT('h8000)
	) name8174 (
		_w370_,
		_w976_,
		_w1341_,
		_w8207_,
		_w8208_
	);
	LUT3 #(
		.INIT('h80)
	) name8175 (
		_w2258_,
		_w2281_,
		_w2744_,
		_w8209_
	);
	LUT4 #(
		.INIT('h8000)
	) name8176 (
		_w2070_,
		_w8206_,
		_w8209_,
		_w8208_,
		_w8210_
	);
	LUT4 #(
		.INIT('h8000)
	) name8177 (
		_w2441_,
		_w2444_,
		_w3923_,
		_w3924_,
		_w8211_
	);
	LUT4 #(
		.INIT('h8000)
	) name8178 (
		_w1018_,
		_w1025_,
		_w8210_,
		_w8211_,
		_w8212_
	);
	LUT2 #(
		.INIT('h8)
	) name8179 (
		_w1272_,
		_w8212_,
		_w8213_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8180 (
		_w377_,
		_w7052_,
		_w7079_,
		_w7080_,
		_w8214_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8181 (
		_w2527_,
		_w6043_,
		_w6933_,
		_w6934_,
		_w8215_
	);
	LUT3 #(
		.INIT('h82)
	) name8182 (
		_w376_,
		_w6929_,
		_w6931_,
		_w8216_
	);
	LUT3 #(
		.INIT('h07)
	) name8183 (
		_w2407_,
		_w7050_,
		_w8216_,
		_w8217_
	);
	LUT2 #(
		.INIT('h4)
	) name8184 (
		_w8215_,
		_w8217_,
		_w8218_
	);
	LUT3 #(
		.INIT('h45)
	) name8185 (
		_w8213_,
		_w8214_,
		_w8218_,
		_w8219_
	);
	LUT4 #(
		.INIT('h1000)
	) name8186 (
		_w237_,
		_w362_,
		_w1589_,
		_w2173_,
		_w8220_
	);
	LUT4 #(
		.INIT('h8000)
	) name8187 (
		_w108_,
		_w1222_,
		_w1278_,
		_w1625_,
		_w8221_
	);
	LUT4 #(
		.INIT('h153f)
	) name8188 (
		_w85_,
		_w44_,
		_w176_,
		_w378_,
		_w8222_
	);
	LUT4 #(
		.INIT('h0800)
	) name8189 (
		_w219_,
		_w222_,
		_w424_,
		_w8222_,
		_w8223_
	);
	LUT4 #(
		.INIT('h8000)
	) name8190 (
		_w3110_,
		_w8221_,
		_w8223_,
		_w8220_,
		_w8224_
	);
	LUT4 #(
		.INIT('h8000)
	) name8191 (
		_w1699_,
		_w1706_,
		_w2142_,
		_w8224_,
		_w8225_
	);
	LUT2 #(
		.INIT('h8)
	) name8192 (
		_w7992_,
		_w8225_,
		_w8226_
	);
	LUT4 #(
		.INIT('h54ab)
	) name8193 (
		_w7054_,
		_w7075_,
		_w7076_,
		_w7078_,
		_w8227_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8194 (
		_w376_,
		_w6645_,
		_w6926_,
		_w6928_,
		_w8228_
	);
	LUT4 #(
		.INIT('h007d)
	) name8195 (
		_w2407_,
		_w6929_,
		_w6931_,
		_w8228_,
		_w8229_
	);
	LUT3 #(
		.INIT('h70)
	) name8196 (
		_w2527_,
		_w7050_,
		_w8229_,
		_w8230_
	);
	LUT4 #(
		.INIT('h2033)
	) name8197 (
		_w377_,
		_w8226_,
		_w8227_,
		_w8230_,
		_w8231_
	);
	LUT4 #(
		.INIT('h0777)
	) name8198 (
		_w122_,
		_w85_,
		_w41_,
		_w184_,
		_w8232_
	);
	LUT4 #(
		.INIT('h135f)
	) name8199 (
		_w38_,
		_w110_,
		_w236_,
		_w166_,
		_w8233_
	);
	LUT4 #(
		.INIT('h8000)
	) name8200 (
		_w216_,
		_w842_,
		_w8232_,
		_w8233_,
		_w8234_
	);
	LUT3 #(
		.INIT('h40)
	) name8201 (
		_w362_,
		_w1589_,
		_w2432_,
		_w8235_
	);
	LUT4 #(
		.INIT('h153f)
	) name8202 (
		_w38_,
		_w43_,
		_w65_,
		_w166_,
		_w8236_
	);
	LUT4 #(
		.INIT('h135f)
	) name8203 (
		_w52_,
		_w46_,
		_w176_,
		_w430_,
		_w8237_
	);
	LUT4 #(
		.INIT('h8000)
	) name8204 (
		_w54_,
		_w1216_,
		_w8236_,
		_w8237_,
		_w8238_
	);
	LUT3 #(
		.INIT('h80)
	) name8205 (
		_w790_,
		_w1414_,
		_w3135_,
		_w8239_
	);
	LUT4 #(
		.INIT('h8000)
	) name8206 (
		_w8238_,
		_w8239_,
		_w8234_,
		_w8235_,
		_w8240_
	);
	LUT4 #(
		.INIT('h8000)
	) name8207 (
		_w500_,
		_w658_,
		_w2827_,
		_w2831_,
		_w8241_
	);
	LUT2 #(
		.INIT('h8)
	) name8208 (
		_w8240_,
		_w8241_,
		_w8242_
	);
	LUT2 #(
		.INIT('h8)
	) name8209 (
		_w2687_,
		_w8242_,
		_w8243_
	);
	LUT3 #(
		.INIT('h82)
	) name8210 (
		_w377_,
		_w7075_,
		_w7077_,
		_w8244_
	);
	LUT3 #(
		.INIT('h82)
	) name8211 (
		_w2527_,
		_w6929_,
		_w6931_,
		_w8245_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8212 (
		_w2407_,
		_w6645_,
		_w6926_,
		_w6928_,
		_w8246_
	);
	LUT2 #(
		.INIT('h8)
	) name8213 (
		_w376_,
		_w7056_,
		_w8247_
	);
	LUT2 #(
		.INIT('h1)
	) name8214 (
		_w8246_,
		_w8247_,
		_w8248_
	);
	LUT2 #(
		.INIT('h4)
	) name8215 (
		_w8245_,
		_w8248_,
		_w8249_
	);
	LUT2 #(
		.INIT('h4)
	) name8216 (
		_w8244_,
		_w8249_,
		_w8250_
	);
	LUT3 #(
		.INIT('h45)
	) name8217 (
		_w8243_,
		_w8244_,
		_w8249_,
		_w8251_
	);
	LUT3 #(
		.INIT('h40)
	) name8218 (
		_w315_,
		_w2432_,
		_w3346_,
		_w8252_
	);
	LUT2 #(
		.INIT('h8)
	) name8219 (
		_w361_,
		_w611_,
		_w8253_
	);
	LUT4 #(
		.INIT('h8000)
	) name8220 (
		_w370_,
		_w361_,
		_w611_,
		_w7596_,
		_w8254_
	);
	LUT2 #(
		.INIT('h8)
	) name8221 (
		_w8252_,
		_w8254_,
		_w8255_
	);
	LUT3 #(
		.INIT('h80)
	) name8222 (
		_w806_,
		_w1992_,
		_w7326_,
		_w8256_
	);
	LUT3 #(
		.INIT('h37)
	) name8223 (
		_w90_,
		_w72_,
		_w50_,
		_w8257_
	);
	LUT4 #(
		.INIT('h8000)
	) name8224 (
		_w96_,
		_w245_,
		_w248_,
		_w8257_,
		_w8258_
	);
	LUT3 #(
		.INIT('h80)
	) name8225 (
		_w229_,
		_w8256_,
		_w8258_,
		_w8259_
	);
	LUT2 #(
		.INIT('h8)
	) name8226 (
		_w8255_,
		_w8259_,
		_w8260_
	);
	LUT4 #(
		.INIT('h153f)
	) name8227 (
		_w47_,
		_w41_,
		_w201_,
		_w158_,
		_w8261_
	);
	LUT4 #(
		.INIT('h4000)
	) name8228 (
		_w425_,
		_w902_,
		_w1502_,
		_w8261_,
		_w8262_
	);
	LUT4 #(
		.INIT('h135f)
	) name8229 (
		_w85_,
		_w110_,
		_w158_,
		_w176_,
		_w8263_
	);
	LUT4 #(
		.INIT('h4000)
	) name8230 (
		_w338_,
		_w1575_,
		_w3022_,
		_w8263_,
		_w8264_
	);
	LUT4 #(
		.INIT('h0777)
	) name8231 (
		_w106_,
		_w47_,
		_w39_,
		_w93_,
		_w8265_
	);
	LUT3 #(
		.INIT('h80)
	) name8232 (
		_w1091_,
		_w2825_,
		_w8265_,
		_w8266_
	);
	LUT4 #(
		.INIT('h8000)
	) name8233 (
		_w2808_,
		_w8266_,
		_w8262_,
		_w8264_,
		_w8267_
	);
	LUT2 #(
		.INIT('h8)
	) name8234 (
		_w4193_,
		_w8267_,
		_w8268_
	);
	LUT3 #(
		.INIT('h80)
	) name8235 (
		_w1360_,
		_w1837_,
		_w7265_,
		_w8269_
	);
	LUT4 #(
		.INIT('h153f)
	) name8236 (
		_w110_,
		_w41_,
		_w39_,
		_w43_,
		_w8270_
	);
	LUT4 #(
		.INIT('h153f)
	) name8237 (
		_w52_,
		_w110_,
		_w419_,
		_w378_,
		_w8271_
	);
	LUT4 #(
		.INIT('h8000)
	) name8238 (
		_w54_,
		_w292_,
		_w8270_,
		_w8271_,
		_w8272_
	);
	LUT4 #(
		.INIT('h8000)
	) name8239 (
		_w188_,
		_w4137_,
		_w8269_,
		_w8272_,
		_w8273_
	);
	LUT2 #(
		.INIT('h8)
	) name8240 (
		_w2477_,
		_w4172_,
		_w8274_
	);
	LUT4 #(
		.INIT('h8000)
	) name8241 (
		_w68_,
		_w1158_,
		_w1411_,
		_w2237_,
		_w8275_
	);
	LUT4 #(
		.INIT('h8000)
	) name8242 (
		_w7450_,
		_w7452_,
		_w8274_,
		_w8275_,
		_w8276_
	);
	LUT4 #(
		.INIT('h8000)
	) name8243 (
		_w4193_,
		_w8267_,
		_w8273_,
		_w8276_,
		_w8277_
	);
	LUT2 #(
		.INIT('h8)
	) name8244 (
		_w8260_,
		_w8277_,
		_w8278_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8245 (
		_w377_,
		_w7058_,
		_w7073_,
		_w7074_,
		_w8279_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8246 (
		_w2527_,
		_w6645_,
		_w6926_,
		_w6928_,
		_w8280_
	);
	LUT3 #(
		.INIT('h82)
	) name8247 (
		_w376_,
		_w6922_,
		_w6924_,
		_w8281_
	);
	LUT3 #(
		.INIT('h07)
	) name8248 (
		_w2407_,
		_w7056_,
		_w8281_,
		_w8282_
	);
	LUT2 #(
		.INIT('h4)
	) name8249 (
		_w8280_,
		_w8282_,
		_w8283_
	);
	LUT3 #(
		.INIT('h45)
	) name8250 (
		_w8278_,
		_w8279_,
		_w8283_,
		_w8284_
	);
	LUT4 #(
		.INIT('h4000)
	) name8251 (
		_w392_,
		_w908_,
		_w1084_,
		_w2489_,
		_w8285_
	);
	LUT3 #(
		.INIT('h80)
	) name8252 (
		_w1761_,
		_w2125_,
		_w7141_,
		_w8286_
	);
	LUT4 #(
		.INIT('h135f)
	) name8253 (
		_w90_,
		_w93_,
		_w201_,
		_w176_,
		_w8287_
	);
	LUT4 #(
		.INIT('h135f)
	) name8254 (
		_w122_,
		_w90_,
		_w56_,
		_w378_,
		_w8288_
	);
	LUT4 #(
		.INIT('h8000)
	) name8255 (
		_w675_,
		_w1334_,
		_w8287_,
		_w8288_,
		_w8289_
	);
	LUT4 #(
		.INIT('h8000)
	) name8256 (
		_w2585_,
		_w8286_,
		_w8289_,
		_w8285_,
		_w8290_
	);
	LUT3 #(
		.INIT('h80)
	) name8257 (
		_w1407_,
		_w7617_,
		_w8290_,
		_w8291_
	);
	LUT4 #(
		.INIT('h8000)
	) name8258 (
		_w1438_,
		_w1921_,
		_w2086_,
		_w2472_,
		_w8292_
	);
	LUT4 #(
		.INIT('h0777)
	) name8259 (
		_w122_,
		_w110_,
		_w90_,
		_w236_,
		_w8293_
	);
	LUT4 #(
		.INIT('h2000)
	) name8260 (
		_w305_,
		_w458_,
		_w793_,
		_w8293_,
		_w8294_
	);
	LUT3 #(
		.INIT('h80)
	) name8261 (
		_w1747_,
		_w8292_,
		_w8294_,
		_w8295_
	);
	LUT3 #(
		.INIT('h80)
	) name8262 (
		_w2572_,
		_w7154_,
		_w8295_,
		_w8296_
	);
	LUT2 #(
		.INIT('h8)
	) name8263 (
		_w8291_,
		_w8296_,
		_w8297_
	);
	LUT4 #(
		.INIT('h54ab)
	) name8264 (
		_w7060_,
		_w7069_,
		_w7070_,
		_w7072_,
		_w8298_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8265 (
		_w376_,
		_w6669_,
		_w6919_,
		_w6921_,
		_w8299_
	);
	LUT4 #(
		.INIT('h007d)
	) name8266 (
		_w2407_,
		_w6922_,
		_w6924_,
		_w8299_,
		_w8300_
	);
	LUT3 #(
		.INIT('h70)
	) name8267 (
		_w2527_,
		_w7056_,
		_w8300_,
		_w8301_
	);
	LUT4 #(
		.INIT('h2033)
	) name8268 (
		_w377_,
		_w8297_,
		_w8298_,
		_w8301_,
		_w8302_
	);
	LUT4 #(
		.INIT('h135f)
	) name8269 (
		_w50_,
		_w93_,
		_w236_,
		_w158_,
		_w8303_
	);
	LUT4 #(
		.INIT('h153f)
	) name8270 (
		_w38_,
		_w78_,
		_w47_,
		_w430_,
		_w8304_
	);
	LUT4 #(
		.INIT('h8000)
	) name8271 (
		_w115_,
		_w116_,
		_w8303_,
		_w8304_,
		_w8305_
	);
	LUT3 #(
		.INIT('h40)
	) name8272 (
		_w276_,
		_w1153_,
		_w7220_,
		_w8306_
	);
	LUT4 #(
		.INIT('h0777)
	) name8273 (
		_w106_,
		_w55_,
		_w43_,
		_w46_,
		_w8307_
	);
	LUT4 #(
		.INIT('h153f)
	) name8274 (
		_w38_,
		_w85_,
		_w78_,
		_w201_,
		_w8308_
	);
	LUT3 #(
		.INIT('h80)
	) name8275 (
		_w909_,
		_w8307_,
		_w8308_,
		_w8309_
	);
	LUT4 #(
		.INIT('h8000)
	) name8276 (
		_w2087_,
		_w8306_,
		_w8309_,
		_w8305_,
		_w8310_
	);
	LUT4 #(
		.INIT('h153f)
	) name8277 (
		_w52_,
		_w67_,
		_w236_,
		_w259_,
		_w8311_
	);
	LUT3 #(
		.INIT('h40)
	) name8278 (
		_w432_,
		_w2809_,
		_w8311_,
		_w8312_
	);
	LUT4 #(
		.INIT('h8000)
	) name8279 (
		_w640_,
		_w7580_,
		_w7581_,
		_w8312_,
		_w8313_
	);
	LUT2 #(
		.INIT('h8)
	) name8280 (
		_w8310_,
		_w8313_,
		_w8314_
	);
	LUT4 #(
		.INIT('h135f)
	) name8281 (
		_w59_,
		_w67_,
		_w259_,
		_w378_,
		_w8315_
	);
	LUT4 #(
		.INIT('h153f)
	) name8282 (
		_w110_,
		_w78_,
		_w50_,
		_w201_,
		_w8316_
	);
	LUT4 #(
		.INIT('h2000)
	) name8283 (
		_w262_,
		_w424_,
		_w8316_,
		_w8315_,
		_w8317_
	);
	LUT2 #(
		.INIT('h8)
	) name8284 (
		_w1357_,
		_w8317_,
		_w8318_
	);
	LUT3 #(
		.INIT('h80)
	) name8285 (
		_w1403_,
		_w1673_,
		_w1978_,
		_w8319_
	);
	LUT3 #(
		.INIT('h80)
	) name8286 (
		_w1002_,
		_w3322_,
		_w8319_,
		_w8320_
	);
	LUT3 #(
		.INIT('h80)
	) name8287 (
		_w2007_,
		_w8318_,
		_w8320_,
		_w8321_
	);
	LUT3 #(
		.INIT('h80)
	) name8288 (
		_w1584_,
		_w8314_,
		_w8321_,
		_w8322_
	);
	LUT3 #(
		.INIT('h82)
	) name8289 (
		_w377_,
		_w7069_,
		_w7071_,
		_w8323_
	);
	LUT3 #(
		.INIT('h82)
	) name8290 (
		_w2527_,
		_w6922_,
		_w6924_,
		_w8324_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8291 (
		_w2407_,
		_w6669_,
		_w6919_,
		_w6921_,
		_w8325_
	);
	LUT2 #(
		.INIT('h8)
	) name8292 (
		_w376_,
		_w7062_,
		_w8326_
	);
	LUT2 #(
		.INIT('h1)
	) name8293 (
		_w8325_,
		_w8326_,
		_w8327_
	);
	LUT2 #(
		.INIT('h4)
	) name8294 (
		_w8324_,
		_w8327_,
		_w8328_
	);
	LUT3 #(
		.INIT('h80)
	) name8295 (
		_w460_,
		_w2195_,
		_w4159_,
		_w8329_
	);
	LUT3 #(
		.INIT('h80)
	) name8296 (
		_w1089_,
		_w1910_,
		_w2823_,
		_w8330_
	);
	LUT4 #(
		.INIT('h135f)
	) name8297 (
		_w67_,
		_w56_,
		_w259_,
		_w176_,
		_w8331_
	);
	LUT4 #(
		.INIT('h0800)
	) name8298 (
		_w216_,
		_w316_,
		_w426_,
		_w8331_,
		_w8332_
	);
	LUT4 #(
		.INIT('h8000)
	) name8299 (
		_w3584_,
		_w3586_,
		_w8330_,
		_w8332_,
		_w8333_
	);
	LUT4 #(
		.INIT('h8000)
	) name8300 (
		_w2387_,
		_w2430_,
		_w8329_,
		_w8333_,
		_w8334_
	);
	LUT2 #(
		.INIT('h8)
	) name8301 (
		_w2800_,
		_w8334_,
		_w8335_
	);
	LUT3 #(
		.INIT('h28)
	) name8302 (
		_w377_,
		_w7065_,
		_w7068_,
		_w8336_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8303 (
		_w2527_,
		_w6669_,
		_w6919_,
		_w6921_,
		_w8337_
	);
	LUT3 #(
		.INIT('h82)
	) name8304 (
		_w376_,
		_w6914_,
		_w6916_,
		_w8338_
	);
	LUT3 #(
		.INIT('h07)
	) name8305 (
		_w2407_,
		_w7062_,
		_w8338_,
		_w8339_
	);
	LUT2 #(
		.INIT('h4)
	) name8306 (
		_w8337_,
		_w8339_,
		_w8340_
	);
	LUT3 #(
		.INIT('h80)
	) name8307 (
		_w529_,
		_w2515_,
		_w8238_,
		_w8341_
	);
	LUT4 #(
		.INIT('h135f)
	) name8308 (
		_w41_,
		_w93_,
		_w201_,
		_w236_,
		_w8342_
	);
	LUT4 #(
		.INIT('h0777)
	) name8309 (
		_w55_,
		_w39_,
		_w50_,
		_w184_,
		_w8343_
	);
	LUT4 #(
		.INIT('h4000)
	) name8310 (
		_w369_,
		_w1975_,
		_w8343_,
		_w8342_,
		_w8344_
	);
	LUT4 #(
		.INIT('h8000)
	) name8311 (
		_w115_,
		_w662_,
		_w713_,
		_w731_,
		_w8345_
	);
	LUT4 #(
		.INIT('h0777)
	) name8312 (
		_w106_,
		_w59_,
		_w56_,
		_w184_,
		_w8346_
	);
	LUT4 #(
		.INIT('h0777)
	) name8313 (
		_w106_,
		_w56_,
		_w46_,
		_w158_,
		_w8347_
	);
	LUT4 #(
		.INIT('h4000)
	) name8314 (
		_w476_,
		_w479_,
		_w8346_,
		_w8347_,
		_w8348_
	);
	LUT4 #(
		.INIT('h8000)
	) name8315 (
		_w1317_,
		_w8344_,
		_w8345_,
		_w8348_,
		_w8349_
	);
	LUT2 #(
		.INIT('h8)
	) name8316 (
		_w8341_,
		_w8349_,
		_w8350_
	);
	LUT2 #(
		.INIT('h2)
	) name8317 (
		_w343_,
		_w469_,
		_w8351_
	);
	LUT4 #(
		.INIT('h135f)
	) name8318 (
		_w52_,
		_w47_,
		_w39_,
		_w184_,
		_w8352_
	);
	LUT4 #(
		.INIT('h8000)
	) name8319 (
		_w1238_,
		_w1529_,
		_w1651_,
		_w8352_,
		_w8353_
	);
	LUT2 #(
		.INIT('h8)
	) name8320 (
		_w8351_,
		_w8353_,
		_w8354_
	);
	LUT4 #(
		.INIT('h8000)
	) name8321 (
		_w603_,
		_w1899_,
		_w1923_,
		_w1940_,
		_w8355_
	);
	LUT3 #(
		.INIT('h80)
	) name8322 (
		_w4221_,
		_w8354_,
		_w8355_,
		_w8356_
	);
	LUT3 #(
		.INIT('h80)
	) name8323 (
		_w2076_,
		_w8350_,
		_w8356_,
		_w8357_
	);
	LUT3 #(
		.INIT('h09)
	) name8324 (
		_w6914_,
		_w6916_,
		_w7067_,
		_w8358_
	);
	LUT4 #(
		.INIT('h2882)
	) name8325 (
		_w377_,
		_w6914_,
		_w6916_,
		_w7067_,
		_w8359_
	);
	LUT4 #(
		.INIT('ha802)
	) name8326 (
		_w2407_,
		_w6689_,
		_w6911_,
		_w6913_,
		_w8360_
	);
	LUT4 #(
		.INIT('h007d)
	) name8327 (
		_w2527_,
		_w6914_,
		_w6916_,
		_w8360_,
		_w8361_
	);
	LUT3 #(
		.INIT('h37)
	) name8328 (
		_w72_,
		_w46_,
		_w166_,
		_w8362_
	);
	LUT4 #(
		.INIT('h8000)
	) name8329 (
		_w143_,
		_w1297_,
		_w1529_,
		_w8362_,
		_w8363_
	);
	LUT3 #(
		.INIT('h37)
	) name8330 (
		_w106_,
		_w44_,
		_w259_,
		_w8364_
	);
	LUT4 #(
		.INIT('h4000)
	) name8331 (
		_w482_,
		_w1147_,
		_w1148_,
		_w8364_,
		_w8365_
	);
	LUT2 #(
		.INIT('h8)
	) name8332 (
		_w1216_,
		_w1438_,
		_w8366_
	);
	LUT4 #(
		.INIT('h135f)
	) name8333 (
		_w85_,
		_w110_,
		_w176_,
		_w378_,
		_w8367_
	);
	LUT2 #(
		.INIT('h4)
	) name8334 (
		_w426_,
		_w8367_,
		_w8368_
	);
	LUT4 #(
		.INIT('h4000)
	) name8335 (
		_w426_,
		_w1216_,
		_w1438_,
		_w8367_,
		_w8369_
	);
	LUT3 #(
		.INIT('h80)
	) name8336 (
		_w8363_,
		_w8365_,
		_w8369_,
		_w8370_
	);
	LUT3 #(
		.INIT('h80)
	) name8337 (
		_w252_,
		_w447_,
		_w921_,
		_w8371_
	);
	LUT4 #(
		.INIT('h2000)
	) name8338 (
		_w283_,
		_w386_,
		_w2379_,
		_w2563_,
		_w8372_
	);
	LUT3 #(
		.INIT('h80)
	) name8339 (
		_w1061_,
		_w1416_,
		_w8352_,
		_w8373_
	);
	LUT3 #(
		.INIT('h57)
	) name8340 (
		_w67_,
		_w158_,
		_w259_,
		_w8374_
	);
	LUT4 #(
		.INIT('h0777)
	) name8341 (
		_w106_,
		_w41_,
		_w65_,
		_w419_,
		_w8375_
	);
	LUT4 #(
		.INIT('h153f)
	) name8342 (
		_w59_,
		_w93_,
		_w184_,
		_w201_,
		_w8376_
	);
	LUT4 #(
		.INIT('h8000)
	) name8343 (
		_w820_,
		_w8376_,
		_w8374_,
		_w8375_,
		_w8377_
	);
	LUT4 #(
		.INIT('h8000)
	) name8344 (
		_w8373_,
		_w8377_,
		_w8371_,
		_w8372_,
		_w8378_
	);
	LUT3 #(
		.INIT('h80)
	) name8345 (
		_w7995_,
		_w8370_,
		_w8378_,
		_w8379_
	);
	LUT2 #(
		.INIT('h8)
	) name8346 (
		_w7579_,
		_w8379_,
		_w8380_
	);
	LUT4 #(
		.INIT('h0045)
	) name8347 (
		_w8357_,
		_w8359_,
		_w8361_,
		_w8380_,
		_w8381_
	);
	LUT4 #(
		.INIT('hba00)
	) name8348 (
		_w8357_,
		_w8359_,
		_w8361_,
		_w8380_,
		_w8382_
	);
	LUT3 #(
		.INIT('h28)
	) name8349 (
		_w377_,
		_w7062_,
		_w8358_,
		_w8383_
	);
	LUT4 #(
		.INIT('ha802)
	) name8350 (
		_w376_,
		_w6689_,
		_w6911_,
		_w6913_,
		_w8384_
	);
	LUT4 #(
		.INIT('h007d)
	) name8351 (
		_w2407_,
		_w6914_,
		_w6916_,
		_w8384_,
		_w8385_
	);
	LUT3 #(
		.INIT('h70)
	) name8352 (
		_w2527_,
		_w7062_,
		_w8385_,
		_w8386_
	);
	LUT4 #(
		.INIT('h4544)
	) name8353 (
		_w8381_,
		_w8382_,
		_w8383_,
		_w8386_,
		_w8387_
	);
	LUT4 #(
		.INIT('hba20)
	) name8354 (
		_w8335_,
		_w8336_,
		_w8340_,
		_w8387_,
		_w8388_
	);
	LUT4 #(
		.INIT('hba20)
	) name8355 (
		_w8322_,
		_w8323_,
		_w8328_,
		_w8388_,
		_w8389_
	);
	LUT4 #(
		.INIT('h4c00)
	) name8356 (
		_w377_,
		_w8297_,
		_w8298_,
		_w8301_,
		_w8390_
	);
	LUT4 #(
		.INIT('h93cc)
	) name8357 (
		_w377_,
		_w8297_,
		_w8298_,
		_w8301_,
		_w8391_
	);
	LUT3 #(
		.INIT('h54)
	) name8358 (
		_w8302_,
		_w8389_,
		_w8390_,
		_w8392_
	);
	LUT3 #(
		.INIT('h20)
	) name8359 (
		_w8278_,
		_w8279_,
		_w8283_,
		_w8393_
	);
	LUT3 #(
		.INIT('h9a)
	) name8360 (
		_w8278_,
		_w8279_,
		_w8283_,
		_w8394_
	);
	LUT3 #(
		.INIT('h54)
	) name8361 (
		_w8284_,
		_w8392_,
		_w8393_,
		_w8395_
	);
	LUT3 #(
		.INIT('h20)
	) name8362 (
		_w8243_,
		_w8244_,
		_w8249_,
		_w8396_
	);
	LUT3 #(
		.INIT('h9a)
	) name8363 (
		_w8243_,
		_w8244_,
		_w8249_,
		_w8397_
	);
	LUT4 #(
		.INIT('h93cc)
	) name8364 (
		_w377_,
		_w8226_,
		_w8227_,
		_w8230_,
		_w8398_
	);
	LUT4 #(
		.INIT('h1700)
	) name8365 (
		_w8243_,
		_w8250_,
		_w8395_,
		_w8398_,
		_w8399_
	);
	LUT3 #(
		.INIT('h9a)
	) name8366 (
		_w8213_,
		_w8214_,
		_w8218_,
		_w8400_
	);
	LUT4 #(
		.INIT('h0155)
	) name8367 (
		_w8219_,
		_w8231_,
		_w8399_,
		_w8400_,
		_w8401_
	);
	LUT3 #(
		.INIT('h20)
	) name8368 (
		_w8196_,
		_w8197_,
		_w8202_,
		_w8402_
	);
	LUT3 #(
		.INIT('h9a)
	) name8369 (
		_w8196_,
		_w8197_,
		_w8202_,
		_w8403_
	);
	LUT3 #(
		.INIT('h54)
	) name8370 (
		_w8203_,
		_w8401_,
		_w8402_,
		_w8404_
	);
	LUT4 #(
		.INIT('h0069)
	) name8371 (
		_w7845_,
		_w8004_,
		_w8009_,
		_w8404_,
		_w8405_
	);
	LUT4 #(
		.INIT('h9600)
	) name8372 (
		_w7845_,
		_w8004_,
		_w8009_,
		_w8404_,
		_w8406_
	);
	LUT4 #(
		.INIT('h6996)
	) name8373 (
		_w7845_,
		_w8004_,
		_w8009_,
		_w8404_,
		_w8407_
	);
	LUT4 #(
		.INIT('h2228)
	) name8374 (
		_w2549_,
		_w5067_,
		_w5282_,
		_w6939_,
		_w8408_
	);
	LUT4 #(
		.INIT('h007d)
	) name8375 (
		_w2617_,
		_w6940_,
		_w6942_,
		_w8408_,
		_w8409_
	);
	LUT3 #(
		.INIT('h70)
	) name8376 (
		_w2854_,
		_w7038_,
		_w8409_,
		_w8410_
	);
	LUT4 #(
		.INIT('h95aa)
	) name8377 (
		\a[29] ,
		_w2550_,
		_w8018_,
		_w8410_,
		_w8411_
	);
	LUT3 #(
		.INIT('h54)
	) name8378 (
		_w8405_,
		_w8406_,
		_w8411_,
		_w8412_
	);
	LUT2 #(
		.INIT('h4)
	) name8379 (
		_w8178_,
		_w8184_,
		_w8413_
	);
	LUT2 #(
		.INIT('h9)
	) name8380 (
		_w8178_,
		_w8184_,
		_w8414_
	);
	LUT3 #(
		.INIT('h96)
	) name8381 (
		_w8010_,
		_w8012_,
		_w8176_,
		_w8415_
	);
	LUT4 #(
		.INIT('h2b00)
	) name8382 (
		_w8178_,
		_w8184_,
		_w8412_,
		_w8415_,
		_w8416_
	);
	LUT2 #(
		.INIT('h9)
	) name8383 (
		_w8017_,
		_w8022_,
		_w8417_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8384 (
		_w2549_,
		_w4695_,
		_w6944_,
		_w6946_,
		_w8418_
	);
	LUT4 #(
		.INIT('h007d)
	) name8385 (
		_w2617_,
		_w6947_,
		_w6949_,
		_w8418_,
		_w8419_
	);
	LUT3 #(
		.INIT('h70)
	) name8386 (
		_w2854_,
		_w7032_,
		_w8419_,
		_w8420_
	);
	LUT4 #(
		.INIT('h95aa)
	) name8387 (
		\a[29] ,
		_w2550_,
		_w7882_,
		_w8420_,
		_w8421_
	);
	LUT4 #(
		.INIT('h1f01)
	) name8388 (
		_w8177_,
		_w8416_,
		_w8417_,
		_w8421_,
		_w8422_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8389 (
		_w2875_,
		_w7028_,
		_w7103_,
		_w7104_,
		_w8423_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8390 (
		_w2986_,
		_w3882_,
		_w6954_,
		_w6956_,
		_w8424_
	);
	LUT3 #(
		.INIT('h82)
	) name8391 (
		_w2874_,
		_w4030_,
		_w6952_,
		_w8425_
	);
	LUT3 #(
		.INIT('h07)
	) name8392 (
		_w2975_,
		_w7026_,
		_w8425_,
		_w8426_
	);
	LUT2 #(
		.INIT('h4)
	) name8393 (
		_w8424_,
		_w8426_,
		_w8427_
	);
	LUT3 #(
		.INIT('h9a)
	) name8394 (
		\a[26] ,
		_w8423_,
		_w8427_,
		_w8428_
	);
	LUT3 #(
		.INIT('hd4)
	) name8395 (
		_w8169_,
		_w8422_,
		_w8428_,
		_w8429_
	);
	LUT3 #(
		.INIT('h82)
	) name8396 (
		_w37_,
		_w7111_,
		_w7113_,
		_w8430_
	);
	LUT3 #(
		.INIT('h82)
	) name8397 (
		_w3262_,
		_w6960_,
		_w6962_,
		_w8431_
	);
	LUT2 #(
		.INIT('h8)
	) name8398 (
		_w3214_,
		_w7020_,
		_w8432_
	);
	LUT4 #(
		.INIT('h2228)
	) name8399 (
		_w3249_,
		_w3409_,
		_w3650_,
		_w6959_,
		_w8433_
	);
	LUT2 #(
		.INIT('h1)
	) name8400 (
		_w8432_,
		_w8433_,
		_w8434_
	);
	LUT2 #(
		.INIT('h4)
	) name8401 (
		_w8431_,
		_w8434_,
		_w8435_
	);
	LUT3 #(
		.INIT('h9a)
	) name8402 (
		\a[23] ,
		_w8430_,
		_w8435_,
		_w8436_
	);
	LUT3 #(
		.INIT('hd4)
	) name8403 (
		_w8168_,
		_w8429_,
		_w8436_,
		_w8437_
	);
	LUT3 #(
		.INIT('h54)
	) name8404 (
		_w8165_,
		_w8166_,
		_w8437_,
		_w8438_
	);
	LUT3 #(
		.INIT('h69)
	) name8405 (
		_w8118_,
		_w8119_,
		_w8125_,
		_w8439_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8406 (
		_w3312_,
		_w7010_,
		_w7121_,
		_w7122_,
		_w8440_
	);
	LUT4 #(
		.INIT('h04c8)
	) name8407 (
		_w2983_,
		_w3654_,
		_w6972_,
		_w6974_,
		_w8441_
	);
	LUT3 #(
		.INIT('h82)
	) name8408 (
		_w3311_,
		_w6967_,
		_w6969_,
		_w8442_
	);
	LUT3 #(
		.INIT('h07)
	) name8409 (
		_w3645_,
		_w7008_,
		_w8442_,
		_w8443_
	);
	LUT2 #(
		.INIT('h4)
	) name8410 (
		_w8441_,
		_w8443_,
		_w8444_
	);
	LUT3 #(
		.INIT('h9a)
	) name8411 (
		\a[20] ,
		_w8440_,
		_w8444_,
		_w8445_
	);
	LUT3 #(
		.INIT('he8)
	) name8412 (
		_w8438_,
		_w8439_,
		_w8445_,
		_w8446_
	);
	LUT3 #(
		.INIT('h82)
	) name8413 (
		_w3710_,
		_w7129_,
		_w7131_,
		_w8447_
	);
	LUT3 #(
		.INIT('h84)
	) name8414 (
		_w2546_,
		_w3886_,
		_w6981_,
		_w8448_
	);
	LUT2 #(
		.INIT('h8)
	) name8415 (
		_w3709_,
		_w7002_,
		_w8449_
	);
	LUT4 #(
		.INIT('h04c8)
	) name8416 (
		_w2622_,
		_w3877_,
		_w6978_,
		_w6980_,
		_w8450_
	);
	LUT2 #(
		.INIT('h1)
	) name8417 (
		_w8449_,
		_w8450_,
		_w8451_
	);
	LUT2 #(
		.INIT('h4)
	) name8418 (
		_w8448_,
		_w8451_,
		_w8452_
	);
	LUT3 #(
		.INIT('h9a)
	) name8419 (
		\a[17] ,
		_w8447_,
		_w8452_,
		_w8453_
	);
	LUT3 #(
		.INIT('hd4)
	) name8420 (
		_w8160_,
		_w8446_,
		_w8453_,
		_w8454_
	);
	LUT3 #(
		.INIT('h54)
	) name8421 (
		_w8157_,
		_w8158_,
		_w8454_,
		_w8455_
	);
	LUT4 #(
		.INIT('h54ab)
	) name8422 (
		_w8090_,
		_w8091_,
		_w8134_,
		_w8136_,
		_w8456_
	);
	LUT2 #(
		.INIT('h6)
	) name8423 (
		_w8144_,
		_w8456_,
		_w8457_
	);
	LUT4 #(
		.INIT('h0a02)
	) name8424 (
		_w4034_,
		_w7169_,
		_w7419_,
		_w7686_,
		_w8458_
	);
	LUT3 #(
		.INIT('h28)
	) name8425 (
		_w4033_,
		_w7136_,
		_w7168_,
		_w8459_
	);
	LUT3 #(
		.INIT('h40)
	) name8426 (
		_w4382_,
		_w7136_,
		_w7167_,
		_w8460_
	);
	LUT3 #(
		.INIT('h31)
	) name8427 (
		_w8081_,
		_w8459_,
		_w8460_,
		_w8461_
	);
	LUT3 #(
		.INIT('h9a)
	) name8428 (
		\a[14] ,
		_w8458_,
		_w8461_,
		_w8462_
	);
	LUT3 #(
		.INIT('he8)
	) name8429 (
		_w8455_,
		_w8457_,
		_w8462_,
		_w8463_
	);
	LUT2 #(
		.INIT('h2)
	) name8430 (
		_w8152_,
		_w8463_,
		_w8464_
	);
	LUT2 #(
		.INIT('h4)
	) name8431 (
		_w8152_,
		_w8463_,
		_w8465_
	);
	LUT2 #(
		.INIT('h9)
	) name8432 (
		_w8152_,
		_w8463_,
		_w8466_
	);
	LUT3 #(
		.INIT('h28)
	) name8433 (
		_w4367_,
		_w7136_,
		_w7168_,
		_w8467_
	);
	LUT4 #(
		.INIT('h028a)
	) name8434 (
		_w4382_,
		_w7136_,
		_w7166_,
		_w7167_,
		_w8468_
	);
	LUT4 #(
		.INIT('h04c8)
	) name8435 (
		_w2411_,
		_w4033_,
		_w6983_,
		_w6993_,
		_w8469_
	);
	LUT3 #(
		.INIT('h01)
	) name8436 (
		_w8468_,
		_w8469_,
		_w8467_,
		_w8470_
	);
	LUT4 #(
		.INIT('h95aa)
	) name8437 (
		\a[14] ,
		_w4034_,
		_w7696_,
		_w8470_,
		_w8471_
	);
	LUT3 #(
		.INIT('h96)
	) name8438 (
		_w8160_,
		_w8446_,
		_w8453_,
		_w8472_
	);
	LUT4 #(
		.INIT('h04c8)
	) name8439 (
		_w3257_,
		_w3311_,
		_w6964_,
		_w6966_,
		_w8473_
	);
	LUT4 #(
		.INIT('h007d)
	) name8440 (
		_w3645_,
		_w6967_,
		_w6969_,
		_w8473_,
		_w8474_
	);
	LUT3 #(
		.INIT('h70)
	) name8441 (
		_w3654_,
		_w7008_,
		_w8474_,
		_w8475_
	);
	LUT4 #(
		.INIT('h95aa)
	) name8442 (
		\a[20] ,
		_w3312_,
		_w7403_,
		_w8475_,
		_w8476_
	);
	LUT3 #(
		.INIT('h09)
	) name8443 (
		_w8167_,
		_w8437_,
		_w8476_,
		_w8477_
	);
	LUT3 #(
		.INIT('h60)
	) name8444 (
		_w8167_,
		_w8437_,
		_w8476_,
		_w8478_
	);
	LUT3 #(
		.INIT('h96)
	) name8445 (
		_w8167_,
		_w8437_,
		_w8476_,
		_w8479_
	);
	LUT3 #(
		.INIT('h96)
	) name8446 (
		_w8168_,
		_w8429_,
		_w8436_,
		_w8480_
	);
	LUT4 #(
		.INIT('h2228)
	) name8447 (
		_w2874_,
		_w4099_,
		_w4378_,
		_w6951_,
		_w8481_
	);
	LUT4 #(
		.INIT('h007d)
	) name8448 (
		_w2975_,
		_w4030_,
		_w6952_,
		_w8481_,
		_w8482_
	);
	LUT3 #(
		.INIT('h70)
	) name8449 (
		_w2986_,
		_w7026_,
		_w8482_,
		_w8483_
	);
	LUT4 #(
		.INIT('h95aa)
	) name8450 (
		\a[26] ,
		_w2875_,
		_w7562_,
		_w8483_,
		_w8484_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name8451 (
		_w8177_,
		_w8416_,
		_w8417_,
		_w8421_,
		_w8485_
	);
	LUT4 #(
		.INIT('h54ab)
	) name8452 (
		_w8185_,
		_w8412_,
		_w8413_,
		_w8415_,
		_w8486_
	);
	LUT3 #(
		.INIT('h82)
	) name8453 (
		_w2550_,
		_w7093_,
		_w7095_,
		_w8487_
	);
	LUT3 #(
		.INIT('h82)
	) name8454 (
		_w2854_,
		_w6947_,
		_w6949_,
		_w8488_
	);
	LUT2 #(
		.INIT('h8)
	) name8455 (
		_w2549_,
		_w7038_,
		_w8489_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8456 (
		_w2617_,
		_w4695_,
		_w6944_,
		_w6946_,
		_w8490_
	);
	LUT2 #(
		.INIT('h1)
	) name8457 (
		_w8489_,
		_w8490_,
		_w8491_
	);
	LUT2 #(
		.INIT('h4)
	) name8458 (
		_w8488_,
		_w8491_,
		_w8492_
	);
	LUT3 #(
		.INIT('h9a)
	) name8459 (
		\a[29] ,
		_w8487_,
		_w8492_,
		_w8493_
	);
	LUT3 #(
		.INIT('h82)
	) name8460 (
		_w2875_,
		_w7099_,
		_w7101_,
		_w8494_
	);
	LUT3 #(
		.INIT('h82)
	) name8461 (
		_w2986_,
		_w4030_,
		_w6952_,
		_w8495_
	);
	LUT2 #(
		.INIT('h8)
	) name8462 (
		_w2874_,
		_w7032_,
		_w8496_
	);
	LUT4 #(
		.INIT('h2228)
	) name8463 (
		_w2975_,
		_w4099_,
		_w4378_,
		_w6951_,
		_w8497_
	);
	LUT2 #(
		.INIT('h1)
	) name8464 (
		_w8496_,
		_w8497_,
		_w8498_
	);
	LUT2 #(
		.INIT('h4)
	) name8465 (
		_w8495_,
		_w8498_,
		_w8499_
	);
	LUT3 #(
		.INIT('h9a)
	) name8466 (
		\a[26] ,
		_w8494_,
		_w8499_,
		_w8500_
	);
	LUT3 #(
		.INIT('hd4)
	) name8467 (
		_w8486_,
		_w8493_,
		_w8500_,
		_w8501_
	);
	LUT3 #(
		.INIT('hb2)
	) name8468 (
		_w8484_,
		_w8485_,
		_w8501_,
		_w8502_
	);
	LUT3 #(
		.INIT('h96)
	) name8469 (
		_w8169_,
		_w8422_,
		_w8428_,
		_w8503_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8470 (
		_w37_,
		_w7022_,
		_w7109_,
		_w7110_,
		_w8504_
	);
	LUT4 #(
		.INIT('h2228)
	) name8471 (
		_w3262_,
		_w3409_,
		_w3650_,
		_w6959_,
		_w8505_
	);
	LUT3 #(
		.INIT('h82)
	) name8472 (
		_w3214_,
		_w3706_,
		_w6957_,
		_w8506_
	);
	LUT3 #(
		.INIT('h07)
	) name8473 (
		_w3249_,
		_w7020_,
		_w8506_,
		_w8507_
	);
	LUT2 #(
		.INIT('h4)
	) name8474 (
		_w8505_,
		_w8507_,
		_w8508_
	);
	LUT3 #(
		.INIT('h9a)
	) name8475 (
		\a[23] ,
		_w8504_,
		_w8508_,
		_w8509_
	);
	LUT3 #(
		.INIT('hb2)
	) name8476 (
		_w8502_,
		_w8503_,
		_w8509_,
		_w8510_
	);
	LUT3 #(
		.INIT('h82)
	) name8477 (
		_w3312_,
		_w7117_,
		_w7119_,
		_w8511_
	);
	LUT3 #(
		.INIT('h82)
	) name8478 (
		_w3654_,
		_w6967_,
		_w6969_,
		_w8512_
	);
	LUT2 #(
		.INIT('h8)
	) name8479 (
		_w3311_,
		_w7014_,
		_w8513_
	);
	LUT4 #(
		.INIT('h04c8)
	) name8480 (
		_w3257_,
		_w3645_,
		_w6964_,
		_w6966_,
		_w8514_
	);
	LUT2 #(
		.INIT('h1)
	) name8481 (
		_w8513_,
		_w8514_,
		_w8515_
	);
	LUT2 #(
		.INIT('h4)
	) name8482 (
		_w8512_,
		_w8515_,
		_w8516_
	);
	LUT3 #(
		.INIT('h9a)
	) name8483 (
		\a[20] ,
		_w8511_,
		_w8516_,
		_w8517_
	);
	LUT3 #(
		.INIT('hd4)
	) name8484 (
		_w8480_,
		_w8510_,
		_w8517_,
		_w8518_
	);
	LUT3 #(
		.INIT('h54)
	) name8485 (
		_w8477_,
		_w8478_,
		_w8518_,
		_w8519_
	);
	LUT3 #(
		.INIT('h69)
	) name8486 (
		_w8438_,
		_w8439_,
		_w8445_,
		_w8520_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8487 (
		_w3710_,
		_w7004_,
		_w7127_,
		_w7128_,
		_w8521_
	);
	LUT4 #(
		.INIT('h04c8)
	) name8488 (
		_w2622_,
		_w3886_,
		_w6978_,
		_w6980_,
		_w8522_
	);
	LUT3 #(
		.INIT('h84)
	) name8489 (
		_w2872_,
		_w3709_,
		_w6975_,
		_w8523_
	);
	LUT3 #(
		.INIT('h07)
	) name8490 (
		_w3877_,
		_w7002_,
		_w8523_,
		_w8524_
	);
	LUT2 #(
		.INIT('h4)
	) name8491 (
		_w8522_,
		_w8524_,
		_w8525_
	);
	LUT3 #(
		.INIT('h9a)
	) name8492 (
		\a[17] ,
		_w8521_,
		_w8525_,
		_w8526_
	);
	LUT3 #(
		.INIT('hb2)
	) name8493 (
		_w8519_,
		_w8520_,
		_w8526_,
		_w8527_
	);
	LUT3 #(
		.INIT('h82)
	) name8494 (
		_w4034_,
		_w7135_,
		_w7172_,
		_w8528_
	);
	LUT3 #(
		.INIT('h28)
	) name8495 (
		_w4382_,
		_w7136_,
		_w7168_,
		_w8529_
	);
	LUT2 #(
		.INIT('h8)
	) name8496 (
		_w4033_,
		_w6996_,
		_w8530_
	);
	LUT4 #(
		.INIT('h04c8)
	) name8497 (
		_w2411_,
		_w4367_,
		_w6983_,
		_w6993_,
		_w8531_
	);
	LUT2 #(
		.INIT('h1)
	) name8498 (
		_w8530_,
		_w8531_,
		_w8532_
	);
	LUT2 #(
		.INIT('h4)
	) name8499 (
		_w8529_,
		_w8532_,
		_w8533_
	);
	LUT3 #(
		.INIT('h9a)
	) name8500 (
		\a[14] ,
		_w8528_,
		_w8533_,
		_w8534_
	);
	LUT4 #(
		.INIT('h0445)
	) name8501 (
		_w8471_,
		_w8472_,
		_w8527_,
		_w8534_,
		_w8535_
	);
	LUT2 #(
		.INIT('h9)
	) name8502 (
		_w8159_,
		_w8454_,
		_w8536_
	);
	LUT4 #(
		.INIT('ha220)
	) name8503 (
		_w8471_,
		_w8472_,
		_w8527_,
		_w8534_,
		_w8537_
	);
	LUT4 #(
		.INIT('h599a)
	) name8504 (
		_w8471_,
		_w8472_,
		_w8527_,
		_w8534_,
		_w8538_
	);
	LUT3 #(
		.INIT('h51)
	) name8505 (
		_w8535_,
		_w8536_,
		_w8537_,
		_w8539_
	);
	LUT3 #(
		.INIT('h69)
	) name8506 (
		_w8455_,
		_w8457_,
		_w8462_,
		_w8540_
	);
	LUT2 #(
		.INIT('h4)
	) name8507 (
		_w8539_,
		_w8540_,
		_w8541_
	);
	LUT2 #(
		.INIT('h6)
	) name8508 (
		_w8536_,
		_w8538_,
		_w8542_
	);
	LUT4 #(
		.INIT('h028a)
	) name8509 (
		_w4458_,
		_w7136_,
		_w7166_,
		_w7167_,
		_w8543_
	);
	LUT4 #(
		.INIT('h781e)
	) name8510 (
		\a[8] ,
		\a[9] ,
		\a[10] ,
		\a[11] ,
		_w8544_
	);
	LUT3 #(
		.INIT('hb0)
	) name8511 (
		_w7136_,
		_w7166_,
		_w8544_,
		_w8545_
	);
	LUT2 #(
		.INIT('h1)
	) name8512 (
		_w8543_,
		_w8545_,
		_w8546_
	);
	LUT4 #(
		.INIT('h5700)
	) name8513 (
		_w4459_,
		_w7418_,
		_w7419_,
		_w8546_,
		_w8547_
	);
	LUT2 #(
		.INIT('h6)
	) name8514 (
		\a[11] ,
		_w8547_,
		_w8548_
	);
	LUT4 #(
		.INIT('h04c8)
	) name8515 (
		_w2983_,
		_w3709_,
		_w6972_,
		_w6974_,
		_w8549_
	);
	LUT4 #(
		.INIT('h007b)
	) name8516 (
		_w2872_,
		_w3877_,
		_w6975_,
		_w8549_,
		_w8550_
	);
	LUT3 #(
		.INIT('h70)
	) name8517 (
		_w3886_,
		_w7002_,
		_w8550_,
		_w8551_
	);
	LUT4 #(
		.INIT('h95aa)
	) name8518 (
		\a[17] ,
		_w3710_,
		_w7426_,
		_w8551_,
		_w8552_
	);
	LUT3 #(
		.INIT('h09)
	) name8519 (
		_w8479_,
		_w8518_,
		_w8552_,
		_w8553_
	);
	LUT3 #(
		.INIT('h60)
	) name8520 (
		_w8479_,
		_w8518_,
		_w8552_,
		_w8554_
	);
	LUT3 #(
		.INIT('h96)
	) name8521 (
		_w8479_,
		_w8518_,
		_w8552_,
		_w8555_
	);
	LUT3 #(
		.INIT('h96)
	) name8522 (
		_w8480_,
		_w8510_,
		_w8517_,
		_w8556_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8523 (
		_w3214_,
		_w3882_,
		_w6954_,
		_w6956_,
		_w8557_
	);
	LUT4 #(
		.INIT('h007d)
	) name8524 (
		_w3249_,
		_w3706_,
		_w6957_,
		_w8557_,
		_w8558_
	);
	LUT3 #(
		.INIT('h70)
	) name8525 (
		_w3262_,
		_w7020_,
		_w8558_,
		_w8559_
	);
	LUT4 #(
		.INIT('h95aa)
	) name8526 (
		\a[23] ,
		_w37_,
		_w7465_,
		_w8559_,
		_w8560_
	);
	LUT4 #(
		.INIT('h0096)
	) name8527 (
		_w8484_,
		_w8485_,
		_w8501_,
		_w8560_,
		_w8561_
	);
	LUT4 #(
		.INIT('h6900)
	) name8528 (
		_w8484_,
		_w8485_,
		_w8501_,
		_w8560_,
		_w8562_
	);
	LUT4 #(
		.INIT('h9669)
	) name8529 (
		_w8484_,
		_w8485_,
		_w8501_,
		_w8560_,
		_w8563_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8530 (
		_w2550_,
		_w7040_,
		_w7091_,
		_w7092_,
		_w8564_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8531 (
		_w2854_,
		_w4695_,
		_w6944_,
		_w6946_,
		_w8565_
	);
	LUT3 #(
		.INIT('h82)
	) name8532 (
		_w2549_,
		_w6940_,
		_w6942_,
		_w8566_
	);
	LUT3 #(
		.INIT('h07)
	) name8533 (
		_w2617_,
		_w7038_,
		_w8566_,
		_w8567_
	);
	LUT2 #(
		.INIT('h4)
	) name8534 (
		_w8565_,
		_w8567_,
		_w8568_
	);
	LUT3 #(
		.INIT('h9a)
	) name8535 (
		\a[29] ,
		_w8564_,
		_w8568_,
		_w8569_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8536 (
		_w2875_,
		_w7034_,
		_w7097_,
		_w7098_,
		_w8570_
	);
	LUT4 #(
		.INIT('h2228)
	) name8537 (
		_w2986_,
		_w4099_,
		_w4378_,
		_w6951_,
		_w8571_
	);
	LUT3 #(
		.INIT('h82)
	) name8538 (
		_w2874_,
		_w6947_,
		_w6949_,
		_w8572_
	);
	LUT3 #(
		.INIT('h07)
	) name8539 (
		_w2975_,
		_w7032_,
		_w8572_,
		_w8573_
	);
	LUT2 #(
		.INIT('h4)
	) name8540 (
		_w8571_,
		_w8573_,
		_w8574_
	);
	LUT3 #(
		.INIT('h9a)
	) name8541 (
		\a[26] ,
		_w8570_,
		_w8574_,
		_w8575_
	);
	LUT4 #(
		.INIT('hf660)
	) name8542 (
		_w8412_,
		_w8414_,
		_w8569_,
		_w8575_,
		_w8576_
	);
	LUT4 #(
		.INIT('h0096)
	) name8543 (
		_w8486_,
		_w8493_,
		_w8500_,
		_w8576_,
		_w8577_
	);
	LUT4 #(
		.INIT('h6900)
	) name8544 (
		_w8486_,
		_w8493_,
		_w8500_,
		_w8576_,
		_w8578_
	);
	LUT3 #(
		.INIT('h82)
	) name8545 (
		_w37_,
		_w7105_,
		_w7107_,
		_w8579_
	);
	LUT3 #(
		.INIT('h82)
	) name8546 (
		_w3262_,
		_w3706_,
		_w6957_,
		_w8580_
	);
	LUT2 #(
		.INIT('h8)
	) name8547 (
		_w3214_,
		_w7026_,
		_w8581_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8548 (
		_w3249_,
		_w3882_,
		_w6954_,
		_w6956_,
		_w8582_
	);
	LUT2 #(
		.INIT('h1)
	) name8549 (
		_w8581_,
		_w8582_,
		_w8583_
	);
	LUT2 #(
		.INIT('h4)
	) name8550 (
		_w8580_,
		_w8583_,
		_w8584_
	);
	LUT3 #(
		.INIT('h9a)
	) name8551 (
		\a[23] ,
		_w8579_,
		_w8584_,
		_w8585_
	);
	LUT3 #(
		.INIT('h54)
	) name8552 (
		_w8577_,
		_w8578_,
		_w8585_,
		_w8586_
	);
	LUT3 #(
		.INIT('h54)
	) name8553 (
		_w8561_,
		_w8562_,
		_w8586_,
		_w8587_
	);
	LUT3 #(
		.INIT('h69)
	) name8554 (
		_w8502_,
		_w8503_,
		_w8509_,
		_w8588_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8555 (
		_w3312_,
		_w7016_,
		_w7115_,
		_w7116_,
		_w8589_
	);
	LUT4 #(
		.INIT('h04c8)
	) name8556 (
		_w3257_,
		_w3654_,
		_w6964_,
		_w6966_,
		_w8590_
	);
	LUT3 #(
		.INIT('h82)
	) name8557 (
		_w3311_,
		_w6960_,
		_w6962_,
		_w8591_
	);
	LUT3 #(
		.INIT('h07)
	) name8558 (
		_w3645_,
		_w7014_,
		_w8591_,
		_w8592_
	);
	LUT2 #(
		.INIT('h4)
	) name8559 (
		_w8590_,
		_w8592_,
		_w8593_
	);
	LUT3 #(
		.INIT('h9a)
	) name8560 (
		\a[20] ,
		_w8589_,
		_w8593_,
		_w8594_
	);
	LUT3 #(
		.INIT('he8)
	) name8561 (
		_w8587_,
		_w8588_,
		_w8594_,
		_w8595_
	);
	LUT3 #(
		.INIT('h82)
	) name8562 (
		_w3710_,
		_w7123_,
		_w7125_,
		_w8596_
	);
	LUT3 #(
		.INIT('h84)
	) name8563 (
		_w2872_,
		_w3886_,
		_w6975_,
		_w8597_
	);
	LUT2 #(
		.INIT('h8)
	) name8564 (
		_w3709_,
		_w7008_,
		_w8598_
	);
	LUT4 #(
		.INIT('h04c8)
	) name8565 (
		_w2983_,
		_w3877_,
		_w6972_,
		_w6974_,
		_w8599_
	);
	LUT2 #(
		.INIT('h1)
	) name8566 (
		_w8598_,
		_w8599_,
		_w8600_
	);
	LUT2 #(
		.INIT('h4)
	) name8567 (
		_w8597_,
		_w8600_,
		_w8601_
	);
	LUT3 #(
		.INIT('h9a)
	) name8568 (
		\a[17] ,
		_w8596_,
		_w8601_,
		_w8602_
	);
	LUT3 #(
		.INIT('hd4)
	) name8569 (
		_w8556_,
		_w8595_,
		_w8602_,
		_w8603_
	);
	LUT3 #(
		.INIT('h54)
	) name8570 (
		_w8553_,
		_w8554_,
		_w8603_,
		_w8604_
	);
	LUT3 #(
		.INIT('h69)
	) name8571 (
		_w8519_,
		_w8520_,
		_w8526_,
		_w8605_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8572 (
		_w4034_,
		_w6998_,
		_w7133_,
		_w7134_,
		_w8606_
	);
	LUT4 #(
		.INIT('h04c8)
	) name8573 (
		_w2411_,
		_w4382_,
		_w6983_,
		_w6993_,
		_w8607_
	);
	LUT3 #(
		.INIT('h84)
	) name8574 (
		_w2546_,
		_w4033_,
		_w6981_,
		_w8608_
	);
	LUT3 #(
		.INIT('h07)
	) name8575 (
		_w4367_,
		_w6996_,
		_w8608_,
		_w8609_
	);
	LUT2 #(
		.INIT('h4)
	) name8576 (
		_w8607_,
		_w8609_,
		_w8610_
	);
	LUT3 #(
		.INIT('h9a)
	) name8577 (
		\a[14] ,
		_w8606_,
		_w8610_,
		_w8611_
	);
	LUT4 #(
		.INIT('h0115)
	) name8578 (
		_w8548_,
		_w8604_,
		_w8605_,
		_w8611_,
		_w8612_
	);
	LUT4 #(
		.INIT('ha880)
	) name8579 (
		_w8548_,
		_w8604_,
		_w8605_,
		_w8611_,
		_w8613_
	);
	LUT3 #(
		.INIT('h96)
	) name8580 (
		_w8472_,
		_w8527_,
		_w8534_,
		_w8614_
	);
	LUT3 #(
		.INIT('h45)
	) name8581 (
		_w8612_,
		_w8613_,
		_w8614_,
		_w8615_
	);
	LUT2 #(
		.INIT('h2)
	) name8582 (
		_w8542_,
		_w8615_,
		_w8616_
	);
	LUT4 #(
		.INIT('h566a)
	) name8583 (
		_w8548_,
		_w8604_,
		_w8605_,
		_w8611_,
		_w8617_
	);
	LUT2 #(
		.INIT('h6)
	) name8584 (
		_w8614_,
		_w8617_,
		_w8618_
	);
	LUT4 #(
		.INIT('h04c8)
	) name8585 (
		_w2622_,
		_w4033_,
		_w6978_,
		_w6980_,
		_w8619_
	);
	LUT4 #(
		.INIT('h007b)
	) name8586 (
		_w2546_,
		_w4367_,
		_w6981_,
		_w8619_,
		_w8620_
	);
	LUT3 #(
		.INIT('h70)
	) name8587 (
		_w4382_,
		_w6996_,
		_w8620_,
		_w8621_
	);
	LUT4 #(
		.INIT('h95aa)
	) name8588 (
		\a[14] ,
		_w4034_,
		_w7500_,
		_w8621_,
		_w8622_
	);
	LUT3 #(
		.INIT('h09)
	) name8589 (
		_w8555_,
		_w8603_,
		_w8622_,
		_w8623_
	);
	LUT3 #(
		.INIT('h60)
	) name8590 (
		_w8555_,
		_w8603_,
		_w8622_,
		_w8624_
	);
	LUT3 #(
		.INIT('h96)
	) name8591 (
		_w8555_,
		_w8603_,
		_w8622_,
		_w8625_
	);
	LUT3 #(
		.INIT('h96)
	) name8592 (
		_w8556_,
		_w8595_,
		_w8602_,
		_w8626_
	);
	LUT4 #(
		.INIT('h2228)
	) name8593 (
		_w3311_,
		_w3409_,
		_w3650_,
		_w6959_,
		_w8627_
	);
	LUT4 #(
		.INIT('h007d)
	) name8594 (
		_w3645_,
		_w6960_,
		_w6962_,
		_w8627_,
		_w8628_
	);
	LUT3 #(
		.INIT('h70)
	) name8595 (
		_w3654_,
		_w7014_,
		_w8628_,
		_w8629_
	);
	LUT4 #(
		.INIT('h95aa)
	) name8596 (
		\a[20] ,
		_w3312_,
		_w7291_,
		_w8629_,
		_w8630_
	);
	LUT4 #(
		.INIT('h9669)
	) name8597 (
		_w8486_,
		_w8493_,
		_w8500_,
		_w8576_,
		_w8631_
	);
	LUT4 #(
		.INIT('h9669)
	) name8598 (
		_w8412_,
		_w8414_,
		_w8569_,
		_w8575_,
		_w8632_
	);
	LUT3 #(
		.INIT('h82)
	) name8599 (
		_w2550_,
		_w7087_,
		_w7089_,
		_w8633_
	);
	LUT3 #(
		.INIT('h82)
	) name8600 (
		_w2854_,
		_w6940_,
		_w6942_,
		_w8634_
	);
	LUT2 #(
		.INIT('h8)
	) name8601 (
		_w2549_,
		_w7044_,
		_w8635_
	);
	LUT4 #(
		.INIT('h2228)
	) name8602 (
		_w2617_,
		_w5067_,
		_w5282_,
		_w6939_,
		_w8636_
	);
	LUT2 #(
		.INIT('h1)
	) name8603 (
		_w8635_,
		_w8636_,
		_w8637_
	);
	LUT2 #(
		.INIT('h4)
	) name8604 (
		_w8634_,
		_w8637_,
		_w8638_
	);
	LUT2 #(
		.INIT('h9)
	) name8605 (
		_w8401_,
		_w8403_,
		_w8639_
	);
	LUT4 #(
		.INIT('h6500)
	) name8606 (
		\a[29] ,
		_w8633_,
		_w8638_,
		_w8639_,
		_w8640_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8607 (
		_w2550_,
		_w7046_,
		_w7085_,
		_w7086_,
		_w8641_
	);
	LUT4 #(
		.INIT('h2228)
	) name8608 (
		_w2854_,
		_w5067_,
		_w5282_,
		_w6939_,
		_w8642_
	);
	LUT3 #(
		.INIT('h82)
	) name8609 (
		_w2549_,
		_w6935_,
		_w6937_,
		_w8643_
	);
	LUT3 #(
		.INIT('h07)
	) name8610 (
		_w2617_,
		_w7044_,
		_w8643_,
		_w8644_
	);
	LUT2 #(
		.INIT('h4)
	) name8611 (
		_w8642_,
		_w8644_,
		_w8645_
	);
	LUT3 #(
		.INIT('h1e)
	) name8612 (
		_w8231_,
		_w8399_,
		_w8400_,
		_w8646_
	);
	LUT4 #(
		.INIT('h6500)
	) name8613 (
		\a[29] ,
		_w8641_,
		_w8645_,
		_w8646_,
		_w8647_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8614 (
		_w2549_,
		_w6043_,
		_w6933_,
		_w6934_,
		_w8648_
	);
	LUT4 #(
		.INIT('h007d)
	) name8615 (
		_w2617_,
		_w6935_,
		_w6937_,
		_w8648_,
		_w8649_
	);
	LUT3 #(
		.INIT('h70)
	) name8616 (
		_w2854_,
		_w7044_,
		_w8649_,
		_w8650_
	);
	LUT4 #(
		.INIT('h95aa)
	) name8617 (
		\a[29] ,
		_w2550_,
		_w8005_,
		_w8650_,
		_w8651_
	);
	LUT4 #(
		.INIT('h54ab)
	) name8618 (
		_w8251_,
		_w8395_,
		_w8396_,
		_w8398_,
		_w8652_
	);
	LUT2 #(
		.INIT('h4)
	) name8619 (
		_w8651_,
		_w8652_,
		_w8653_
	);
	LUT3 #(
		.INIT('h82)
	) name8620 (
		_w2550_,
		_w7081_,
		_w7083_,
		_w8654_
	);
	LUT3 #(
		.INIT('h82)
	) name8621 (
		_w2854_,
		_w6935_,
		_w6937_,
		_w8655_
	);
	LUT2 #(
		.INIT('h8)
	) name8622 (
		_w2549_,
		_w7050_,
		_w8656_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8623 (
		_w2617_,
		_w6043_,
		_w6933_,
		_w6934_,
		_w8657_
	);
	LUT2 #(
		.INIT('h1)
	) name8624 (
		_w8656_,
		_w8657_,
		_w8658_
	);
	LUT2 #(
		.INIT('h4)
	) name8625 (
		_w8655_,
		_w8658_,
		_w8659_
	);
	LUT2 #(
		.INIT('h9)
	) name8626 (
		_w8395_,
		_w8397_,
		_w8660_
	);
	LUT4 #(
		.INIT('h6500)
	) name8627 (
		\a[29] ,
		_w8654_,
		_w8659_,
		_w8660_,
		_w8661_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8628 (
		_w2550_,
		_w7052_,
		_w7079_,
		_w7080_,
		_w8662_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8629 (
		_w2854_,
		_w6043_,
		_w6933_,
		_w6934_,
		_w8663_
	);
	LUT3 #(
		.INIT('h82)
	) name8630 (
		_w2549_,
		_w6929_,
		_w6931_,
		_w8664_
	);
	LUT3 #(
		.INIT('h07)
	) name8631 (
		_w2617_,
		_w7050_,
		_w8664_,
		_w8665_
	);
	LUT2 #(
		.INIT('h4)
	) name8632 (
		_w8663_,
		_w8665_,
		_w8666_
	);
	LUT2 #(
		.INIT('h9)
	) name8633 (
		_w8392_,
		_w8394_,
		_w8667_
	);
	LUT4 #(
		.INIT('h6500)
	) name8634 (
		\a[29] ,
		_w8662_,
		_w8666_,
		_w8667_,
		_w8668_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8635 (
		_w2549_,
		_w6645_,
		_w6926_,
		_w6928_,
		_w8669_
	);
	LUT4 #(
		.INIT('h007d)
	) name8636 (
		_w2617_,
		_w6929_,
		_w6931_,
		_w8669_,
		_w8670_
	);
	LUT3 #(
		.INIT('h70)
	) name8637 (
		_w2854_,
		_w7050_,
		_w8670_,
		_w8671_
	);
	LUT4 #(
		.INIT('h95aa)
	) name8638 (
		\a[29] ,
		_w2550_,
		_w8227_,
		_w8671_,
		_w8672_
	);
	LUT2 #(
		.INIT('h9)
	) name8639 (
		_w8389_,
		_w8391_,
		_w8673_
	);
	LUT2 #(
		.INIT('h4)
	) name8640 (
		_w8672_,
		_w8673_,
		_w8674_
	);
	LUT3 #(
		.INIT('h82)
	) name8641 (
		_w2550_,
		_w7075_,
		_w7077_,
		_w8675_
	);
	LUT3 #(
		.INIT('h82)
	) name8642 (
		_w2854_,
		_w6929_,
		_w6931_,
		_w8676_
	);
	LUT2 #(
		.INIT('h8)
	) name8643 (
		_w2549_,
		_w7056_,
		_w8677_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8644 (
		_w2617_,
		_w6645_,
		_w6926_,
		_w6928_,
		_w8678_
	);
	LUT2 #(
		.INIT('h1)
	) name8645 (
		_w8677_,
		_w8678_,
		_w8679_
	);
	LUT2 #(
		.INIT('h4)
	) name8646 (
		_w8676_,
		_w8679_,
		_w8680_
	);
	LUT4 #(
		.INIT('h9a65)
	) name8647 (
		_w8322_,
		_w8323_,
		_w8328_,
		_w8388_,
		_w8681_
	);
	LUT4 #(
		.INIT('h6500)
	) name8648 (
		\a[29] ,
		_w8675_,
		_w8680_,
		_w8681_,
		_w8682_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8649 (
		_w2550_,
		_w7058_,
		_w7073_,
		_w7074_,
		_w8683_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8650 (
		_w2854_,
		_w6645_,
		_w6926_,
		_w6928_,
		_w8684_
	);
	LUT3 #(
		.INIT('h82)
	) name8651 (
		_w2549_,
		_w6922_,
		_w6924_,
		_w8685_
	);
	LUT3 #(
		.INIT('h07)
	) name8652 (
		_w2617_,
		_w7056_,
		_w8685_,
		_w8686_
	);
	LUT2 #(
		.INIT('h4)
	) name8653 (
		_w8684_,
		_w8686_,
		_w8687_
	);
	LUT4 #(
		.INIT('h9a65)
	) name8654 (
		_w8335_,
		_w8336_,
		_w8340_,
		_w8387_,
		_w8688_
	);
	LUT4 #(
		.INIT('h6500)
	) name8655 (
		\a[29] ,
		_w8683_,
		_w8687_,
		_w8688_,
		_w8689_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8656 (
		_w2549_,
		_w6669_,
		_w6919_,
		_w6921_,
		_w8690_
	);
	LUT4 #(
		.INIT('h007d)
	) name8657 (
		_w2617_,
		_w6922_,
		_w6924_,
		_w8690_,
		_w8691_
	);
	LUT3 #(
		.INIT('h70)
	) name8658 (
		_w2854_,
		_w7056_,
		_w8691_,
		_w8692_
	);
	LUT4 #(
		.INIT('h95aa)
	) name8659 (
		\a[29] ,
		_w2550_,
		_w8298_,
		_w8692_,
		_w8693_
	);
	LUT4 #(
		.INIT('h45ba)
	) name8660 (
		_w8357_,
		_w8359_,
		_w8361_,
		_w8380_,
		_w8694_
	);
	LUT3 #(
		.INIT('h4b)
	) name8661 (
		_w8383_,
		_w8386_,
		_w8694_,
		_w8695_
	);
	LUT2 #(
		.INIT('h4)
	) name8662 (
		_w8693_,
		_w8695_,
		_w8696_
	);
	LUT3 #(
		.INIT('h82)
	) name8663 (
		_w2550_,
		_w7069_,
		_w7071_,
		_w8697_
	);
	LUT3 #(
		.INIT('h82)
	) name8664 (
		_w2854_,
		_w6922_,
		_w6924_,
		_w8698_
	);
	LUT2 #(
		.INIT('h8)
	) name8665 (
		_w2549_,
		_w7062_,
		_w8699_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8666 (
		_w2617_,
		_w6669_,
		_w6919_,
		_w6921_,
		_w8700_
	);
	LUT2 #(
		.INIT('h1)
	) name8667 (
		_w8699_,
		_w8700_,
		_w8701_
	);
	LUT2 #(
		.INIT('h4)
	) name8668 (
		_w8698_,
		_w8701_,
		_w8702_
	);
	LUT3 #(
		.INIT('h9a)
	) name8669 (
		_w8357_,
		_w8359_,
		_w8361_,
		_w8703_
	);
	LUT4 #(
		.INIT('h6500)
	) name8670 (
		\a[29] ,
		_w8697_,
		_w8702_,
		_w8703_,
		_w8704_
	);
	LUT4 #(
		.INIT('h5401)
	) name8671 (
		_w375_,
		_w6689_,
		_w6911_,
		_w6913_,
		_w8705_
	);
	LUT4 #(
		.INIT('h2882)
	) name8672 (
		_w2550_,
		_w6914_,
		_w6916_,
		_w7067_,
		_w8706_
	);
	LUT4 #(
		.INIT('ha802)
	) name8673 (
		_w2617_,
		_w6689_,
		_w6911_,
		_w6913_,
		_w8707_
	);
	LUT4 #(
		.INIT('h007d)
	) name8674 (
		_w2854_,
		_w6914_,
		_w6916_,
		_w8707_,
		_w8708_
	);
	LUT4 #(
		.INIT('h5401)
	) name8675 (
		_w2548_,
		_w6689_,
		_w6911_,
		_w6913_,
		_w8709_
	);
	LUT2 #(
		.INIT('h2)
	) name8676 (
		\a[29] ,
		_w8709_,
		_w8710_
	);
	LUT3 #(
		.INIT('h40)
	) name8677 (
		_w8706_,
		_w8708_,
		_w8710_,
		_w8711_
	);
	LUT3 #(
		.INIT('h28)
	) name8678 (
		_w2550_,
		_w7062_,
		_w8358_,
		_w8712_
	);
	LUT4 #(
		.INIT('ha802)
	) name8679 (
		_w2549_,
		_w6689_,
		_w6911_,
		_w6913_,
		_w8713_
	);
	LUT4 #(
		.INIT('h007d)
	) name8680 (
		_w2617_,
		_w6914_,
		_w6916_,
		_w8713_,
		_w8714_
	);
	LUT3 #(
		.INIT('h70)
	) name8681 (
		_w2854_,
		_w7062_,
		_w8714_,
		_w8715_
	);
	LUT4 #(
		.INIT('h0800)
	) name8682 (
		_w8705_,
		_w8711_,
		_w8712_,
		_w8715_,
		_w8716_
	);
	LUT3 #(
		.INIT('h28)
	) name8683 (
		_w2550_,
		_w7065_,
		_w7068_,
		_w8717_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8684 (
		_w2854_,
		_w6669_,
		_w6919_,
		_w6921_,
		_w8718_
	);
	LUT3 #(
		.INIT('h82)
	) name8685 (
		_w2549_,
		_w6914_,
		_w6916_,
		_w8719_
	);
	LUT3 #(
		.INIT('h07)
	) name8686 (
		_w2617_,
		_w7062_,
		_w8719_,
		_w8720_
	);
	LUT2 #(
		.INIT('h4)
	) name8687 (
		_w8718_,
		_w8720_,
		_w8721_
	);
	LUT4 #(
		.INIT('ha6aa)
	) name8688 (
		_w8705_,
		_w8711_,
		_w8712_,
		_w8715_,
		_w8722_
	);
	LUT4 #(
		.INIT('h6500)
	) name8689 (
		\a[29] ,
		_w8717_,
		_w8721_,
		_w8722_,
		_w8723_
	);
	LUT2 #(
		.INIT('h1)
	) name8690 (
		_w8716_,
		_w8723_,
		_w8724_
	);
	LUT4 #(
		.INIT('h009a)
	) name8691 (
		\a[29] ,
		_w8697_,
		_w8702_,
		_w8703_,
		_w8725_
	);
	LUT4 #(
		.INIT('h9a65)
	) name8692 (
		\a[29] ,
		_w8697_,
		_w8702_,
		_w8703_,
		_w8726_
	);
	LUT3 #(
		.INIT('h54)
	) name8693 (
		_w8704_,
		_w8724_,
		_w8725_,
		_w8727_
	);
	LUT2 #(
		.INIT('h2)
	) name8694 (
		_w8693_,
		_w8695_,
		_w8728_
	);
	LUT2 #(
		.INIT('h9)
	) name8695 (
		_w8693_,
		_w8695_,
		_w8729_
	);
	LUT4 #(
		.INIT('h9a65)
	) name8696 (
		\a[29] ,
		_w8683_,
		_w8687_,
		_w8688_,
		_w8730_
	);
	LUT4 #(
		.INIT('h4d00)
	) name8697 (
		_w8693_,
		_w8695_,
		_w8727_,
		_w8730_,
		_w8731_
	);
	LUT4 #(
		.INIT('h9a65)
	) name8698 (
		\a[29] ,
		_w8675_,
		_w8680_,
		_w8681_,
		_w8732_
	);
	LUT4 #(
		.INIT('h0155)
	) name8699 (
		_w8682_,
		_w8689_,
		_w8731_,
		_w8732_,
		_w8733_
	);
	LUT2 #(
		.INIT('h2)
	) name8700 (
		_w8672_,
		_w8673_,
		_w8734_
	);
	LUT2 #(
		.INIT('h9)
	) name8701 (
		_w8672_,
		_w8673_,
		_w8735_
	);
	LUT4 #(
		.INIT('h9a65)
	) name8702 (
		\a[29] ,
		_w8662_,
		_w8666_,
		_w8667_,
		_w8736_
	);
	LUT4 #(
		.INIT('h4d00)
	) name8703 (
		_w8672_,
		_w8673_,
		_w8733_,
		_w8736_,
		_w8737_
	);
	LUT4 #(
		.INIT('h9a65)
	) name8704 (
		\a[29] ,
		_w8654_,
		_w8659_,
		_w8660_,
		_w8738_
	);
	LUT4 #(
		.INIT('h0155)
	) name8705 (
		_w8661_,
		_w8668_,
		_w8737_,
		_w8738_,
		_w8739_
	);
	LUT2 #(
		.INIT('h2)
	) name8706 (
		_w8651_,
		_w8652_,
		_w8740_
	);
	LUT2 #(
		.INIT('h9)
	) name8707 (
		_w8651_,
		_w8652_,
		_w8741_
	);
	LUT4 #(
		.INIT('h9a65)
	) name8708 (
		\a[29] ,
		_w8641_,
		_w8645_,
		_w8646_,
		_w8742_
	);
	LUT4 #(
		.INIT('h4d00)
	) name8709 (
		_w8651_,
		_w8652_,
		_w8739_,
		_w8742_,
		_w8743_
	);
	LUT4 #(
		.INIT('h9a65)
	) name8710 (
		\a[29] ,
		_w8633_,
		_w8638_,
		_w8639_,
		_w8744_
	);
	LUT4 #(
		.INIT('h0155)
	) name8711 (
		_w8640_,
		_w8647_,
		_w8743_,
		_w8744_,
		_w8745_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8712 (
		_w2874_,
		_w4695_,
		_w6944_,
		_w6946_,
		_w8746_
	);
	LUT4 #(
		.INIT('h007d)
	) name8713 (
		_w2975_,
		_w6947_,
		_w6949_,
		_w8746_,
		_w8747_
	);
	LUT3 #(
		.INIT('h70)
	) name8714 (
		_w2986_,
		_w7032_,
		_w8747_,
		_w8748_
	);
	LUT4 #(
		.INIT('h95aa)
	) name8715 (
		\a[26] ,
		_w2875_,
		_w7882_,
		_w8748_,
		_w8749_
	);
	LUT4 #(
		.INIT('hf660)
	) name8716 (
		_w8407_,
		_w8411_,
		_w8745_,
		_w8749_,
		_w8750_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8717 (
		_w37_,
		_w7028_,
		_w7103_,
		_w7104_,
		_w8751_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8718 (
		_w3262_,
		_w3882_,
		_w6954_,
		_w6956_,
		_w8752_
	);
	LUT3 #(
		.INIT('h82)
	) name8719 (
		_w3214_,
		_w4030_,
		_w6952_,
		_w8753_
	);
	LUT3 #(
		.INIT('h07)
	) name8720 (
		_w3249_,
		_w7026_,
		_w8753_,
		_w8754_
	);
	LUT2 #(
		.INIT('h4)
	) name8721 (
		_w8752_,
		_w8754_,
		_w8755_
	);
	LUT3 #(
		.INIT('h9a)
	) name8722 (
		\a[23] ,
		_w8751_,
		_w8755_,
		_w8756_
	);
	LUT3 #(
		.INIT('hd4)
	) name8723 (
		_w8632_,
		_w8750_,
		_w8756_,
		_w8757_
	);
	LUT3 #(
		.INIT('h82)
	) name8724 (
		_w3312_,
		_w7111_,
		_w7113_,
		_w8758_
	);
	LUT3 #(
		.INIT('h82)
	) name8725 (
		_w3654_,
		_w6960_,
		_w6962_,
		_w8759_
	);
	LUT2 #(
		.INIT('h8)
	) name8726 (
		_w3311_,
		_w7020_,
		_w8760_
	);
	LUT4 #(
		.INIT('h4448)
	) name8727 (
		_w3409_,
		_w3645_,
		_w3650_,
		_w6959_,
		_w8761_
	);
	LUT2 #(
		.INIT('h1)
	) name8728 (
		_w8760_,
		_w8761_,
		_w8762_
	);
	LUT2 #(
		.INIT('h4)
	) name8729 (
		_w8759_,
		_w8762_,
		_w8763_
	);
	LUT3 #(
		.INIT('h9a)
	) name8730 (
		\a[20] ,
		_w8758_,
		_w8763_,
		_w8764_
	);
	LUT4 #(
		.INIT('hf660)
	) name8731 (
		_w8585_,
		_w8631_,
		_w8757_,
		_w8764_,
		_w8765_
	);
	LUT4 #(
		.INIT('hf660)
	) name8732 (
		_w8563_,
		_w8586_,
		_w8630_,
		_w8765_,
		_w8766_
	);
	LUT4 #(
		.INIT('h0069)
	) name8733 (
		_w8587_,
		_w8588_,
		_w8594_,
		_w8766_,
		_w8767_
	);
	LUT4 #(
		.INIT('h9600)
	) name8734 (
		_w8587_,
		_w8588_,
		_w8594_,
		_w8766_,
		_w8768_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8735 (
		_w3710_,
		_w7010_,
		_w7121_,
		_w7122_,
		_w8769_
	);
	LUT4 #(
		.INIT('h04c8)
	) name8736 (
		_w2983_,
		_w3886_,
		_w6972_,
		_w6974_,
		_w8770_
	);
	LUT3 #(
		.INIT('h82)
	) name8737 (
		_w3709_,
		_w6967_,
		_w6969_,
		_w8771_
	);
	LUT3 #(
		.INIT('h07)
	) name8738 (
		_w3877_,
		_w7008_,
		_w8771_,
		_w8772_
	);
	LUT2 #(
		.INIT('h4)
	) name8739 (
		_w8770_,
		_w8772_,
		_w8773_
	);
	LUT3 #(
		.INIT('h9a)
	) name8740 (
		\a[17] ,
		_w8769_,
		_w8773_,
		_w8774_
	);
	LUT3 #(
		.INIT('h54)
	) name8741 (
		_w8767_,
		_w8768_,
		_w8774_,
		_w8775_
	);
	LUT3 #(
		.INIT('h82)
	) name8742 (
		_w4034_,
		_w7129_,
		_w7131_,
		_w8776_
	);
	LUT3 #(
		.INIT('h84)
	) name8743 (
		_w2546_,
		_w4382_,
		_w6981_,
		_w8777_
	);
	LUT2 #(
		.INIT('h8)
	) name8744 (
		_w4033_,
		_w7002_,
		_w8778_
	);
	LUT4 #(
		.INIT('h04c8)
	) name8745 (
		_w2622_,
		_w4367_,
		_w6978_,
		_w6980_,
		_w8779_
	);
	LUT2 #(
		.INIT('h1)
	) name8746 (
		_w8778_,
		_w8779_,
		_w8780_
	);
	LUT2 #(
		.INIT('h4)
	) name8747 (
		_w8777_,
		_w8780_,
		_w8781_
	);
	LUT3 #(
		.INIT('h9a)
	) name8748 (
		\a[14] ,
		_w8776_,
		_w8781_,
		_w8782_
	);
	LUT3 #(
		.INIT('hd4)
	) name8749 (
		_w8626_,
		_w8775_,
		_w8782_,
		_w8783_
	);
	LUT3 #(
		.INIT('h54)
	) name8750 (
		_w8623_,
		_w8624_,
		_w8783_,
		_w8784_
	);
	LUT3 #(
		.INIT('h69)
	) name8751 (
		_w8604_,
		_w8605_,
		_w8611_,
		_w8785_
	);
	LUT4 #(
		.INIT('h0a02)
	) name8752 (
		_w4459_,
		_w7169_,
		_w7419_,
		_w7686_,
		_w8786_
	);
	LUT3 #(
		.INIT('h28)
	) name8753 (
		_w4458_,
		_w7136_,
		_w7168_,
		_w8787_
	);
	LUT3 #(
		.INIT('h40)
	) name8754 (
		_w4700_,
		_w7136_,
		_w7167_,
		_w8788_
	);
	LUT3 #(
		.INIT('h31)
	) name8755 (
		_w8545_,
		_w8787_,
		_w8788_,
		_w8789_
	);
	LUT3 #(
		.INIT('h9a)
	) name8756 (
		\a[11] ,
		_w8786_,
		_w8789_,
		_w8790_
	);
	LUT3 #(
		.INIT('hb2)
	) name8757 (
		_w8784_,
		_w8785_,
		_w8790_,
		_w8791_
	);
	LUT2 #(
		.INIT('h2)
	) name8758 (
		_w8618_,
		_w8791_,
		_w8792_
	);
	LUT2 #(
		.INIT('h4)
	) name8759 (
		_w8618_,
		_w8791_,
		_w8793_
	);
	LUT2 #(
		.INIT('h9)
	) name8760 (
		_w8618_,
		_w8791_,
		_w8794_
	);
	LUT3 #(
		.INIT('h28)
	) name8761 (
		_w4684_,
		_w7136_,
		_w7168_,
		_w8795_
	);
	LUT4 #(
		.INIT('h028a)
	) name8762 (
		_w4700_,
		_w7136_,
		_w7166_,
		_w7167_,
		_w8796_
	);
	LUT4 #(
		.INIT('h04c8)
	) name8763 (
		_w2411_,
		_w4458_,
		_w6983_,
		_w6993_,
		_w8797_
	);
	LUT3 #(
		.INIT('h01)
	) name8764 (
		_w8796_,
		_w8797_,
		_w8795_,
		_w8798_
	);
	LUT4 #(
		.INIT('h95aa)
	) name8765 (
		\a[11] ,
		_w4459_,
		_w7696_,
		_w8798_,
		_w8799_
	);
	LUT3 #(
		.INIT('h96)
	) name8766 (
		_w8626_,
		_w8775_,
		_w8782_,
		_w8800_
	);
	LUT4 #(
		.INIT('h9669)
	) name8767 (
		_w8563_,
		_w8586_,
		_w8630_,
		_w8765_,
		_w8801_
	);
	LUT4 #(
		.INIT('h04c8)
	) name8768 (
		_w3257_,
		_w3709_,
		_w6964_,
		_w6966_,
		_w8802_
	);
	LUT4 #(
		.INIT('h007d)
	) name8769 (
		_w3877_,
		_w6967_,
		_w6969_,
		_w8802_,
		_w8803_
	);
	LUT3 #(
		.INIT('h70)
	) name8770 (
		_w3886_,
		_w7008_,
		_w8803_,
		_w8804_
	);
	LUT4 #(
		.INIT('h95aa)
	) name8771 (
		\a[17] ,
		_w3710_,
		_w7403_,
		_w8804_,
		_w8805_
	);
	LUT4 #(
		.INIT('h9669)
	) name8772 (
		_w8585_,
		_w8631_,
		_w8757_,
		_w8764_,
		_w8806_
	);
	LUT3 #(
		.INIT('h1e)
	) name8773 (
		_w8647_,
		_w8743_,
		_w8744_,
		_w8807_
	);
	LUT3 #(
		.INIT('h82)
	) name8774 (
		_w2875_,
		_w7093_,
		_w7095_,
		_w8808_
	);
	LUT3 #(
		.INIT('h82)
	) name8775 (
		_w2986_,
		_w6947_,
		_w6949_,
		_w8809_
	);
	LUT2 #(
		.INIT('h8)
	) name8776 (
		_w2874_,
		_w7038_,
		_w8810_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8777 (
		_w2975_,
		_w4695_,
		_w6944_,
		_w6946_,
		_w8811_
	);
	LUT2 #(
		.INIT('h1)
	) name8778 (
		_w8810_,
		_w8811_,
		_w8812_
	);
	LUT2 #(
		.INIT('h4)
	) name8779 (
		_w8809_,
		_w8812_,
		_w8813_
	);
	LUT4 #(
		.INIT('h4844)
	) name8780 (
		\a[26] ,
		_w8807_,
		_w8808_,
		_w8813_,
		_w8814_
	);
	LUT4 #(
		.INIT('h54ab)
	) name8781 (
		_w8653_,
		_w8739_,
		_w8740_,
		_w8742_,
		_w8815_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8782 (
		_w2875_,
		_w7040_,
		_w7091_,
		_w7092_,
		_w8816_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8783 (
		_w2986_,
		_w4695_,
		_w6944_,
		_w6946_,
		_w8817_
	);
	LUT3 #(
		.INIT('h82)
	) name8784 (
		_w2874_,
		_w6940_,
		_w6942_,
		_w8818_
	);
	LUT3 #(
		.INIT('h07)
	) name8785 (
		_w2975_,
		_w7038_,
		_w8818_,
		_w8819_
	);
	LUT2 #(
		.INIT('h4)
	) name8786 (
		_w8817_,
		_w8819_,
		_w8820_
	);
	LUT4 #(
		.INIT('h4844)
	) name8787 (
		\a[26] ,
		_w8815_,
		_w8816_,
		_w8820_,
		_w8821_
	);
	LUT2 #(
		.INIT('h9)
	) name8788 (
		_w8739_,
		_w8741_,
		_w8822_
	);
	LUT4 #(
		.INIT('h2228)
	) name8789 (
		_w2874_,
		_w5067_,
		_w5282_,
		_w6939_,
		_w8823_
	);
	LUT4 #(
		.INIT('h007d)
	) name8790 (
		_w2975_,
		_w6940_,
		_w6942_,
		_w8823_,
		_w8824_
	);
	LUT3 #(
		.INIT('h70)
	) name8791 (
		_w2986_,
		_w7038_,
		_w8824_,
		_w8825_
	);
	LUT4 #(
		.INIT('h95aa)
	) name8792 (
		\a[26] ,
		_w2875_,
		_w8018_,
		_w8825_,
		_w8826_
	);
	LUT2 #(
		.INIT('h2)
	) name8793 (
		_w8822_,
		_w8826_,
		_w8827_
	);
	LUT3 #(
		.INIT('h1e)
	) name8794 (
		_w8668_,
		_w8737_,
		_w8738_,
		_w8828_
	);
	LUT3 #(
		.INIT('h82)
	) name8795 (
		_w2875_,
		_w7087_,
		_w7089_,
		_w8829_
	);
	LUT3 #(
		.INIT('h82)
	) name8796 (
		_w2986_,
		_w6940_,
		_w6942_,
		_w8830_
	);
	LUT2 #(
		.INIT('h8)
	) name8797 (
		_w2874_,
		_w7044_,
		_w8831_
	);
	LUT4 #(
		.INIT('h2228)
	) name8798 (
		_w2975_,
		_w5067_,
		_w5282_,
		_w6939_,
		_w8832_
	);
	LUT2 #(
		.INIT('h1)
	) name8799 (
		_w8831_,
		_w8832_,
		_w8833_
	);
	LUT2 #(
		.INIT('h4)
	) name8800 (
		_w8830_,
		_w8833_,
		_w8834_
	);
	LUT4 #(
		.INIT('h4844)
	) name8801 (
		\a[26] ,
		_w8828_,
		_w8829_,
		_w8834_,
		_w8835_
	);
	LUT4 #(
		.INIT('h54ab)
	) name8802 (
		_w8674_,
		_w8733_,
		_w8734_,
		_w8736_,
		_w8836_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8803 (
		_w2875_,
		_w7046_,
		_w7085_,
		_w7086_,
		_w8837_
	);
	LUT4 #(
		.INIT('h2228)
	) name8804 (
		_w2986_,
		_w5067_,
		_w5282_,
		_w6939_,
		_w8838_
	);
	LUT3 #(
		.INIT('h82)
	) name8805 (
		_w2874_,
		_w6935_,
		_w6937_,
		_w8839_
	);
	LUT3 #(
		.INIT('h07)
	) name8806 (
		_w2975_,
		_w7044_,
		_w8839_,
		_w8840_
	);
	LUT2 #(
		.INIT('h4)
	) name8807 (
		_w8838_,
		_w8840_,
		_w8841_
	);
	LUT4 #(
		.INIT('h4844)
	) name8808 (
		\a[26] ,
		_w8836_,
		_w8837_,
		_w8841_,
		_w8842_
	);
	LUT2 #(
		.INIT('h9)
	) name8809 (
		_w8733_,
		_w8735_,
		_w8843_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8810 (
		_w2874_,
		_w6043_,
		_w6933_,
		_w6934_,
		_w8844_
	);
	LUT4 #(
		.INIT('h007d)
	) name8811 (
		_w2975_,
		_w6935_,
		_w6937_,
		_w8844_,
		_w8845_
	);
	LUT3 #(
		.INIT('h70)
	) name8812 (
		_w2986_,
		_w7044_,
		_w8845_,
		_w8846_
	);
	LUT4 #(
		.INIT('h95aa)
	) name8813 (
		\a[26] ,
		_w2875_,
		_w8005_,
		_w8846_,
		_w8847_
	);
	LUT2 #(
		.INIT('h2)
	) name8814 (
		_w8843_,
		_w8847_,
		_w8848_
	);
	LUT3 #(
		.INIT('h1e)
	) name8815 (
		_w8689_,
		_w8731_,
		_w8732_,
		_w8849_
	);
	LUT3 #(
		.INIT('h82)
	) name8816 (
		_w2875_,
		_w7081_,
		_w7083_,
		_w8850_
	);
	LUT3 #(
		.INIT('h82)
	) name8817 (
		_w2986_,
		_w6935_,
		_w6937_,
		_w8851_
	);
	LUT2 #(
		.INIT('h8)
	) name8818 (
		_w2874_,
		_w7050_,
		_w8852_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8819 (
		_w2975_,
		_w6043_,
		_w6933_,
		_w6934_,
		_w8853_
	);
	LUT2 #(
		.INIT('h1)
	) name8820 (
		_w8852_,
		_w8853_,
		_w8854_
	);
	LUT2 #(
		.INIT('h4)
	) name8821 (
		_w8851_,
		_w8854_,
		_w8855_
	);
	LUT4 #(
		.INIT('h4844)
	) name8822 (
		\a[26] ,
		_w8849_,
		_w8850_,
		_w8855_,
		_w8856_
	);
	LUT4 #(
		.INIT('h54ab)
	) name8823 (
		_w8696_,
		_w8727_,
		_w8728_,
		_w8730_,
		_w8857_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8824 (
		_w2875_,
		_w7052_,
		_w7079_,
		_w7080_,
		_w8858_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8825 (
		_w2986_,
		_w6043_,
		_w6933_,
		_w6934_,
		_w8859_
	);
	LUT3 #(
		.INIT('h82)
	) name8826 (
		_w2874_,
		_w6929_,
		_w6931_,
		_w8860_
	);
	LUT3 #(
		.INIT('h07)
	) name8827 (
		_w2975_,
		_w7050_,
		_w8860_,
		_w8861_
	);
	LUT2 #(
		.INIT('h4)
	) name8828 (
		_w8859_,
		_w8861_,
		_w8862_
	);
	LUT4 #(
		.INIT('h4844)
	) name8829 (
		\a[26] ,
		_w8857_,
		_w8858_,
		_w8862_,
		_w8863_
	);
	LUT2 #(
		.INIT('h9)
	) name8830 (
		_w8727_,
		_w8729_,
		_w8864_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8831 (
		_w2874_,
		_w6645_,
		_w6926_,
		_w6928_,
		_w8865_
	);
	LUT4 #(
		.INIT('h007d)
	) name8832 (
		_w2975_,
		_w6929_,
		_w6931_,
		_w8865_,
		_w8866_
	);
	LUT3 #(
		.INIT('h70)
	) name8833 (
		_w2986_,
		_w7050_,
		_w8866_,
		_w8867_
	);
	LUT4 #(
		.INIT('h95aa)
	) name8834 (
		\a[26] ,
		_w2875_,
		_w8227_,
		_w8867_,
		_w8868_
	);
	LUT2 #(
		.INIT('h2)
	) name8835 (
		_w8864_,
		_w8868_,
		_w8869_
	);
	LUT3 #(
		.INIT('h82)
	) name8836 (
		_w2875_,
		_w7075_,
		_w7077_,
		_w8870_
	);
	LUT3 #(
		.INIT('h82)
	) name8837 (
		_w2986_,
		_w6929_,
		_w6931_,
		_w8871_
	);
	LUT2 #(
		.INIT('h8)
	) name8838 (
		_w2874_,
		_w7056_,
		_w8872_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8839 (
		_w2975_,
		_w6645_,
		_w6926_,
		_w6928_,
		_w8873_
	);
	LUT2 #(
		.INIT('h1)
	) name8840 (
		_w8872_,
		_w8873_,
		_w8874_
	);
	LUT2 #(
		.INIT('h4)
	) name8841 (
		_w8871_,
		_w8874_,
		_w8875_
	);
	LUT2 #(
		.INIT('h9)
	) name8842 (
		_w8724_,
		_w8726_,
		_w8876_
	);
	LUT4 #(
		.INIT('h6500)
	) name8843 (
		\a[26] ,
		_w8870_,
		_w8875_,
		_w8876_,
		_w8877_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8844 (
		_w2875_,
		_w7058_,
		_w7073_,
		_w7074_,
		_w8878_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8845 (
		_w2986_,
		_w6645_,
		_w6926_,
		_w6928_,
		_w8879_
	);
	LUT3 #(
		.INIT('h82)
	) name8846 (
		_w2874_,
		_w6922_,
		_w6924_,
		_w8880_
	);
	LUT3 #(
		.INIT('h07)
	) name8847 (
		_w2975_,
		_w7056_,
		_w8880_,
		_w8881_
	);
	LUT2 #(
		.INIT('h4)
	) name8848 (
		_w8879_,
		_w8881_,
		_w8882_
	);
	LUT4 #(
		.INIT('h9a65)
	) name8849 (
		\a[29] ,
		_w8717_,
		_w8721_,
		_w8722_,
		_w8883_
	);
	LUT4 #(
		.INIT('h6500)
	) name8850 (
		\a[26] ,
		_w8878_,
		_w8882_,
		_w8883_,
		_w8884_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8851 (
		_w2874_,
		_w6669_,
		_w6919_,
		_w6921_,
		_w8885_
	);
	LUT4 #(
		.INIT('h007d)
	) name8852 (
		_w2975_,
		_w6922_,
		_w6924_,
		_w8885_,
		_w8886_
	);
	LUT3 #(
		.INIT('h70)
	) name8853 (
		_w2986_,
		_w7056_,
		_w8886_,
		_w8887_
	);
	LUT4 #(
		.INIT('h95aa)
	) name8854 (
		\a[26] ,
		_w2875_,
		_w8298_,
		_w8887_,
		_w8888_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name8855 (
		\a[29] ,
		_w8709_,
		_w8706_,
		_w8708_,
		_w8889_
	);
	LUT3 #(
		.INIT('h4b)
	) name8856 (
		_w8712_,
		_w8715_,
		_w8889_,
		_w8890_
	);
	LUT2 #(
		.INIT('h4)
	) name8857 (
		_w8888_,
		_w8890_,
		_w8891_
	);
	LUT3 #(
		.INIT('h82)
	) name8858 (
		_w2875_,
		_w7069_,
		_w7071_,
		_w8892_
	);
	LUT3 #(
		.INIT('h82)
	) name8859 (
		_w2986_,
		_w6922_,
		_w6924_,
		_w8893_
	);
	LUT2 #(
		.INIT('h8)
	) name8860 (
		_w2874_,
		_w7062_,
		_w8894_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8861 (
		_w2975_,
		_w6669_,
		_w6919_,
		_w6921_,
		_w8895_
	);
	LUT2 #(
		.INIT('h1)
	) name8862 (
		_w8894_,
		_w8895_,
		_w8896_
	);
	LUT2 #(
		.INIT('h4)
	) name8863 (
		_w8893_,
		_w8896_,
		_w8897_
	);
	LUT2 #(
		.INIT('h8)
	) name8864 (
		\a[29] ,
		_w8709_,
		_w8898_
	);
	LUT3 #(
		.INIT('h4b)
	) name8865 (
		_w8706_,
		_w8708_,
		_w8898_,
		_w8899_
	);
	LUT4 #(
		.INIT('h6500)
	) name8866 (
		\a[26] ,
		_w8892_,
		_w8897_,
		_w8899_,
		_w8900_
	);
	LUT4 #(
		.INIT('h2882)
	) name8867 (
		_w2875_,
		_w6914_,
		_w6916_,
		_w7067_,
		_w8901_
	);
	LUT4 #(
		.INIT('ha802)
	) name8868 (
		_w2975_,
		_w6689_,
		_w6911_,
		_w6913_,
		_w8902_
	);
	LUT4 #(
		.INIT('h007d)
	) name8869 (
		_w2986_,
		_w6914_,
		_w6916_,
		_w8902_,
		_w8903_
	);
	LUT4 #(
		.INIT('h5401)
	) name8870 (
		_w2873_,
		_w6689_,
		_w6911_,
		_w6913_,
		_w8904_
	);
	LUT2 #(
		.INIT('h2)
	) name8871 (
		\a[26] ,
		_w8904_,
		_w8905_
	);
	LUT3 #(
		.INIT('h40)
	) name8872 (
		_w8901_,
		_w8903_,
		_w8905_,
		_w8906_
	);
	LUT3 #(
		.INIT('h28)
	) name8873 (
		_w2875_,
		_w7062_,
		_w8358_,
		_w8907_
	);
	LUT4 #(
		.INIT('ha802)
	) name8874 (
		_w2874_,
		_w6689_,
		_w6911_,
		_w6913_,
		_w8908_
	);
	LUT4 #(
		.INIT('h007d)
	) name8875 (
		_w2975_,
		_w6914_,
		_w6916_,
		_w8908_,
		_w8909_
	);
	LUT3 #(
		.INIT('h70)
	) name8876 (
		_w2986_,
		_w7062_,
		_w8909_,
		_w8910_
	);
	LUT4 #(
		.INIT('h0800)
	) name8877 (
		_w8709_,
		_w8906_,
		_w8907_,
		_w8910_,
		_w8911_
	);
	LUT3 #(
		.INIT('h28)
	) name8878 (
		_w2875_,
		_w7065_,
		_w7068_,
		_w8912_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8879 (
		_w2986_,
		_w6669_,
		_w6919_,
		_w6921_,
		_w8913_
	);
	LUT3 #(
		.INIT('h82)
	) name8880 (
		_w2874_,
		_w6914_,
		_w6916_,
		_w8914_
	);
	LUT3 #(
		.INIT('h07)
	) name8881 (
		_w2975_,
		_w7062_,
		_w8914_,
		_w8915_
	);
	LUT2 #(
		.INIT('h4)
	) name8882 (
		_w8913_,
		_w8915_,
		_w8916_
	);
	LUT4 #(
		.INIT('ha6aa)
	) name8883 (
		_w8709_,
		_w8906_,
		_w8907_,
		_w8910_,
		_w8917_
	);
	LUT4 #(
		.INIT('h6500)
	) name8884 (
		\a[26] ,
		_w8912_,
		_w8916_,
		_w8917_,
		_w8918_
	);
	LUT2 #(
		.INIT('h1)
	) name8885 (
		_w8911_,
		_w8918_,
		_w8919_
	);
	LUT4 #(
		.INIT('h009a)
	) name8886 (
		\a[26] ,
		_w8892_,
		_w8897_,
		_w8899_,
		_w8920_
	);
	LUT4 #(
		.INIT('h9a65)
	) name8887 (
		\a[26] ,
		_w8892_,
		_w8897_,
		_w8899_,
		_w8921_
	);
	LUT3 #(
		.INIT('h54)
	) name8888 (
		_w8900_,
		_w8919_,
		_w8920_,
		_w8922_
	);
	LUT2 #(
		.INIT('h2)
	) name8889 (
		_w8888_,
		_w8890_,
		_w8923_
	);
	LUT2 #(
		.INIT('h9)
	) name8890 (
		_w8888_,
		_w8890_,
		_w8924_
	);
	LUT4 #(
		.INIT('h9a65)
	) name8891 (
		\a[26] ,
		_w8878_,
		_w8882_,
		_w8883_,
		_w8925_
	);
	LUT4 #(
		.INIT('h4d00)
	) name8892 (
		_w8888_,
		_w8890_,
		_w8922_,
		_w8925_,
		_w8926_
	);
	LUT4 #(
		.INIT('h9a65)
	) name8893 (
		\a[26] ,
		_w8870_,
		_w8875_,
		_w8876_,
		_w8927_
	);
	LUT4 #(
		.INIT('h0155)
	) name8894 (
		_w8877_,
		_w8884_,
		_w8926_,
		_w8927_,
		_w8928_
	);
	LUT2 #(
		.INIT('h4)
	) name8895 (
		_w8864_,
		_w8868_,
		_w8929_
	);
	LUT2 #(
		.INIT('h9)
	) name8896 (
		_w8864_,
		_w8868_,
		_w8930_
	);
	LUT4 #(
		.INIT('h9699)
	) name8897 (
		\a[26] ,
		_w8857_,
		_w8858_,
		_w8862_,
		_w8931_
	);
	LUT4 #(
		.INIT('h2b00)
	) name8898 (
		_w8864_,
		_w8868_,
		_w8928_,
		_w8931_,
		_w8932_
	);
	LUT4 #(
		.INIT('h9699)
	) name8899 (
		\a[26] ,
		_w8849_,
		_w8850_,
		_w8855_,
		_w8933_
	);
	LUT4 #(
		.INIT('h0155)
	) name8900 (
		_w8856_,
		_w8863_,
		_w8932_,
		_w8933_,
		_w8934_
	);
	LUT2 #(
		.INIT('h4)
	) name8901 (
		_w8843_,
		_w8847_,
		_w8935_
	);
	LUT2 #(
		.INIT('h9)
	) name8902 (
		_w8843_,
		_w8847_,
		_w8936_
	);
	LUT4 #(
		.INIT('h9699)
	) name8903 (
		\a[26] ,
		_w8836_,
		_w8837_,
		_w8841_,
		_w8937_
	);
	LUT4 #(
		.INIT('h2b00)
	) name8904 (
		_w8843_,
		_w8847_,
		_w8934_,
		_w8937_,
		_w8938_
	);
	LUT4 #(
		.INIT('h9699)
	) name8905 (
		\a[26] ,
		_w8828_,
		_w8829_,
		_w8834_,
		_w8939_
	);
	LUT4 #(
		.INIT('h0155)
	) name8906 (
		_w8835_,
		_w8842_,
		_w8938_,
		_w8939_,
		_w8940_
	);
	LUT2 #(
		.INIT('h4)
	) name8907 (
		_w8822_,
		_w8826_,
		_w8941_
	);
	LUT2 #(
		.INIT('h9)
	) name8908 (
		_w8822_,
		_w8826_,
		_w8942_
	);
	LUT4 #(
		.INIT('h9699)
	) name8909 (
		\a[26] ,
		_w8815_,
		_w8816_,
		_w8820_,
		_w8943_
	);
	LUT4 #(
		.INIT('h2b00)
	) name8910 (
		_w8822_,
		_w8826_,
		_w8940_,
		_w8943_,
		_w8944_
	);
	LUT4 #(
		.INIT('h9699)
	) name8911 (
		\a[26] ,
		_w8807_,
		_w8808_,
		_w8813_,
		_w8945_
	);
	LUT4 #(
		.INIT('h0155)
	) name8912 (
		_w8814_,
		_w8821_,
		_w8944_,
		_w8945_,
		_w8946_
	);
	LUT4 #(
		.INIT('h9669)
	) name8913 (
		_w8407_,
		_w8411_,
		_w8745_,
		_w8749_,
		_w8947_
	);
	LUT4 #(
		.INIT('h2228)
	) name8914 (
		_w3214_,
		_w4099_,
		_w4378_,
		_w6951_,
		_w8948_
	);
	LUT4 #(
		.INIT('h007d)
	) name8915 (
		_w3249_,
		_w4030_,
		_w6952_,
		_w8948_,
		_w8949_
	);
	LUT3 #(
		.INIT('h70)
	) name8916 (
		_w3262_,
		_w7026_,
		_w8949_,
		_w8950_
	);
	LUT4 #(
		.INIT('h95aa)
	) name8917 (
		\a[23] ,
		_w37_,
		_w7562_,
		_w8950_,
		_w8951_
	);
	LUT3 #(
		.INIT('hb2)
	) name8918 (
		_w8946_,
		_w8947_,
		_w8951_,
		_w8952_
	);
	LUT4 #(
		.INIT('h0096)
	) name8919 (
		_w8632_,
		_w8750_,
		_w8756_,
		_w8952_,
		_w8953_
	);
	LUT4 #(
		.INIT('h6900)
	) name8920 (
		_w8632_,
		_w8750_,
		_w8756_,
		_w8952_,
		_w8954_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8921 (
		_w3312_,
		_w7022_,
		_w7109_,
		_w7110_,
		_w8955_
	);
	LUT4 #(
		.INIT('h5060)
	) name8922 (
		_w3409_,
		_w3650_,
		_w3654_,
		_w6959_,
		_w8956_
	);
	LUT3 #(
		.INIT('h82)
	) name8923 (
		_w3311_,
		_w3706_,
		_w6957_,
		_w8957_
	);
	LUT3 #(
		.INIT('h07)
	) name8924 (
		_w3645_,
		_w7020_,
		_w8957_,
		_w8958_
	);
	LUT2 #(
		.INIT('h4)
	) name8925 (
		_w8956_,
		_w8958_,
		_w8959_
	);
	LUT3 #(
		.INIT('h9a)
	) name8926 (
		\a[20] ,
		_w8955_,
		_w8959_,
		_w8960_
	);
	LUT3 #(
		.INIT('h54)
	) name8927 (
		_w8953_,
		_w8954_,
		_w8960_,
		_w8961_
	);
	LUT3 #(
		.INIT('h82)
	) name8928 (
		_w3710_,
		_w7117_,
		_w7119_,
		_w8962_
	);
	LUT3 #(
		.INIT('h82)
	) name8929 (
		_w3886_,
		_w6967_,
		_w6969_,
		_w8963_
	);
	LUT2 #(
		.INIT('h8)
	) name8930 (
		_w3709_,
		_w7014_,
		_w8964_
	);
	LUT4 #(
		.INIT('h04c8)
	) name8931 (
		_w3257_,
		_w3877_,
		_w6964_,
		_w6966_,
		_w8965_
	);
	LUT2 #(
		.INIT('h1)
	) name8932 (
		_w8964_,
		_w8965_,
		_w8966_
	);
	LUT2 #(
		.INIT('h4)
	) name8933 (
		_w8963_,
		_w8966_,
		_w8967_
	);
	LUT3 #(
		.INIT('h9a)
	) name8934 (
		\a[17] ,
		_w8962_,
		_w8967_,
		_w8968_
	);
	LUT3 #(
		.INIT('hd4)
	) name8935 (
		_w8806_,
		_w8961_,
		_w8968_,
		_w8969_
	);
	LUT3 #(
		.INIT('hd4)
	) name8936 (
		_w8801_,
		_w8805_,
		_w8969_,
		_w8970_
	);
	LUT4 #(
		.INIT('h6996)
	) name8937 (
		_w8587_,
		_w8588_,
		_w8594_,
		_w8766_,
		_w8971_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8938 (
		_w4034_,
		_w7004_,
		_w7127_,
		_w7128_,
		_w8972_
	);
	LUT4 #(
		.INIT('h04c8)
	) name8939 (
		_w2622_,
		_w4382_,
		_w6978_,
		_w6980_,
		_w8973_
	);
	LUT3 #(
		.INIT('h84)
	) name8940 (
		_w2872_,
		_w4033_,
		_w6975_,
		_w8974_
	);
	LUT3 #(
		.INIT('h07)
	) name8941 (
		_w4367_,
		_w7002_,
		_w8974_,
		_w8975_
	);
	LUT2 #(
		.INIT('h4)
	) name8942 (
		_w8973_,
		_w8975_,
		_w8976_
	);
	LUT3 #(
		.INIT('h9a)
	) name8943 (
		\a[14] ,
		_w8972_,
		_w8976_,
		_w8977_
	);
	LUT4 #(
		.INIT('hde48)
	) name8944 (
		_w8774_,
		_w8970_,
		_w8971_,
		_w8977_,
		_w8978_
	);
	LUT4 #(
		.INIT('h0096)
	) name8945 (
		_w8626_,
		_w8775_,
		_w8782_,
		_w8978_,
		_w8979_
	);
	LUT4 #(
		.INIT('h6900)
	) name8946 (
		_w8626_,
		_w8775_,
		_w8782_,
		_w8978_,
		_w8980_
	);
	LUT3 #(
		.INIT('h82)
	) name8947 (
		_w4459_,
		_w7135_,
		_w7172_,
		_w8981_
	);
	LUT3 #(
		.INIT('h28)
	) name8948 (
		_w4700_,
		_w7136_,
		_w7168_,
		_w8982_
	);
	LUT2 #(
		.INIT('h8)
	) name8949 (
		_w4458_,
		_w6996_,
		_w8983_
	);
	LUT4 #(
		.INIT('h04c8)
	) name8950 (
		_w2411_,
		_w4684_,
		_w6983_,
		_w6993_,
		_w8984_
	);
	LUT2 #(
		.INIT('h1)
	) name8951 (
		_w8983_,
		_w8984_,
		_w8985_
	);
	LUT2 #(
		.INIT('h4)
	) name8952 (
		_w8982_,
		_w8985_,
		_w8986_
	);
	LUT3 #(
		.INIT('h9a)
	) name8953 (
		\a[11] ,
		_w8981_,
		_w8986_,
		_w8987_
	);
	LUT4 #(
		.INIT('h0445)
	) name8954 (
		_w8799_,
		_w8800_,
		_w8978_,
		_w8987_,
		_w8988_
	);
	LUT2 #(
		.INIT('h9)
	) name8955 (
		_w8625_,
		_w8783_,
		_w8989_
	);
	LUT4 #(
		.INIT('ha220)
	) name8956 (
		_w8799_,
		_w8800_,
		_w8978_,
		_w8987_,
		_w8990_
	);
	LUT4 #(
		.INIT('h999a)
	) name8957 (
		_w8799_,
		_w8979_,
		_w8980_,
		_w8987_,
		_w8991_
	);
	LUT3 #(
		.INIT('h51)
	) name8958 (
		_w8988_,
		_w8989_,
		_w8990_,
		_w8992_
	);
	LUT3 #(
		.INIT('h69)
	) name8959 (
		_w8784_,
		_w8785_,
		_w8790_,
		_w8993_
	);
	LUT2 #(
		.INIT('h1)
	) name8960 (
		_w8992_,
		_w8993_,
		_w8994_
	);
	LUT4 #(
		.INIT('h028a)
	) name8961 (
		_w4875_,
		_w7136_,
		_w7166_,
		_w7167_,
		_w8995_
	);
	LUT4 #(
		.INIT('h781e)
	) name8962 (
		\a[5] ,
		\a[6] ,
		\a[7] ,
		\a[8] ,
		_w8996_
	);
	LUT3 #(
		.INIT('hb0)
	) name8963 (
		_w7136_,
		_w7166_,
		_w8996_,
		_w8997_
	);
	LUT2 #(
		.INIT('h1)
	) name8964 (
		_w8995_,
		_w8997_,
		_w8998_
	);
	LUT4 #(
		.INIT('h5700)
	) name8965 (
		_w4876_,
		_w7418_,
		_w7419_,
		_w8998_,
		_w8999_
	);
	LUT2 #(
		.INIT('h6)
	) name8966 (
		\a[8] ,
		_w8999_,
		_w9000_
	);
	LUT4 #(
		.INIT('h04c8)
	) name8967 (
		_w2983_,
		_w4033_,
		_w6972_,
		_w6974_,
		_w9001_
	);
	LUT4 #(
		.INIT('h007b)
	) name8968 (
		_w2872_,
		_w4367_,
		_w6975_,
		_w9001_,
		_w9002_
	);
	LUT3 #(
		.INIT('h70)
	) name8969 (
		_w4382_,
		_w7002_,
		_w9002_,
		_w9003_
	);
	LUT4 #(
		.INIT('h95aa)
	) name8970 (
		\a[14] ,
		_w4034_,
		_w7426_,
		_w9003_,
		_w9004_
	);
	LUT4 #(
		.INIT('h0096)
	) name8971 (
		_w8801_,
		_w8805_,
		_w8969_,
		_w9004_,
		_w9005_
	);
	LUT4 #(
		.INIT('h6900)
	) name8972 (
		_w8801_,
		_w8805_,
		_w8969_,
		_w9004_,
		_w9006_
	);
	LUT4 #(
		.INIT('h9669)
	) name8973 (
		_w8801_,
		_w8805_,
		_w8969_,
		_w9004_,
		_w9007_
	);
	LUT4 #(
		.INIT('h9669)
	) name8974 (
		_w8632_,
		_w8750_,
		_w8756_,
		_w8952_,
		_w9008_
	);
	LUT3 #(
		.INIT('h82)
	) name8975 (
		_w37_,
		_w7099_,
		_w7101_,
		_w9009_
	);
	LUT3 #(
		.INIT('h82)
	) name8976 (
		_w3262_,
		_w4030_,
		_w6952_,
		_w9010_
	);
	LUT2 #(
		.INIT('h8)
	) name8977 (
		_w3214_,
		_w7032_,
		_w9011_
	);
	LUT4 #(
		.INIT('h2228)
	) name8978 (
		_w3249_,
		_w4099_,
		_w4378_,
		_w6951_,
		_w9012_
	);
	LUT2 #(
		.INIT('h1)
	) name8979 (
		_w9011_,
		_w9012_,
		_w9013_
	);
	LUT2 #(
		.INIT('h4)
	) name8980 (
		_w9010_,
		_w9013_,
		_w9014_
	);
	LUT3 #(
		.INIT('h1e)
	) name8981 (
		_w8821_,
		_w8944_,
		_w8945_,
		_w9015_
	);
	LUT4 #(
		.INIT('h6500)
	) name8982 (
		\a[23] ,
		_w9009_,
		_w9014_,
		_w9015_,
		_w9016_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8983 (
		_w37_,
		_w7034_,
		_w7097_,
		_w7098_,
		_w9017_
	);
	LUT4 #(
		.INIT('h2228)
	) name8984 (
		_w3262_,
		_w4099_,
		_w4378_,
		_w6951_,
		_w9018_
	);
	LUT3 #(
		.INIT('h82)
	) name8985 (
		_w3214_,
		_w6947_,
		_w6949_,
		_w9019_
	);
	LUT3 #(
		.INIT('h07)
	) name8986 (
		_w3249_,
		_w7032_,
		_w9019_,
		_w9020_
	);
	LUT2 #(
		.INIT('h4)
	) name8987 (
		_w9018_,
		_w9020_,
		_w9021_
	);
	LUT4 #(
		.INIT('h54ab)
	) name8988 (
		_w8827_,
		_w8940_,
		_w8941_,
		_w8943_,
		_w9022_
	);
	LUT4 #(
		.INIT('h6500)
	) name8989 (
		\a[23] ,
		_w9017_,
		_w9021_,
		_w9022_,
		_w9023_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8990 (
		_w3214_,
		_w4695_,
		_w6944_,
		_w6946_,
		_w9024_
	);
	LUT4 #(
		.INIT('h007d)
	) name8991 (
		_w3249_,
		_w6947_,
		_w6949_,
		_w9024_,
		_w9025_
	);
	LUT3 #(
		.INIT('h70)
	) name8992 (
		_w3262_,
		_w7032_,
		_w9025_,
		_w9026_
	);
	LUT4 #(
		.INIT('h95aa)
	) name8993 (
		\a[23] ,
		_w37_,
		_w7882_,
		_w9026_,
		_w9027_
	);
	LUT2 #(
		.INIT('h9)
	) name8994 (
		_w8940_,
		_w8942_,
		_w9028_
	);
	LUT2 #(
		.INIT('h4)
	) name8995 (
		_w9027_,
		_w9028_,
		_w9029_
	);
	LUT3 #(
		.INIT('h82)
	) name8996 (
		_w37_,
		_w7093_,
		_w7095_,
		_w9030_
	);
	LUT3 #(
		.INIT('h82)
	) name8997 (
		_w3262_,
		_w6947_,
		_w6949_,
		_w9031_
	);
	LUT2 #(
		.INIT('h8)
	) name8998 (
		_w3214_,
		_w7038_,
		_w9032_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8999 (
		_w3249_,
		_w4695_,
		_w6944_,
		_w6946_,
		_w9033_
	);
	LUT2 #(
		.INIT('h1)
	) name9000 (
		_w9032_,
		_w9033_,
		_w9034_
	);
	LUT2 #(
		.INIT('h4)
	) name9001 (
		_w9031_,
		_w9034_,
		_w9035_
	);
	LUT3 #(
		.INIT('h1e)
	) name9002 (
		_w8842_,
		_w8938_,
		_w8939_,
		_w9036_
	);
	LUT4 #(
		.INIT('h6500)
	) name9003 (
		\a[23] ,
		_w9030_,
		_w9035_,
		_w9036_,
		_w9037_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9004 (
		_w37_,
		_w7040_,
		_w7091_,
		_w7092_,
		_w9038_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9005 (
		_w3262_,
		_w4695_,
		_w6944_,
		_w6946_,
		_w9039_
	);
	LUT3 #(
		.INIT('h82)
	) name9006 (
		_w3214_,
		_w6940_,
		_w6942_,
		_w9040_
	);
	LUT3 #(
		.INIT('h07)
	) name9007 (
		_w3249_,
		_w7038_,
		_w9040_,
		_w9041_
	);
	LUT2 #(
		.INIT('h4)
	) name9008 (
		_w9039_,
		_w9041_,
		_w9042_
	);
	LUT4 #(
		.INIT('h54ab)
	) name9009 (
		_w8848_,
		_w8934_,
		_w8935_,
		_w8937_,
		_w9043_
	);
	LUT4 #(
		.INIT('h6500)
	) name9010 (
		\a[23] ,
		_w9038_,
		_w9042_,
		_w9043_,
		_w9044_
	);
	LUT4 #(
		.INIT('h2228)
	) name9011 (
		_w3214_,
		_w5067_,
		_w5282_,
		_w6939_,
		_w9045_
	);
	LUT4 #(
		.INIT('h007d)
	) name9012 (
		_w3249_,
		_w6940_,
		_w6942_,
		_w9045_,
		_w9046_
	);
	LUT3 #(
		.INIT('h70)
	) name9013 (
		_w3262_,
		_w7038_,
		_w9046_,
		_w9047_
	);
	LUT4 #(
		.INIT('h95aa)
	) name9014 (
		\a[23] ,
		_w37_,
		_w8018_,
		_w9047_,
		_w9048_
	);
	LUT2 #(
		.INIT('h9)
	) name9015 (
		_w8934_,
		_w8936_,
		_w9049_
	);
	LUT2 #(
		.INIT('h4)
	) name9016 (
		_w9048_,
		_w9049_,
		_w9050_
	);
	LUT3 #(
		.INIT('h82)
	) name9017 (
		_w37_,
		_w7087_,
		_w7089_,
		_w9051_
	);
	LUT3 #(
		.INIT('h82)
	) name9018 (
		_w3262_,
		_w6940_,
		_w6942_,
		_w9052_
	);
	LUT2 #(
		.INIT('h8)
	) name9019 (
		_w3214_,
		_w7044_,
		_w9053_
	);
	LUT4 #(
		.INIT('h2228)
	) name9020 (
		_w3249_,
		_w5067_,
		_w5282_,
		_w6939_,
		_w9054_
	);
	LUT2 #(
		.INIT('h1)
	) name9021 (
		_w9053_,
		_w9054_,
		_w9055_
	);
	LUT2 #(
		.INIT('h4)
	) name9022 (
		_w9052_,
		_w9055_,
		_w9056_
	);
	LUT3 #(
		.INIT('h1e)
	) name9023 (
		_w8863_,
		_w8932_,
		_w8933_,
		_w9057_
	);
	LUT4 #(
		.INIT('h6500)
	) name9024 (
		\a[23] ,
		_w9051_,
		_w9056_,
		_w9057_,
		_w9058_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9025 (
		_w37_,
		_w7046_,
		_w7085_,
		_w7086_,
		_w9059_
	);
	LUT4 #(
		.INIT('h2228)
	) name9026 (
		_w3262_,
		_w5067_,
		_w5282_,
		_w6939_,
		_w9060_
	);
	LUT3 #(
		.INIT('h82)
	) name9027 (
		_w3214_,
		_w6935_,
		_w6937_,
		_w9061_
	);
	LUT3 #(
		.INIT('h07)
	) name9028 (
		_w3249_,
		_w7044_,
		_w9061_,
		_w9062_
	);
	LUT2 #(
		.INIT('h4)
	) name9029 (
		_w9060_,
		_w9062_,
		_w9063_
	);
	LUT4 #(
		.INIT('h54ab)
	) name9030 (
		_w8869_,
		_w8928_,
		_w8929_,
		_w8931_,
		_w9064_
	);
	LUT4 #(
		.INIT('h6500)
	) name9031 (
		\a[23] ,
		_w9059_,
		_w9063_,
		_w9064_,
		_w9065_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9032 (
		_w3214_,
		_w6043_,
		_w6933_,
		_w6934_,
		_w9066_
	);
	LUT4 #(
		.INIT('h007d)
	) name9033 (
		_w3249_,
		_w6935_,
		_w6937_,
		_w9066_,
		_w9067_
	);
	LUT3 #(
		.INIT('h70)
	) name9034 (
		_w3262_,
		_w7044_,
		_w9067_,
		_w9068_
	);
	LUT4 #(
		.INIT('h95aa)
	) name9035 (
		\a[23] ,
		_w37_,
		_w8005_,
		_w9068_,
		_w9069_
	);
	LUT2 #(
		.INIT('h9)
	) name9036 (
		_w8928_,
		_w8930_,
		_w9070_
	);
	LUT2 #(
		.INIT('h4)
	) name9037 (
		_w9069_,
		_w9070_,
		_w9071_
	);
	LUT3 #(
		.INIT('h82)
	) name9038 (
		_w37_,
		_w7081_,
		_w7083_,
		_w9072_
	);
	LUT3 #(
		.INIT('h82)
	) name9039 (
		_w3262_,
		_w6935_,
		_w6937_,
		_w9073_
	);
	LUT2 #(
		.INIT('h8)
	) name9040 (
		_w3214_,
		_w7050_,
		_w9074_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9041 (
		_w3249_,
		_w6043_,
		_w6933_,
		_w6934_,
		_w9075_
	);
	LUT2 #(
		.INIT('h1)
	) name9042 (
		_w9074_,
		_w9075_,
		_w9076_
	);
	LUT2 #(
		.INIT('h4)
	) name9043 (
		_w9073_,
		_w9076_,
		_w9077_
	);
	LUT3 #(
		.INIT('h1e)
	) name9044 (
		_w8884_,
		_w8926_,
		_w8927_,
		_w9078_
	);
	LUT4 #(
		.INIT('h6500)
	) name9045 (
		\a[23] ,
		_w9072_,
		_w9077_,
		_w9078_,
		_w9079_
	);
	LUT4 #(
		.INIT('h54ab)
	) name9046 (
		_w8891_,
		_w8922_,
		_w8923_,
		_w8925_,
		_w9080_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9047 (
		_w37_,
		_w7052_,
		_w7079_,
		_w7080_,
		_w9081_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9048 (
		_w3262_,
		_w6043_,
		_w6933_,
		_w6934_,
		_w9082_
	);
	LUT3 #(
		.INIT('h82)
	) name9049 (
		_w3214_,
		_w6929_,
		_w6931_,
		_w9083_
	);
	LUT3 #(
		.INIT('h07)
	) name9050 (
		_w3249_,
		_w7050_,
		_w9083_,
		_w9084_
	);
	LUT2 #(
		.INIT('h4)
	) name9051 (
		_w9082_,
		_w9084_,
		_w9085_
	);
	LUT4 #(
		.INIT('h4844)
	) name9052 (
		\a[23] ,
		_w9080_,
		_w9081_,
		_w9085_,
		_w9086_
	);
	LUT2 #(
		.INIT('h9)
	) name9053 (
		_w8922_,
		_w8924_,
		_w9087_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9054 (
		_w3214_,
		_w6645_,
		_w6926_,
		_w6928_,
		_w9088_
	);
	LUT4 #(
		.INIT('h007d)
	) name9055 (
		_w3249_,
		_w6929_,
		_w6931_,
		_w9088_,
		_w9089_
	);
	LUT3 #(
		.INIT('h70)
	) name9056 (
		_w3262_,
		_w7050_,
		_w9089_,
		_w9090_
	);
	LUT4 #(
		.INIT('h95aa)
	) name9057 (
		\a[23] ,
		_w37_,
		_w8227_,
		_w9090_,
		_w9091_
	);
	LUT2 #(
		.INIT('h2)
	) name9058 (
		_w9087_,
		_w9091_,
		_w9092_
	);
	LUT3 #(
		.INIT('h82)
	) name9059 (
		_w37_,
		_w7075_,
		_w7077_,
		_w9093_
	);
	LUT3 #(
		.INIT('h82)
	) name9060 (
		_w3262_,
		_w6929_,
		_w6931_,
		_w9094_
	);
	LUT2 #(
		.INIT('h8)
	) name9061 (
		_w3214_,
		_w7056_,
		_w9095_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9062 (
		_w3249_,
		_w6645_,
		_w6926_,
		_w6928_,
		_w9096_
	);
	LUT2 #(
		.INIT('h1)
	) name9063 (
		_w9095_,
		_w9096_,
		_w9097_
	);
	LUT2 #(
		.INIT('h4)
	) name9064 (
		_w9094_,
		_w9097_,
		_w9098_
	);
	LUT2 #(
		.INIT('h9)
	) name9065 (
		_w8919_,
		_w8921_,
		_w9099_
	);
	LUT4 #(
		.INIT('h6500)
	) name9066 (
		\a[23] ,
		_w9093_,
		_w9098_,
		_w9099_,
		_w9100_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9067 (
		_w37_,
		_w7058_,
		_w7073_,
		_w7074_,
		_w9101_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9068 (
		_w3262_,
		_w6645_,
		_w6926_,
		_w6928_,
		_w9102_
	);
	LUT3 #(
		.INIT('h82)
	) name9069 (
		_w3214_,
		_w6922_,
		_w6924_,
		_w9103_
	);
	LUT3 #(
		.INIT('h07)
	) name9070 (
		_w3249_,
		_w7056_,
		_w9103_,
		_w9104_
	);
	LUT2 #(
		.INIT('h4)
	) name9071 (
		_w9102_,
		_w9104_,
		_w9105_
	);
	LUT4 #(
		.INIT('h9a65)
	) name9072 (
		\a[26] ,
		_w8912_,
		_w8916_,
		_w8917_,
		_w9106_
	);
	LUT4 #(
		.INIT('h6500)
	) name9073 (
		\a[23] ,
		_w9101_,
		_w9105_,
		_w9106_,
		_w9107_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9074 (
		_w3214_,
		_w6669_,
		_w6919_,
		_w6921_,
		_w9108_
	);
	LUT4 #(
		.INIT('h007d)
	) name9075 (
		_w3249_,
		_w6922_,
		_w6924_,
		_w9108_,
		_w9109_
	);
	LUT3 #(
		.INIT('h70)
	) name9076 (
		_w3262_,
		_w7056_,
		_w9109_,
		_w9110_
	);
	LUT4 #(
		.INIT('h95aa)
	) name9077 (
		\a[23] ,
		_w37_,
		_w8298_,
		_w9110_,
		_w9111_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name9078 (
		\a[26] ,
		_w8904_,
		_w8901_,
		_w8903_,
		_w9112_
	);
	LUT3 #(
		.INIT('h4b)
	) name9079 (
		_w8907_,
		_w8910_,
		_w9112_,
		_w9113_
	);
	LUT2 #(
		.INIT('h4)
	) name9080 (
		_w9111_,
		_w9113_,
		_w9114_
	);
	LUT3 #(
		.INIT('h82)
	) name9081 (
		_w37_,
		_w7069_,
		_w7071_,
		_w9115_
	);
	LUT3 #(
		.INIT('h82)
	) name9082 (
		_w3262_,
		_w6922_,
		_w6924_,
		_w9116_
	);
	LUT2 #(
		.INIT('h8)
	) name9083 (
		_w3214_,
		_w7062_,
		_w9117_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9084 (
		_w3249_,
		_w6669_,
		_w6919_,
		_w6921_,
		_w9118_
	);
	LUT2 #(
		.INIT('h1)
	) name9085 (
		_w9117_,
		_w9118_,
		_w9119_
	);
	LUT2 #(
		.INIT('h4)
	) name9086 (
		_w9116_,
		_w9119_,
		_w9120_
	);
	LUT2 #(
		.INIT('h8)
	) name9087 (
		\a[26] ,
		_w8904_,
		_w9121_
	);
	LUT3 #(
		.INIT('h4b)
	) name9088 (
		_w8901_,
		_w8903_,
		_w9121_,
		_w9122_
	);
	LUT4 #(
		.INIT('h6500)
	) name9089 (
		\a[23] ,
		_w9115_,
		_w9120_,
		_w9122_,
		_w9123_
	);
	LUT4 #(
		.INIT('h2882)
	) name9090 (
		_w37_,
		_w6914_,
		_w6916_,
		_w7067_,
		_w9124_
	);
	LUT4 #(
		.INIT('ha802)
	) name9091 (
		_w3249_,
		_w6689_,
		_w6911_,
		_w6913_,
		_w9125_
	);
	LUT4 #(
		.INIT('h007d)
	) name9092 (
		_w3262_,
		_w6914_,
		_w6916_,
		_w9125_,
		_w9126_
	);
	LUT4 #(
		.INIT('h5401)
	) name9093 (
		_w36_,
		_w6689_,
		_w6911_,
		_w6913_,
		_w9127_
	);
	LUT2 #(
		.INIT('h2)
	) name9094 (
		\a[23] ,
		_w9127_,
		_w9128_
	);
	LUT3 #(
		.INIT('h40)
	) name9095 (
		_w9124_,
		_w9126_,
		_w9128_,
		_w9129_
	);
	LUT3 #(
		.INIT('h28)
	) name9096 (
		_w37_,
		_w7062_,
		_w8358_,
		_w9130_
	);
	LUT4 #(
		.INIT('ha802)
	) name9097 (
		_w3214_,
		_w6689_,
		_w6911_,
		_w6913_,
		_w9131_
	);
	LUT4 #(
		.INIT('h007d)
	) name9098 (
		_w3249_,
		_w6914_,
		_w6916_,
		_w9131_,
		_w9132_
	);
	LUT3 #(
		.INIT('h70)
	) name9099 (
		_w3262_,
		_w7062_,
		_w9132_,
		_w9133_
	);
	LUT4 #(
		.INIT('h0800)
	) name9100 (
		_w8904_,
		_w9129_,
		_w9130_,
		_w9133_,
		_w9134_
	);
	LUT3 #(
		.INIT('h28)
	) name9101 (
		_w37_,
		_w7065_,
		_w7068_,
		_w9135_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9102 (
		_w3262_,
		_w6669_,
		_w6919_,
		_w6921_,
		_w9136_
	);
	LUT3 #(
		.INIT('h82)
	) name9103 (
		_w3214_,
		_w6914_,
		_w6916_,
		_w9137_
	);
	LUT3 #(
		.INIT('h07)
	) name9104 (
		_w3249_,
		_w7062_,
		_w9137_,
		_w9138_
	);
	LUT2 #(
		.INIT('h4)
	) name9105 (
		_w9136_,
		_w9138_,
		_w9139_
	);
	LUT4 #(
		.INIT('ha6aa)
	) name9106 (
		_w8904_,
		_w9129_,
		_w9130_,
		_w9133_,
		_w9140_
	);
	LUT4 #(
		.INIT('h6500)
	) name9107 (
		\a[23] ,
		_w9135_,
		_w9139_,
		_w9140_,
		_w9141_
	);
	LUT2 #(
		.INIT('h1)
	) name9108 (
		_w9134_,
		_w9141_,
		_w9142_
	);
	LUT4 #(
		.INIT('h009a)
	) name9109 (
		\a[23] ,
		_w9115_,
		_w9120_,
		_w9122_,
		_w9143_
	);
	LUT4 #(
		.INIT('h9a65)
	) name9110 (
		\a[23] ,
		_w9115_,
		_w9120_,
		_w9122_,
		_w9144_
	);
	LUT3 #(
		.INIT('h54)
	) name9111 (
		_w9123_,
		_w9142_,
		_w9143_,
		_w9145_
	);
	LUT2 #(
		.INIT('h2)
	) name9112 (
		_w9111_,
		_w9113_,
		_w9146_
	);
	LUT2 #(
		.INIT('h9)
	) name9113 (
		_w9111_,
		_w9113_,
		_w9147_
	);
	LUT4 #(
		.INIT('h9a65)
	) name9114 (
		\a[23] ,
		_w9101_,
		_w9105_,
		_w9106_,
		_w9148_
	);
	LUT4 #(
		.INIT('h4d00)
	) name9115 (
		_w9111_,
		_w9113_,
		_w9145_,
		_w9148_,
		_w9149_
	);
	LUT4 #(
		.INIT('h9a65)
	) name9116 (
		\a[23] ,
		_w9093_,
		_w9098_,
		_w9099_,
		_w9150_
	);
	LUT4 #(
		.INIT('h0155)
	) name9117 (
		_w9100_,
		_w9107_,
		_w9149_,
		_w9150_,
		_w9151_
	);
	LUT2 #(
		.INIT('h4)
	) name9118 (
		_w9087_,
		_w9091_,
		_w9152_
	);
	LUT2 #(
		.INIT('h9)
	) name9119 (
		_w9087_,
		_w9091_,
		_w9153_
	);
	LUT4 #(
		.INIT('h9699)
	) name9120 (
		\a[23] ,
		_w9080_,
		_w9081_,
		_w9085_,
		_w9154_
	);
	LUT4 #(
		.INIT('h2b00)
	) name9121 (
		_w9087_,
		_w9091_,
		_w9151_,
		_w9154_,
		_w9155_
	);
	LUT4 #(
		.INIT('h9a65)
	) name9122 (
		\a[23] ,
		_w9072_,
		_w9077_,
		_w9078_,
		_w9156_
	);
	LUT4 #(
		.INIT('h0155)
	) name9123 (
		_w9079_,
		_w9086_,
		_w9155_,
		_w9156_,
		_w9157_
	);
	LUT2 #(
		.INIT('h2)
	) name9124 (
		_w9069_,
		_w9070_,
		_w9158_
	);
	LUT2 #(
		.INIT('h9)
	) name9125 (
		_w9069_,
		_w9070_,
		_w9159_
	);
	LUT4 #(
		.INIT('h9a65)
	) name9126 (
		\a[23] ,
		_w9059_,
		_w9063_,
		_w9064_,
		_w9160_
	);
	LUT4 #(
		.INIT('h4d00)
	) name9127 (
		_w9069_,
		_w9070_,
		_w9157_,
		_w9160_,
		_w9161_
	);
	LUT4 #(
		.INIT('h9a65)
	) name9128 (
		\a[23] ,
		_w9051_,
		_w9056_,
		_w9057_,
		_w9162_
	);
	LUT4 #(
		.INIT('h0155)
	) name9129 (
		_w9058_,
		_w9065_,
		_w9161_,
		_w9162_,
		_w9163_
	);
	LUT2 #(
		.INIT('h2)
	) name9130 (
		_w9048_,
		_w9049_,
		_w9164_
	);
	LUT2 #(
		.INIT('h9)
	) name9131 (
		_w9048_,
		_w9049_,
		_w9165_
	);
	LUT4 #(
		.INIT('h9a65)
	) name9132 (
		\a[23] ,
		_w9038_,
		_w9042_,
		_w9043_,
		_w9166_
	);
	LUT4 #(
		.INIT('h4d00)
	) name9133 (
		_w9048_,
		_w9049_,
		_w9163_,
		_w9166_,
		_w9167_
	);
	LUT4 #(
		.INIT('h9a65)
	) name9134 (
		\a[23] ,
		_w9030_,
		_w9035_,
		_w9036_,
		_w9168_
	);
	LUT4 #(
		.INIT('h0155)
	) name9135 (
		_w9037_,
		_w9044_,
		_w9167_,
		_w9168_,
		_w9169_
	);
	LUT2 #(
		.INIT('h2)
	) name9136 (
		_w9027_,
		_w9028_,
		_w9170_
	);
	LUT2 #(
		.INIT('h9)
	) name9137 (
		_w9027_,
		_w9028_,
		_w9171_
	);
	LUT4 #(
		.INIT('h9a65)
	) name9138 (
		\a[23] ,
		_w9017_,
		_w9021_,
		_w9022_,
		_w9172_
	);
	LUT4 #(
		.INIT('h4d00)
	) name9139 (
		_w9027_,
		_w9028_,
		_w9169_,
		_w9172_,
		_w9173_
	);
	LUT4 #(
		.INIT('h9a65)
	) name9140 (
		\a[23] ,
		_w9009_,
		_w9014_,
		_w9015_,
		_w9174_
	);
	LUT4 #(
		.INIT('h0155)
	) name9141 (
		_w9016_,
		_w9023_,
		_w9173_,
		_w9174_,
		_w9175_
	);
	LUT4 #(
		.INIT('h0096)
	) name9142 (
		_w8946_,
		_w8947_,
		_w8951_,
		_w9175_,
		_w9176_
	);
	LUT4 #(
		.INIT('h6900)
	) name9143 (
		_w8946_,
		_w8947_,
		_w8951_,
		_w9175_,
		_w9177_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9144 (
		_w3311_,
		_w3882_,
		_w6954_,
		_w6956_,
		_w9178_
	);
	LUT4 #(
		.INIT('h007d)
	) name9145 (
		_w3645_,
		_w3706_,
		_w6957_,
		_w9178_,
		_w9179_
	);
	LUT3 #(
		.INIT('h70)
	) name9146 (
		_w3654_,
		_w7020_,
		_w9179_,
		_w9180_
	);
	LUT4 #(
		.INIT('h95aa)
	) name9147 (
		\a[20] ,
		_w3312_,
		_w7465_,
		_w9180_,
		_w9181_
	);
	LUT3 #(
		.INIT('h54)
	) name9148 (
		_w9176_,
		_w9177_,
		_w9181_,
		_w9182_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9149 (
		_w3710_,
		_w7016_,
		_w7115_,
		_w7116_,
		_w9183_
	);
	LUT4 #(
		.INIT('h04c8)
	) name9150 (
		_w3257_,
		_w3886_,
		_w6964_,
		_w6966_,
		_w9184_
	);
	LUT3 #(
		.INIT('h82)
	) name9151 (
		_w3709_,
		_w6960_,
		_w6962_,
		_w9185_
	);
	LUT3 #(
		.INIT('h07)
	) name9152 (
		_w3877_,
		_w7014_,
		_w9185_,
		_w9186_
	);
	LUT2 #(
		.INIT('h4)
	) name9153 (
		_w9184_,
		_w9186_,
		_w9187_
	);
	LUT3 #(
		.INIT('h9a)
	) name9154 (
		\a[17] ,
		_w9183_,
		_w9187_,
		_w9188_
	);
	LUT4 #(
		.INIT('hf660)
	) name9155 (
		_w8960_,
		_w9008_,
		_w9182_,
		_w9188_,
		_w9189_
	);
	LUT4 #(
		.INIT('h0096)
	) name9156 (
		_w8806_,
		_w8961_,
		_w8968_,
		_w9189_,
		_w9190_
	);
	LUT4 #(
		.INIT('h6900)
	) name9157 (
		_w8806_,
		_w8961_,
		_w8968_,
		_w9189_,
		_w9191_
	);
	LUT3 #(
		.INIT('h82)
	) name9158 (
		_w4034_,
		_w7123_,
		_w7125_,
		_w9192_
	);
	LUT3 #(
		.INIT('h84)
	) name9159 (
		_w2872_,
		_w4382_,
		_w6975_,
		_w9193_
	);
	LUT2 #(
		.INIT('h8)
	) name9160 (
		_w4033_,
		_w7008_,
		_w9194_
	);
	LUT4 #(
		.INIT('h04c8)
	) name9161 (
		_w2983_,
		_w4367_,
		_w6972_,
		_w6974_,
		_w9195_
	);
	LUT2 #(
		.INIT('h1)
	) name9162 (
		_w9194_,
		_w9195_,
		_w9196_
	);
	LUT2 #(
		.INIT('h4)
	) name9163 (
		_w9193_,
		_w9196_,
		_w9197_
	);
	LUT3 #(
		.INIT('h9a)
	) name9164 (
		\a[14] ,
		_w9192_,
		_w9197_,
		_w9198_
	);
	LUT3 #(
		.INIT('h54)
	) name9165 (
		_w9190_,
		_w9191_,
		_w9198_,
		_w9199_
	);
	LUT3 #(
		.INIT('h54)
	) name9166 (
		_w9005_,
		_w9006_,
		_w9199_,
		_w9200_
	);
	LUT4 #(
		.INIT('h9669)
	) name9167 (
		_w8774_,
		_w8970_,
		_w8971_,
		_w8977_,
		_w9201_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9168 (
		_w4459_,
		_w6998_,
		_w7133_,
		_w7134_,
		_w9202_
	);
	LUT4 #(
		.INIT('h04c8)
	) name9169 (
		_w2411_,
		_w4700_,
		_w6983_,
		_w6993_,
		_w9203_
	);
	LUT3 #(
		.INIT('h84)
	) name9170 (
		_w2546_,
		_w4458_,
		_w6981_,
		_w9204_
	);
	LUT3 #(
		.INIT('h07)
	) name9171 (
		_w4684_,
		_w6996_,
		_w9204_,
		_w9205_
	);
	LUT2 #(
		.INIT('h4)
	) name9172 (
		_w9203_,
		_w9205_,
		_w9206_
	);
	LUT3 #(
		.INIT('h9a)
	) name9173 (
		\a[11] ,
		_w9202_,
		_w9206_,
		_w9207_
	);
	LUT4 #(
		.INIT('h1051)
	) name9174 (
		_w9000_,
		_w9200_,
		_w9201_,
		_w9207_,
		_w9208_
	);
	LUT4 #(
		.INIT('h8a08)
	) name9175 (
		_w9000_,
		_w9200_,
		_w9201_,
		_w9207_,
		_w9209_
	);
	LUT4 #(
		.INIT('h9669)
	) name9176 (
		_w8626_,
		_w8775_,
		_w8782_,
		_w8978_,
		_w9210_
	);
	LUT4 #(
		.INIT('h3132)
	) name9177 (
		_w8987_,
		_w9208_,
		_w9209_,
		_w9210_,
		_w9211_
	);
	LUT3 #(
		.INIT('h06)
	) name9178 (
		_w8989_,
		_w8991_,
		_w9211_,
		_w9212_
	);
	LUT4 #(
		.INIT('h65a6)
	) name9179 (
		_w9000_,
		_w9200_,
		_w9201_,
		_w9207_,
		_w9213_
	);
	LUT3 #(
		.INIT('h69)
	) name9180 (
		_w8987_,
		_w9210_,
		_w9213_,
		_w9214_
	);
	LUT4 #(
		.INIT('h04c8)
	) name9181 (
		_w2622_,
		_w4458_,
		_w6978_,
		_w6980_,
		_w9215_
	);
	LUT4 #(
		.INIT('h007b)
	) name9182 (
		_w2546_,
		_w4684_,
		_w6981_,
		_w9215_,
		_w9216_
	);
	LUT3 #(
		.INIT('h70)
	) name9183 (
		_w4700_,
		_w6996_,
		_w9216_,
		_w9217_
	);
	LUT4 #(
		.INIT('h95aa)
	) name9184 (
		\a[11] ,
		_w4459_,
		_w7500_,
		_w9217_,
		_w9218_
	);
	LUT4 #(
		.INIT('h9669)
	) name9185 (
		_w8806_,
		_w8961_,
		_w8968_,
		_w9189_,
		_w9219_
	);
	LUT4 #(
		.INIT('h9669)
	) name9186 (
		_w8960_,
		_w9008_,
		_w9182_,
		_w9188_,
		_w9220_
	);
	LUT3 #(
		.INIT('h1e)
	) name9187 (
		_w9023_,
		_w9173_,
		_w9174_,
		_w9221_
	);
	LUT3 #(
		.INIT('h82)
	) name9188 (
		_w3312_,
		_w7105_,
		_w7107_,
		_w9222_
	);
	LUT3 #(
		.INIT('h82)
	) name9189 (
		_w3654_,
		_w3706_,
		_w6957_,
		_w9223_
	);
	LUT2 #(
		.INIT('h8)
	) name9190 (
		_w3311_,
		_w7026_,
		_w9224_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9191 (
		_w3645_,
		_w3882_,
		_w6954_,
		_w6956_,
		_w9225_
	);
	LUT2 #(
		.INIT('h1)
	) name9192 (
		_w9224_,
		_w9225_,
		_w9226_
	);
	LUT2 #(
		.INIT('h4)
	) name9193 (
		_w9223_,
		_w9226_,
		_w9227_
	);
	LUT4 #(
		.INIT('h4844)
	) name9194 (
		\a[20] ,
		_w9221_,
		_w9222_,
		_w9227_,
		_w9228_
	);
	LUT4 #(
		.INIT('h54ab)
	) name9195 (
		_w9029_,
		_w9169_,
		_w9170_,
		_w9172_,
		_w9229_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9196 (
		_w3312_,
		_w7028_,
		_w7103_,
		_w7104_,
		_w9230_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9197 (
		_w3654_,
		_w3882_,
		_w6954_,
		_w6956_,
		_w9231_
	);
	LUT3 #(
		.INIT('h82)
	) name9198 (
		_w3311_,
		_w4030_,
		_w6952_,
		_w9232_
	);
	LUT3 #(
		.INIT('h07)
	) name9199 (
		_w3645_,
		_w7026_,
		_w9232_,
		_w9233_
	);
	LUT2 #(
		.INIT('h4)
	) name9200 (
		_w9231_,
		_w9233_,
		_w9234_
	);
	LUT4 #(
		.INIT('h4844)
	) name9201 (
		\a[20] ,
		_w9229_,
		_w9230_,
		_w9234_,
		_w9235_
	);
	LUT2 #(
		.INIT('h9)
	) name9202 (
		_w9169_,
		_w9171_,
		_w9236_
	);
	LUT4 #(
		.INIT('h2228)
	) name9203 (
		_w3311_,
		_w4099_,
		_w4378_,
		_w6951_,
		_w9237_
	);
	LUT4 #(
		.INIT('h007d)
	) name9204 (
		_w3645_,
		_w4030_,
		_w6952_,
		_w9237_,
		_w9238_
	);
	LUT3 #(
		.INIT('h70)
	) name9205 (
		_w3654_,
		_w7026_,
		_w9238_,
		_w9239_
	);
	LUT4 #(
		.INIT('h95aa)
	) name9206 (
		\a[20] ,
		_w3312_,
		_w7562_,
		_w9239_,
		_w9240_
	);
	LUT2 #(
		.INIT('h2)
	) name9207 (
		_w9236_,
		_w9240_,
		_w9241_
	);
	LUT3 #(
		.INIT('h1e)
	) name9208 (
		_w9044_,
		_w9167_,
		_w9168_,
		_w9242_
	);
	LUT3 #(
		.INIT('h82)
	) name9209 (
		_w3312_,
		_w7099_,
		_w7101_,
		_w9243_
	);
	LUT3 #(
		.INIT('h82)
	) name9210 (
		_w3654_,
		_w4030_,
		_w6952_,
		_w9244_
	);
	LUT2 #(
		.INIT('h8)
	) name9211 (
		_w3311_,
		_w7032_,
		_w9245_
	);
	LUT4 #(
		.INIT('h2228)
	) name9212 (
		_w3645_,
		_w4099_,
		_w4378_,
		_w6951_,
		_w9246_
	);
	LUT2 #(
		.INIT('h1)
	) name9213 (
		_w9245_,
		_w9246_,
		_w9247_
	);
	LUT2 #(
		.INIT('h4)
	) name9214 (
		_w9244_,
		_w9247_,
		_w9248_
	);
	LUT4 #(
		.INIT('h4844)
	) name9215 (
		\a[20] ,
		_w9242_,
		_w9243_,
		_w9248_,
		_w9249_
	);
	LUT4 #(
		.INIT('h54ab)
	) name9216 (
		_w9050_,
		_w9163_,
		_w9164_,
		_w9166_,
		_w9250_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9217 (
		_w3312_,
		_w7034_,
		_w7097_,
		_w7098_,
		_w9251_
	);
	LUT4 #(
		.INIT('h2228)
	) name9218 (
		_w3654_,
		_w4099_,
		_w4378_,
		_w6951_,
		_w9252_
	);
	LUT3 #(
		.INIT('h82)
	) name9219 (
		_w3311_,
		_w6947_,
		_w6949_,
		_w9253_
	);
	LUT3 #(
		.INIT('h07)
	) name9220 (
		_w3645_,
		_w7032_,
		_w9253_,
		_w9254_
	);
	LUT2 #(
		.INIT('h4)
	) name9221 (
		_w9252_,
		_w9254_,
		_w9255_
	);
	LUT4 #(
		.INIT('h4844)
	) name9222 (
		\a[20] ,
		_w9250_,
		_w9251_,
		_w9255_,
		_w9256_
	);
	LUT2 #(
		.INIT('h9)
	) name9223 (
		_w9163_,
		_w9165_,
		_w9257_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9224 (
		_w3311_,
		_w4695_,
		_w6944_,
		_w6946_,
		_w9258_
	);
	LUT4 #(
		.INIT('h007d)
	) name9225 (
		_w3645_,
		_w6947_,
		_w6949_,
		_w9258_,
		_w9259_
	);
	LUT3 #(
		.INIT('h70)
	) name9226 (
		_w3654_,
		_w7032_,
		_w9259_,
		_w9260_
	);
	LUT4 #(
		.INIT('h95aa)
	) name9227 (
		\a[20] ,
		_w3312_,
		_w7882_,
		_w9260_,
		_w9261_
	);
	LUT2 #(
		.INIT('h2)
	) name9228 (
		_w9257_,
		_w9261_,
		_w9262_
	);
	LUT3 #(
		.INIT('h1e)
	) name9229 (
		_w9065_,
		_w9161_,
		_w9162_,
		_w9263_
	);
	LUT3 #(
		.INIT('h82)
	) name9230 (
		_w3312_,
		_w7093_,
		_w7095_,
		_w9264_
	);
	LUT3 #(
		.INIT('h82)
	) name9231 (
		_w3654_,
		_w6947_,
		_w6949_,
		_w9265_
	);
	LUT2 #(
		.INIT('h8)
	) name9232 (
		_w3311_,
		_w7038_,
		_w9266_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9233 (
		_w3645_,
		_w4695_,
		_w6944_,
		_w6946_,
		_w9267_
	);
	LUT2 #(
		.INIT('h1)
	) name9234 (
		_w9266_,
		_w9267_,
		_w9268_
	);
	LUT2 #(
		.INIT('h4)
	) name9235 (
		_w9265_,
		_w9268_,
		_w9269_
	);
	LUT4 #(
		.INIT('h4844)
	) name9236 (
		\a[20] ,
		_w9263_,
		_w9264_,
		_w9269_,
		_w9270_
	);
	LUT4 #(
		.INIT('h54ab)
	) name9237 (
		_w9071_,
		_w9157_,
		_w9158_,
		_w9160_,
		_w9271_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9238 (
		_w3312_,
		_w7040_,
		_w7091_,
		_w7092_,
		_w9272_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9239 (
		_w3654_,
		_w4695_,
		_w6944_,
		_w6946_,
		_w9273_
	);
	LUT3 #(
		.INIT('h82)
	) name9240 (
		_w3311_,
		_w6940_,
		_w6942_,
		_w9274_
	);
	LUT3 #(
		.INIT('h07)
	) name9241 (
		_w3645_,
		_w7038_,
		_w9274_,
		_w9275_
	);
	LUT2 #(
		.INIT('h4)
	) name9242 (
		_w9273_,
		_w9275_,
		_w9276_
	);
	LUT4 #(
		.INIT('h4844)
	) name9243 (
		\a[20] ,
		_w9271_,
		_w9272_,
		_w9276_,
		_w9277_
	);
	LUT2 #(
		.INIT('h9)
	) name9244 (
		_w9157_,
		_w9159_,
		_w9278_
	);
	LUT4 #(
		.INIT('h2228)
	) name9245 (
		_w3311_,
		_w5067_,
		_w5282_,
		_w6939_,
		_w9279_
	);
	LUT4 #(
		.INIT('h007d)
	) name9246 (
		_w3645_,
		_w6940_,
		_w6942_,
		_w9279_,
		_w9280_
	);
	LUT3 #(
		.INIT('h70)
	) name9247 (
		_w3654_,
		_w7038_,
		_w9280_,
		_w9281_
	);
	LUT4 #(
		.INIT('h95aa)
	) name9248 (
		\a[20] ,
		_w3312_,
		_w8018_,
		_w9281_,
		_w9282_
	);
	LUT2 #(
		.INIT('h2)
	) name9249 (
		_w9278_,
		_w9282_,
		_w9283_
	);
	LUT3 #(
		.INIT('h1e)
	) name9250 (
		_w9086_,
		_w9155_,
		_w9156_,
		_w9284_
	);
	LUT3 #(
		.INIT('h82)
	) name9251 (
		_w3312_,
		_w7087_,
		_w7089_,
		_w9285_
	);
	LUT3 #(
		.INIT('h82)
	) name9252 (
		_w3654_,
		_w6940_,
		_w6942_,
		_w9286_
	);
	LUT2 #(
		.INIT('h8)
	) name9253 (
		_w3311_,
		_w7044_,
		_w9287_
	);
	LUT4 #(
		.INIT('h2228)
	) name9254 (
		_w3645_,
		_w5067_,
		_w5282_,
		_w6939_,
		_w9288_
	);
	LUT2 #(
		.INIT('h1)
	) name9255 (
		_w9287_,
		_w9288_,
		_w9289_
	);
	LUT2 #(
		.INIT('h4)
	) name9256 (
		_w9286_,
		_w9289_,
		_w9290_
	);
	LUT4 #(
		.INIT('h4844)
	) name9257 (
		\a[20] ,
		_w9284_,
		_w9285_,
		_w9290_,
		_w9291_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9258 (
		_w3312_,
		_w7046_,
		_w7085_,
		_w7086_,
		_w9292_
	);
	LUT4 #(
		.INIT('h2228)
	) name9259 (
		_w3654_,
		_w5067_,
		_w5282_,
		_w6939_,
		_w9293_
	);
	LUT3 #(
		.INIT('h82)
	) name9260 (
		_w3311_,
		_w6935_,
		_w6937_,
		_w9294_
	);
	LUT3 #(
		.INIT('h07)
	) name9261 (
		_w3645_,
		_w7044_,
		_w9294_,
		_w9295_
	);
	LUT2 #(
		.INIT('h4)
	) name9262 (
		_w9293_,
		_w9295_,
		_w9296_
	);
	LUT4 #(
		.INIT('h54ab)
	) name9263 (
		_w9092_,
		_w9151_,
		_w9152_,
		_w9154_,
		_w9297_
	);
	LUT4 #(
		.INIT('h6500)
	) name9264 (
		\a[20] ,
		_w9292_,
		_w9296_,
		_w9297_,
		_w9298_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9265 (
		_w3311_,
		_w6043_,
		_w6933_,
		_w6934_,
		_w9299_
	);
	LUT4 #(
		.INIT('h007d)
	) name9266 (
		_w3645_,
		_w6935_,
		_w6937_,
		_w9299_,
		_w9300_
	);
	LUT3 #(
		.INIT('h70)
	) name9267 (
		_w3654_,
		_w7044_,
		_w9300_,
		_w9301_
	);
	LUT4 #(
		.INIT('h95aa)
	) name9268 (
		\a[20] ,
		_w3312_,
		_w8005_,
		_w9301_,
		_w9302_
	);
	LUT2 #(
		.INIT('h9)
	) name9269 (
		_w9151_,
		_w9153_,
		_w9303_
	);
	LUT2 #(
		.INIT('h4)
	) name9270 (
		_w9302_,
		_w9303_,
		_w9304_
	);
	LUT3 #(
		.INIT('h1e)
	) name9271 (
		_w9107_,
		_w9149_,
		_w9150_,
		_w9305_
	);
	LUT3 #(
		.INIT('h82)
	) name9272 (
		_w3312_,
		_w7081_,
		_w7083_,
		_w9306_
	);
	LUT3 #(
		.INIT('h82)
	) name9273 (
		_w3654_,
		_w6935_,
		_w6937_,
		_w9307_
	);
	LUT2 #(
		.INIT('h8)
	) name9274 (
		_w3311_,
		_w7050_,
		_w9308_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9275 (
		_w3645_,
		_w6043_,
		_w6933_,
		_w6934_,
		_w9309_
	);
	LUT2 #(
		.INIT('h1)
	) name9276 (
		_w9308_,
		_w9309_,
		_w9310_
	);
	LUT2 #(
		.INIT('h4)
	) name9277 (
		_w9307_,
		_w9310_,
		_w9311_
	);
	LUT4 #(
		.INIT('h4844)
	) name9278 (
		\a[20] ,
		_w9305_,
		_w9306_,
		_w9311_,
		_w9312_
	);
	LUT4 #(
		.INIT('h54ab)
	) name9279 (
		_w9114_,
		_w9145_,
		_w9146_,
		_w9148_,
		_w9313_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9280 (
		_w3312_,
		_w7052_,
		_w7079_,
		_w7080_,
		_w9314_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9281 (
		_w3654_,
		_w6043_,
		_w6933_,
		_w6934_,
		_w9315_
	);
	LUT3 #(
		.INIT('h82)
	) name9282 (
		_w3311_,
		_w6929_,
		_w6931_,
		_w9316_
	);
	LUT3 #(
		.INIT('h07)
	) name9283 (
		_w3645_,
		_w7050_,
		_w9316_,
		_w9317_
	);
	LUT2 #(
		.INIT('h4)
	) name9284 (
		_w9315_,
		_w9317_,
		_w9318_
	);
	LUT4 #(
		.INIT('h4844)
	) name9285 (
		\a[20] ,
		_w9313_,
		_w9314_,
		_w9318_,
		_w9319_
	);
	LUT2 #(
		.INIT('h9)
	) name9286 (
		_w9145_,
		_w9147_,
		_w9320_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9287 (
		_w3311_,
		_w6645_,
		_w6926_,
		_w6928_,
		_w9321_
	);
	LUT4 #(
		.INIT('h007d)
	) name9288 (
		_w3645_,
		_w6929_,
		_w6931_,
		_w9321_,
		_w9322_
	);
	LUT3 #(
		.INIT('h70)
	) name9289 (
		_w3654_,
		_w7050_,
		_w9322_,
		_w9323_
	);
	LUT4 #(
		.INIT('h95aa)
	) name9290 (
		\a[20] ,
		_w3312_,
		_w8227_,
		_w9323_,
		_w9324_
	);
	LUT2 #(
		.INIT('h2)
	) name9291 (
		_w9320_,
		_w9324_,
		_w9325_
	);
	LUT3 #(
		.INIT('h82)
	) name9292 (
		_w3312_,
		_w7075_,
		_w7077_,
		_w9326_
	);
	LUT3 #(
		.INIT('h82)
	) name9293 (
		_w3654_,
		_w6929_,
		_w6931_,
		_w9327_
	);
	LUT2 #(
		.INIT('h8)
	) name9294 (
		_w3311_,
		_w7056_,
		_w9328_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9295 (
		_w3645_,
		_w6645_,
		_w6926_,
		_w6928_,
		_w9329_
	);
	LUT2 #(
		.INIT('h1)
	) name9296 (
		_w9328_,
		_w9329_,
		_w9330_
	);
	LUT2 #(
		.INIT('h4)
	) name9297 (
		_w9327_,
		_w9330_,
		_w9331_
	);
	LUT2 #(
		.INIT('h9)
	) name9298 (
		_w9142_,
		_w9144_,
		_w9332_
	);
	LUT4 #(
		.INIT('h6500)
	) name9299 (
		\a[20] ,
		_w9326_,
		_w9331_,
		_w9332_,
		_w9333_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9300 (
		_w3312_,
		_w7058_,
		_w7073_,
		_w7074_,
		_w9334_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9301 (
		_w3654_,
		_w6645_,
		_w6926_,
		_w6928_,
		_w9335_
	);
	LUT3 #(
		.INIT('h82)
	) name9302 (
		_w3311_,
		_w6922_,
		_w6924_,
		_w9336_
	);
	LUT3 #(
		.INIT('h07)
	) name9303 (
		_w3645_,
		_w7056_,
		_w9336_,
		_w9337_
	);
	LUT2 #(
		.INIT('h4)
	) name9304 (
		_w9335_,
		_w9337_,
		_w9338_
	);
	LUT4 #(
		.INIT('h9a65)
	) name9305 (
		\a[23] ,
		_w9135_,
		_w9139_,
		_w9140_,
		_w9339_
	);
	LUT4 #(
		.INIT('h6500)
	) name9306 (
		\a[20] ,
		_w9334_,
		_w9338_,
		_w9339_,
		_w9340_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9307 (
		_w3311_,
		_w6669_,
		_w6919_,
		_w6921_,
		_w9341_
	);
	LUT4 #(
		.INIT('h007d)
	) name9308 (
		_w3645_,
		_w6922_,
		_w6924_,
		_w9341_,
		_w9342_
	);
	LUT3 #(
		.INIT('h70)
	) name9309 (
		_w3654_,
		_w7056_,
		_w9342_,
		_w9343_
	);
	LUT4 #(
		.INIT('h95aa)
	) name9310 (
		\a[20] ,
		_w3312_,
		_w8298_,
		_w9343_,
		_w9344_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name9311 (
		\a[23] ,
		_w9127_,
		_w9124_,
		_w9126_,
		_w9345_
	);
	LUT3 #(
		.INIT('h4b)
	) name9312 (
		_w9130_,
		_w9133_,
		_w9345_,
		_w9346_
	);
	LUT2 #(
		.INIT('h4)
	) name9313 (
		_w9344_,
		_w9346_,
		_w9347_
	);
	LUT3 #(
		.INIT('h82)
	) name9314 (
		_w3312_,
		_w7069_,
		_w7071_,
		_w9348_
	);
	LUT3 #(
		.INIT('h82)
	) name9315 (
		_w3654_,
		_w6922_,
		_w6924_,
		_w9349_
	);
	LUT2 #(
		.INIT('h8)
	) name9316 (
		_w3311_,
		_w7062_,
		_w9350_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9317 (
		_w3645_,
		_w6669_,
		_w6919_,
		_w6921_,
		_w9351_
	);
	LUT2 #(
		.INIT('h1)
	) name9318 (
		_w9350_,
		_w9351_,
		_w9352_
	);
	LUT2 #(
		.INIT('h4)
	) name9319 (
		_w9349_,
		_w9352_,
		_w9353_
	);
	LUT2 #(
		.INIT('h8)
	) name9320 (
		\a[23] ,
		_w9127_,
		_w9354_
	);
	LUT3 #(
		.INIT('h4b)
	) name9321 (
		_w9124_,
		_w9126_,
		_w9354_,
		_w9355_
	);
	LUT4 #(
		.INIT('h6500)
	) name9322 (
		\a[20] ,
		_w9348_,
		_w9353_,
		_w9355_,
		_w9356_
	);
	LUT4 #(
		.INIT('h2882)
	) name9323 (
		_w3312_,
		_w6914_,
		_w6916_,
		_w7067_,
		_w9357_
	);
	LUT4 #(
		.INIT('ha802)
	) name9324 (
		_w3645_,
		_w6689_,
		_w6911_,
		_w6913_,
		_w9358_
	);
	LUT4 #(
		.INIT('h007d)
	) name9325 (
		_w3654_,
		_w6914_,
		_w6916_,
		_w9358_,
		_w9359_
	);
	LUT4 #(
		.INIT('h5401)
	) name9326 (
		_w3310_,
		_w6689_,
		_w6911_,
		_w6913_,
		_w9360_
	);
	LUT2 #(
		.INIT('h2)
	) name9327 (
		\a[20] ,
		_w9360_,
		_w9361_
	);
	LUT3 #(
		.INIT('h40)
	) name9328 (
		_w9357_,
		_w9359_,
		_w9361_,
		_w9362_
	);
	LUT3 #(
		.INIT('h28)
	) name9329 (
		_w3312_,
		_w7062_,
		_w8358_,
		_w9363_
	);
	LUT4 #(
		.INIT('ha802)
	) name9330 (
		_w3311_,
		_w6689_,
		_w6911_,
		_w6913_,
		_w9364_
	);
	LUT4 #(
		.INIT('h007d)
	) name9331 (
		_w3645_,
		_w6914_,
		_w6916_,
		_w9364_,
		_w9365_
	);
	LUT3 #(
		.INIT('h70)
	) name9332 (
		_w3654_,
		_w7062_,
		_w9365_,
		_w9366_
	);
	LUT4 #(
		.INIT('h0800)
	) name9333 (
		_w9127_,
		_w9362_,
		_w9363_,
		_w9366_,
		_w9367_
	);
	LUT3 #(
		.INIT('h28)
	) name9334 (
		_w3312_,
		_w7065_,
		_w7068_,
		_w9368_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9335 (
		_w3654_,
		_w6669_,
		_w6919_,
		_w6921_,
		_w9369_
	);
	LUT3 #(
		.INIT('h82)
	) name9336 (
		_w3311_,
		_w6914_,
		_w6916_,
		_w9370_
	);
	LUT3 #(
		.INIT('h07)
	) name9337 (
		_w3645_,
		_w7062_,
		_w9370_,
		_w9371_
	);
	LUT2 #(
		.INIT('h4)
	) name9338 (
		_w9369_,
		_w9371_,
		_w9372_
	);
	LUT4 #(
		.INIT('ha6aa)
	) name9339 (
		_w9127_,
		_w9362_,
		_w9363_,
		_w9366_,
		_w9373_
	);
	LUT4 #(
		.INIT('h6500)
	) name9340 (
		\a[20] ,
		_w9368_,
		_w9372_,
		_w9373_,
		_w9374_
	);
	LUT2 #(
		.INIT('h1)
	) name9341 (
		_w9367_,
		_w9374_,
		_w9375_
	);
	LUT4 #(
		.INIT('h009a)
	) name9342 (
		\a[20] ,
		_w9348_,
		_w9353_,
		_w9355_,
		_w9376_
	);
	LUT4 #(
		.INIT('h9a65)
	) name9343 (
		\a[20] ,
		_w9348_,
		_w9353_,
		_w9355_,
		_w9377_
	);
	LUT3 #(
		.INIT('h54)
	) name9344 (
		_w9356_,
		_w9375_,
		_w9376_,
		_w9378_
	);
	LUT2 #(
		.INIT('h2)
	) name9345 (
		_w9344_,
		_w9346_,
		_w9379_
	);
	LUT2 #(
		.INIT('h9)
	) name9346 (
		_w9344_,
		_w9346_,
		_w9380_
	);
	LUT4 #(
		.INIT('h9a65)
	) name9347 (
		\a[20] ,
		_w9334_,
		_w9338_,
		_w9339_,
		_w9381_
	);
	LUT4 #(
		.INIT('h4d00)
	) name9348 (
		_w9344_,
		_w9346_,
		_w9378_,
		_w9381_,
		_w9382_
	);
	LUT4 #(
		.INIT('h9a65)
	) name9349 (
		\a[20] ,
		_w9326_,
		_w9331_,
		_w9332_,
		_w9383_
	);
	LUT4 #(
		.INIT('h0155)
	) name9350 (
		_w9333_,
		_w9340_,
		_w9382_,
		_w9383_,
		_w9384_
	);
	LUT2 #(
		.INIT('h4)
	) name9351 (
		_w9320_,
		_w9324_,
		_w9385_
	);
	LUT2 #(
		.INIT('h9)
	) name9352 (
		_w9320_,
		_w9324_,
		_w9386_
	);
	LUT4 #(
		.INIT('h9699)
	) name9353 (
		\a[20] ,
		_w9313_,
		_w9314_,
		_w9318_,
		_w9387_
	);
	LUT4 #(
		.INIT('h2b00)
	) name9354 (
		_w9320_,
		_w9324_,
		_w9384_,
		_w9387_,
		_w9388_
	);
	LUT4 #(
		.INIT('h9699)
	) name9355 (
		\a[20] ,
		_w9305_,
		_w9306_,
		_w9311_,
		_w9389_
	);
	LUT4 #(
		.INIT('h0155)
	) name9356 (
		_w9312_,
		_w9319_,
		_w9388_,
		_w9389_,
		_w9390_
	);
	LUT2 #(
		.INIT('h2)
	) name9357 (
		_w9302_,
		_w9303_,
		_w9391_
	);
	LUT2 #(
		.INIT('h9)
	) name9358 (
		_w9302_,
		_w9303_,
		_w9392_
	);
	LUT4 #(
		.INIT('h9a65)
	) name9359 (
		\a[20] ,
		_w9292_,
		_w9296_,
		_w9297_,
		_w9393_
	);
	LUT4 #(
		.INIT('h4d00)
	) name9360 (
		_w9302_,
		_w9303_,
		_w9390_,
		_w9393_,
		_w9394_
	);
	LUT4 #(
		.INIT('h9699)
	) name9361 (
		\a[20] ,
		_w9284_,
		_w9285_,
		_w9290_,
		_w9395_
	);
	LUT4 #(
		.INIT('h0155)
	) name9362 (
		_w9291_,
		_w9298_,
		_w9394_,
		_w9395_,
		_w9396_
	);
	LUT2 #(
		.INIT('h4)
	) name9363 (
		_w9278_,
		_w9282_,
		_w9397_
	);
	LUT2 #(
		.INIT('h9)
	) name9364 (
		_w9278_,
		_w9282_,
		_w9398_
	);
	LUT4 #(
		.INIT('h9699)
	) name9365 (
		\a[20] ,
		_w9271_,
		_w9272_,
		_w9276_,
		_w9399_
	);
	LUT4 #(
		.INIT('h2b00)
	) name9366 (
		_w9278_,
		_w9282_,
		_w9396_,
		_w9399_,
		_w9400_
	);
	LUT4 #(
		.INIT('h9699)
	) name9367 (
		\a[20] ,
		_w9263_,
		_w9264_,
		_w9269_,
		_w9401_
	);
	LUT4 #(
		.INIT('h0155)
	) name9368 (
		_w9270_,
		_w9277_,
		_w9400_,
		_w9401_,
		_w9402_
	);
	LUT2 #(
		.INIT('h4)
	) name9369 (
		_w9257_,
		_w9261_,
		_w9403_
	);
	LUT2 #(
		.INIT('h9)
	) name9370 (
		_w9257_,
		_w9261_,
		_w9404_
	);
	LUT4 #(
		.INIT('h9699)
	) name9371 (
		\a[20] ,
		_w9250_,
		_w9251_,
		_w9255_,
		_w9405_
	);
	LUT4 #(
		.INIT('h2b00)
	) name9372 (
		_w9257_,
		_w9261_,
		_w9402_,
		_w9405_,
		_w9406_
	);
	LUT4 #(
		.INIT('h9699)
	) name9373 (
		\a[20] ,
		_w9242_,
		_w9243_,
		_w9248_,
		_w9407_
	);
	LUT4 #(
		.INIT('h0155)
	) name9374 (
		_w9249_,
		_w9256_,
		_w9406_,
		_w9407_,
		_w9408_
	);
	LUT2 #(
		.INIT('h4)
	) name9375 (
		_w9236_,
		_w9240_,
		_w9409_
	);
	LUT2 #(
		.INIT('h9)
	) name9376 (
		_w9236_,
		_w9240_,
		_w9410_
	);
	LUT4 #(
		.INIT('h9699)
	) name9377 (
		\a[20] ,
		_w9229_,
		_w9230_,
		_w9234_,
		_w9411_
	);
	LUT4 #(
		.INIT('h2b00)
	) name9378 (
		_w9236_,
		_w9240_,
		_w9408_,
		_w9411_,
		_w9412_
	);
	LUT4 #(
		.INIT('h9699)
	) name9379 (
		\a[20] ,
		_w9221_,
		_w9222_,
		_w9227_,
		_w9413_
	);
	LUT4 #(
		.INIT('h0155)
	) name9380 (
		_w9228_,
		_w9235_,
		_w9412_,
		_w9413_,
		_w9414_
	);
	LUT4 #(
		.INIT('h9669)
	) name9381 (
		_w8946_,
		_w8947_,
		_w8951_,
		_w9175_,
		_w9415_
	);
	LUT4 #(
		.INIT('h5060)
	) name9382 (
		_w3409_,
		_w3650_,
		_w3709_,
		_w6959_,
		_w9416_
	);
	LUT4 #(
		.INIT('h007d)
	) name9383 (
		_w3877_,
		_w6960_,
		_w6962_,
		_w9416_,
		_w9417_
	);
	LUT3 #(
		.INIT('h70)
	) name9384 (
		_w3886_,
		_w7014_,
		_w9417_,
		_w9418_
	);
	LUT4 #(
		.INIT('h95aa)
	) name9385 (
		\a[17] ,
		_w3710_,
		_w7291_,
		_w9418_,
		_w9419_
	);
	LUT4 #(
		.INIT('hde48)
	) name9386 (
		_w9181_,
		_w9414_,
		_w9415_,
		_w9419_,
		_w9420_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9387 (
		_w4034_,
		_w7010_,
		_w7121_,
		_w7122_,
		_w9421_
	);
	LUT4 #(
		.INIT('h04c8)
	) name9388 (
		_w2983_,
		_w4382_,
		_w6972_,
		_w6974_,
		_w9422_
	);
	LUT3 #(
		.INIT('h82)
	) name9389 (
		_w4033_,
		_w6967_,
		_w6969_,
		_w9423_
	);
	LUT3 #(
		.INIT('h07)
	) name9390 (
		_w4367_,
		_w7008_,
		_w9423_,
		_w9424_
	);
	LUT2 #(
		.INIT('h4)
	) name9391 (
		_w9422_,
		_w9424_,
		_w9425_
	);
	LUT3 #(
		.INIT('h9a)
	) name9392 (
		\a[14] ,
		_w9421_,
		_w9425_,
		_w9426_
	);
	LUT3 #(
		.INIT('hd4)
	) name9393 (
		_w9220_,
		_w9420_,
		_w9426_,
		_w9427_
	);
	LUT3 #(
		.INIT('h82)
	) name9394 (
		_w4459_,
		_w7129_,
		_w7131_,
		_w9428_
	);
	LUT3 #(
		.INIT('h84)
	) name9395 (
		_w2546_,
		_w4700_,
		_w6981_,
		_w9429_
	);
	LUT2 #(
		.INIT('h8)
	) name9396 (
		_w4458_,
		_w7002_,
		_w9430_
	);
	LUT4 #(
		.INIT('h04c8)
	) name9397 (
		_w2622_,
		_w4684_,
		_w6978_,
		_w6980_,
		_w9431_
	);
	LUT2 #(
		.INIT('h1)
	) name9398 (
		_w9430_,
		_w9431_,
		_w9432_
	);
	LUT2 #(
		.INIT('h4)
	) name9399 (
		_w9429_,
		_w9432_,
		_w9433_
	);
	LUT3 #(
		.INIT('h9a)
	) name9400 (
		\a[11] ,
		_w9428_,
		_w9433_,
		_w9434_
	);
	LUT4 #(
		.INIT('hf660)
	) name9401 (
		_w9198_,
		_w9219_,
		_w9427_,
		_w9434_,
		_w9435_
	);
	LUT4 #(
		.INIT('hf660)
	) name9402 (
		_w9007_,
		_w9199_,
		_w9218_,
		_w9435_,
		_w9436_
	);
	LUT4 #(
		.INIT('h0096)
	) name9403 (
		_w9200_,
		_w9201_,
		_w9207_,
		_w9436_,
		_w9437_
	);
	LUT4 #(
		.INIT('h6900)
	) name9404 (
		_w9200_,
		_w9201_,
		_w9207_,
		_w9436_,
		_w9438_
	);
	LUT4 #(
		.INIT('h0a02)
	) name9405 (
		_w4876_,
		_w7169_,
		_w7419_,
		_w7686_,
		_w9439_
	);
	LUT3 #(
		.INIT('h28)
	) name9406 (
		_w4875_,
		_w7136_,
		_w7168_,
		_w9440_
	);
	LUT3 #(
		.INIT('h40)
	) name9407 (
		_w5286_,
		_w7136_,
		_w7167_,
		_w9441_
	);
	LUT3 #(
		.INIT('h31)
	) name9408 (
		_w8997_,
		_w9440_,
		_w9441_,
		_w9442_
	);
	LUT3 #(
		.INIT('h9a)
	) name9409 (
		\a[8] ,
		_w9439_,
		_w9442_,
		_w9443_
	);
	LUT3 #(
		.INIT('h54)
	) name9410 (
		_w9437_,
		_w9438_,
		_w9443_,
		_w9444_
	);
	LUT2 #(
		.INIT('h2)
	) name9411 (
		_w9214_,
		_w9444_,
		_w9445_
	);
	LUT2 #(
		.INIT('h9)
	) name9412 (
		_w9214_,
		_w9444_,
		_w9446_
	);
	LUT3 #(
		.INIT('h28)
	) name9413 (
		_w5271_,
		_w7136_,
		_w7168_,
		_w9447_
	);
	LUT4 #(
		.INIT('h028a)
	) name9414 (
		_w5286_,
		_w7136_,
		_w7166_,
		_w7167_,
		_w9448_
	);
	LUT4 #(
		.INIT('h04c8)
	) name9415 (
		_w2411_,
		_w4875_,
		_w6983_,
		_w6993_,
		_w9449_
	);
	LUT3 #(
		.INIT('h01)
	) name9416 (
		_w9448_,
		_w9449_,
		_w9447_,
		_w9450_
	);
	LUT4 #(
		.INIT('h95aa)
	) name9417 (
		\a[8] ,
		_w4876_,
		_w7696_,
		_w9450_,
		_w9451_
	);
	LUT4 #(
		.INIT('h9669)
	) name9418 (
		_w9198_,
		_w9219_,
		_w9427_,
		_w9434_,
		_w9452_
	);
	LUT3 #(
		.INIT('h82)
	) name9419 (
		_w3710_,
		_w7111_,
		_w7113_,
		_w9453_
	);
	LUT3 #(
		.INIT('h82)
	) name9420 (
		_w3886_,
		_w6960_,
		_w6962_,
		_w9454_
	);
	LUT2 #(
		.INIT('h8)
	) name9421 (
		_w3709_,
		_w7020_,
		_w9455_
	);
	LUT4 #(
		.INIT('h5060)
	) name9422 (
		_w3409_,
		_w3650_,
		_w3877_,
		_w6959_,
		_w9456_
	);
	LUT2 #(
		.INIT('h1)
	) name9423 (
		_w9455_,
		_w9456_,
		_w9457_
	);
	LUT2 #(
		.INIT('h4)
	) name9424 (
		_w9454_,
		_w9457_,
		_w9458_
	);
	LUT3 #(
		.INIT('h1e)
	) name9425 (
		_w9235_,
		_w9412_,
		_w9413_,
		_w9459_
	);
	LUT4 #(
		.INIT('h6500)
	) name9426 (
		\a[17] ,
		_w9453_,
		_w9458_,
		_w9459_,
		_w9460_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9427 (
		_w3710_,
		_w7022_,
		_w7109_,
		_w7110_,
		_w9461_
	);
	LUT4 #(
		.INIT('h5060)
	) name9428 (
		_w3409_,
		_w3650_,
		_w3886_,
		_w6959_,
		_w9462_
	);
	LUT3 #(
		.INIT('h84)
	) name9429 (
		_w3706_,
		_w3709_,
		_w6957_,
		_w9463_
	);
	LUT3 #(
		.INIT('h07)
	) name9430 (
		_w3877_,
		_w7020_,
		_w9463_,
		_w9464_
	);
	LUT2 #(
		.INIT('h4)
	) name9431 (
		_w9462_,
		_w9464_,
		_w9465_
	);
	LUT4 #(
		.INIT('h54ab)
	) name9432 (
		_w9241_,
		_w9408_,
		_w9409_,
		_w9411_,
		_w9466_
	);
	LUT4 #(
		.INIT('h6500)
	) name9433 (
		\a[17] ,
		_w9461_,
		_w9465_,
		_w9466_,
		_w9467_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9434 (
		_w3709_,
		_w3882_,
		_w6954_,
		_w6956_,
		_w9468_
	);
	LUT4 #(
		.INIT('h007b)
	) name9435 (
		_w3706_,
		_w3877_,
		_w6957_,
		_w9468_,
		_w9469_
	);
	LUT3 #(
		.INIT('h70)
	) name9436 (
		_w3886_,
		_w7020_,
		_w9469_,
		_w9470_
	);
	LUT4 #(
		.INIT('h95aa)
	) name9437 (
		\a[17] ,
		_w3710_,
		_w7465_,
		_w9470_,
		_w9471_
	);
	LUT2 #(
		.INIT('h9)
	) name9438 (
		_w9408_,
		_w9410_,
		_w9472_
	);
	LUT2 #(
		.INIT('h4)
	) name9439 (
		_w9471_,
		_w9472_,
		_w9473_
	);
	LUT3 #(
		.INIT('h82)
	) name9440 (
		_w3710_,
		_w7105_,
		_w7107_,
		_w9474_
	);
	LUT3 #(
		.INIT('h84)
	) name9441 (
		_w3706_,
		_w3886_,
		_w6957_,
		_w9475_
	);
	LUT2 #(
		.INIT('h8)
	) name9442 (
		_w3709_,
		_w7026_,
		_w9476_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9443 (
		_w3877_,
		_w3882_,
		_w6954_,
		_w6956_,
		_w9477_
	);
	LUT2 #(
		.INIT('h1)
	) name9444 (
		_w9476_,
		_w9477_,
		_w9478_
	);
	LUT2 #(
		.INIT('h4)
	) name9445 (
		_w9475_,
		_w9478_,
		_w9479_
	);
	LUT3 #(
		.INIT('h1e)
	) name9446 (
		_w9256_,
		_w9406_,
		_w9407_,
		_w9480_
	);
	LUT4 #(
		.INIT('h6500)
	) name9447 (
		\a[17] ,
		_w9474_,
		_w9479_,
		_w9480_,
		_w9481_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9448 (
		_w3710_,
		_w7028_,
		_w7103_,
		_w7104_,
		_w9482_
	);
	LUT4 #(
		.INIT('h04c8)
	) name9449 (
		_w3882_,
		_w3886_,
		_w6954_,
		_w6956_,
		_w9483_
	);
	LUT3 #(
		.INIT('h82)
	) name9450 (
		_w3709_,
		_w4030_,
		_w6952_,
		_w9484_
	);
	LUT3 #(
		.INIT('h07)
	) name9451 (
		_w3877_,
		_w7026_,
		_w9484_,
		_w9485_
	);
	LUT2 #(
		.INIT('h4)
	) name9452 (
		_w9483_,
		_w9485_,
		_w9486_
	);
	LUT4 #(
		.INIT('h54ab)
	) name9453 (
		_w9262_,
		_w9402_,
		_w9403_,
		_w9405_,
		_w9487_
	);
	LUT4 #(
		.INIT('h6500)
	) name9454 (
		\a[17] ,
		_w9482_,
		_w9486_,
		_w9487_,
		_w9488_
	);
	LUT4 #(
		.INIT('h2228)
	) name9455 (
		_w3709_,
		_w4099_,
		_w4378_,
		_w6951_,
		_w9489_
	);
	LUT4 #(
		.INIT('h007d)
	) name9456 (
		_w3877_,
		_w4030_,
		_w6952_,
		_w9489_,
		_w9490_
	);
	LUT3 #(
		.INIT('h70)
	) name9457 (
		_w3886_,
		_w7026_,
		_w9490_,
		_w9491_
	);
	LUT4 #(
		.INIT('h95aa)
	) name9458 (
		\a[17] ,
		_w3710_,
		_w7562_,
		_w9491_,
		_w9492_
	);
	LUT2 #(
		.INIT('h9)
	) name9459 (
		_w9402_,
		_w9404_,
		_w9493_
	);
	LUT2 #(
		.INIT('h4)
	) name9460 (
		_w9492_,
		_w9493_,
		_w9494_
	);
	LUT3 #(
		.INIT('h82)
	) name9461 (
		_w3710_,
		_w7099_,
		_w7101_,
		_w9495_
	);
	LUT3 #(
		.INIT('h82)
	) name9462 (
		_w3886_,
		_w4030_,
		_w6952_,
		_w9496_
	);
	LUT2 #(
		.INIT('h8)
	) name9463 (
		_w3709_,
		_w7032_,
		_w9497_
	);
	LUT4 #(
		.INIT('h2228)
	) name9464 (
		_w3877_,
		_w4099_,
		_w4378_,
		_w6951_,
		_w9498_
	);
	LUT2 #(
		.INIT('h1)
	) name9465 (
		_w9497_,
		_w9498_,
		_w9499_
	);
	LUT2 #(
		.INIT('h4)
	) name9466 (
		_w9496_,
		_w9499_,
		_w9500_
	);
	LUT3 #(
		.INIT('h1e)
	) name9467 (
		_w9277_,
		_w9400_,
		_w9401_,
		_w9501_
	);
	LUT4 #(
		.INIT('h6500)
	) name9468 (
		\a[17] ,
		_w9495_,
		_w9500_,
		_w9501_,
		_w9502_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9469 (
		_w3710_,
		_w7034_,
		_w7097_,
		_w7098_,
		_w9503_
	);
	LUT4 #(
		.INIT('h2228)
	) name9470 (
		_w3886_,
		_w4099_,
		_w4378_,
		_w6951_,
		_w9504_
	);
	LUT3 #(
		.INIT('h82)
	) name9471 (
		_w3709_,
		_w6947_,
		_w6949_,
		_w9505_
	);
	LUT3 #(
		.INIT('h07)
	) name9472 (
		_w3877_,
		_w7032_,
		_w9505_,
		_w9506_
	);
	LUT2 #(
		.INIT('h4)
	) name9473 (
		_w9504_,
		_w9506_,
		_w9507_
	);
	LUT4 #(
		.INIT('h54ab)
	) name9474 (
		_w9283_,
		_w9396_,
		_w9397_,
		_w9399_,
		_w9508_
	);
	LUT4 #(
		.INIT('h6500)
	) name9475 (
		\a[17] ,
		_w9503_,
		_w9507_,
		_w9508_,
		_w9509_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9476 (
		_w3709_,
		_w4695_,
		_w6944_,
		_w6946_,
		_w9510_
	);
	LUT4 #(
		.INIT('h007d)
	) name9477 (
		_w3877_,
		_w6947_,
		_w6949_,
		_w9510_,
		_w9511_
	);
	LUT3 #(
		.INIT('h70)
	) name9478 (
		_w3886_,
		_w7032_,
		_w9511_,
		_w9512_
	);
	LUT4 #(
		.INIT('h95aa)
	) name9479 (
		\a[17] ,
		_w3710_,
		_w7882_,
		_w9512_,
		_w9513_
	);
	LUT2 #(
		.INIT('h9)
	) name9480 (
		_w9396_,
		_w9398_,
		_w9514_
	);
	LUT2 #(
		.INIT('h4)
	) name9481 (
		_w9513_,
		_w9514_,
		_w9515_
	);
	LUT3 #(
		.INIT('h82)
	) name9482 (
		_w3710_,
		_w7093_,
		_w7095_,
		_w9516_
	);
	LUT3 #(
		.INIT('h82)
	) name9483 (
		_w3886_,
		_w6947_,
		_w6949_,
		_w9517_
	);
	LUT2 #(
		.INIT('h8)
	) name9484 (
		_w3709_,
		_w7038_,
		_w9518_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9485 (
		_w3877_,
		_w4695_,
		_w6944_,
		_w6946_,
		_w9519_
	);
	LUT2 #(
		.INIT('h1)
	) name9486 (
		_w9518_,
		_w9519_,
		_w9520_
	);
	LUT2 #(
		.INIT('h4)
	) name9487 (
		_w9517_,
		_w9520_,
		_w9521_
	);
	LUT3 #(
		.INIT('h1e)
	) name9488 (
		_w9298_,
		_w9394_,
		_w9395_,
		_w9522_
	);
	LUT4 #(
		.INIT('h6500)
	) name9489 (
		\a[17] ,
		_w9516_,
		_w9521_,
		_w9522_,
		_w9523_
	);
	LUT4 #(
		.INIT('h54ab)
	) name9490 (
		_w9304_,
		_w9390_,
		_w9391_,
		_w9393_,
		_w9524_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9491 (
		_w3710_,
		_w7040_,
		_w7091_,
		_w7092_,
		_w9525_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9492 (
		_w3886_,
		_w4695_,
		_w6944_,
		_w6946_,
		_w9526_
	);
	LUT3 #(
		.INIT('h82)
	) name9493 (
		_w3709_,
		_w6940_,
		_w6942_,
		_w9527_
	);
	LUT3 #(
		.INIT('h07)
	) name9494 (
		_w3877_,
		_w7038_,
		_w9527_,
		_w9528_
	);
	LUT2 #(
		.INIT('h4)
	) name9495 (
		_w9526_,
		_w9528_,
		_w9529_
	);
	LUT4 #(
		.INIT('h4844)
	) name9496 (
		\a[17] ,
		_w9524_,
		_w9525_,
		_w9529_,
		_w9530_
	);
	LUT2 #(
		.INIT('h9)
	) name9497 (
		_w9390_,
		_w9392_,
		_w9531_
	);
	LUT4 #(
		.INIT('h2228)
	) name9498 (
		_w3709_,
		_w5067_,
		_w5282_,
		_w6939_,
		_w9532_
	);
	LUT4 #(
		.INIT('h007d)
	) name9499 (
		_w3877_,
		_w6940_,
		_w6942_,
		_w9532_,
		_w9533_
	);
	LUT3 #(
		.INIT('h70)
	) name9500 (
		_w3886_,
		_w7038_,
		_w9533_,
		_w9534_
	);
	LUT4 #(
		.INIT('h95aa)
	) name9501 (
		\a[17] ,
		_w3710_,
		_w8018_,
		_w9534_,
		_w9535_
	);
	LUT2 #(
		.INIT('h2)
	) name9502 (
		_w9531_,
		_w9535_,
		_w9536_
	);
	LUT3 #(
		.INIT('h82)
	) name9503 (
		_w3710_,
		_w7087_,
		_w7089_,
		_w9537_
	);
	LUT3 #(
		.INIT('h82)
	) name9504 (
		_w3886_,
		_w6940_,
		_w6942_,
		_w9538_
	);
	LUT2 #(
		.INIT('h8)
	) name9505 (
		_w3709_,
		_w7044_,
		_w9539_
	);
	LUT4 #(
		.INIT('h2228)
	) name9506 (
		_w3877_,
		_w5067_,
		_w5282_,
		_w6939_,
		_w9540_
	);
	LUT2 #(
		.INIT('h1)
	) name9507 (
		_w9539_,
		_w9540_,
		_w9541_
	);
	LUT2 #(
		.INIT('h4)
	) name9508 (
		_w9538_,
		_w9541_,
		_w9542_
	);
	LUT3 #(
		.INIT('h1e)
	) name9509 (
		_w9319_,
		_w9388_,
		_w9389_,
		_w9543_
	);
	LUT4 #(
		.INIT('h6500)
	) name9510 (
		\a[17] ,
		_w9537_,
		_w9542_,
		_w9543_,
		_w9544_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9511 (
		_w3710_,
		_w7046_,
		_w7085_,
		_w7086_,
		_w9545_
	);
	LUT4 #(
		.INIT('h2228)
	) name9512 (
		_w3886_,
		_w5067_,
		_w5282_,
		_w6939_,
		_w9546_
	);
	LUT3 #(
		.INIT('h82)
	) name9513 (
		_w3709_,
		_w6935_,
		_w6937_,
		_w9547_
	);
	LUT3 #(
		.INIT('h07)
	) name9514 (
		_w3877_,
		_w7044_,
		_w9547_,
		_w9548_
	);
	LUT2 #(
		.INIT('h4)
	) name9515 (
		_w9546_,
		_w9548_,
		_w9549_
	);
	LUT4 #(
		.INIT('h54ab)
	) name9516 (
		_w9325_,
		_w9384_,
		_w9385_,
		_w9387_,
		_w9550_
	);
	LUT4 #(
		.INIT('h6500)
	) name9517 (
		\a[17] ,
		_w9545_,
		_w9549_,
		_w9550_,
		_w9551_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9518 (
		_w3709_,
		_w6043_,
		_w6933_,
		_w6934_,
		_w9552_
	);
	LUT4 #(
		.INIT('h007d)
	) name9519 (
		_w3877_,
		_w6935_,
		_w6937_,
		_w9552_,
		_w9553_
	);
	LUT3 #(
		.INIT('h70)
	) name9520 (
		_w3886_,
		_w7044_,
		_w9553_,
		_w9554_
	);
	LUT4 #(
		.INIT('h95aa)
	) name9521 (
		\a[17] ,
		_w3710_,
		_w8005_,
		_w9554_,
		_w9555_
	);
	LUT2 #(
		.INIT('h9)
	) name9522 (
		_w9384_,
		_w9386_,
		_w9556_
	);
	LUT2 #(
		.INIT('h4)
	) name9523 (
		_w9555_,
		_w9556_,
		_w9557_
	);
	LUT3 #(
		.INIT('h1e)
	) name9524 (
		_w9340_,
		_w9382_,
		_w9383_,
		_w9558_
	);
	LUT3 #(
		.INIT('h82)
	) name9525 (
		_w3710_,
		_w7081_,
		_w7083_,
		_w9559_
	);
	LUT3 #(
		.INIT('h82)
	) name9526 (
		_w3886_,
		_w6935_,
		_w6937_,
		_w9560_
	);
	LUT2 #(
		.INIT('h8)
	) name9527 (
		_w3709_,
		_w7050_,
		_w9561_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9528 (
		_w3877_,
		_w6043_,
		_w6933_,
		_w6934_,
		_w9562_
	);
	LUT2 #(
		.INIT('h1)
	) name9529 (
		_w9561_,
		_w9562_,
		_w9563_
	);
	LUT2 #(
		.INIT('h4)
	) name9530 (
		_w9560_,
		_w9563_,
		_w9564_
	);
	LUT4 #(
		.INIT('h4844)
	) name9531 (
		\a[17] ,
		_w9558_,
		_w9559_,
		_w9564_,
		_w9565_
	);
	LUT4 #(
		.INIT('h54ab)
	) name9532 (
		_w9347_,
		_w9378_,
		_w9379_,
		_w9381_,
		_w9566_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9533 (
		_w3710_,
		_w7052_,
		_w7079_,
		_w7080_,
		_w9567_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9534 (
		_w3886_,
		_w6043_,
		_w6933_,
		_w6934_,
		_w9568_
	);
	LUT3 #(
		.INIT('h82)
	) name9535 (
		_w3709_,
		_w6929_,
		_w6931_,
		_w9569_
	);
	LUT3 #(
		.INIT('h07)
	) name9536 (
		_w3877_,
		_w7050_,
		_w9569_,
		_w9570_
	);
	LUT2 #(
		.INIT('h4)
	) name9537 (
		_w9568_,
		_w9570_,
		_w9571_
	);
	LUT4 #(
		.INIT('h4844)
	) name9538 (
		\a[17] ,
		_w9566_,
		_w9567_,
		_w9571_,
		_w9572_
	);
	LUT2 #(
		.INIT('h9)
	) name9539 (
		_w9378_,
		_w9380_,
		_w9573_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9540 (
		_w3709_,
		_w6645_,
		_w6926_,
		_w6928_,
		_w9574_
	);
	LUT4 #(
		.INIT('h007d)
	) name9541 (
		_w3877_,
		_w6929_,
		_w6931_,
		_w9574_,
		_w9575_
	);
	LUT3 #(
		.INIT('h70)
	) name9542 (
		_w3886_,
		_w7050_,
		_w9575_,
		_w9576_
	);
	LUT4 #(
		.INIT('h95aa)
	) name9543 (
		\a[17] ,
		_w3710_,
		_w8227_,
		_w9576_,
		_w9577_
	);
	LUT2 #(
		.INIT('h2)
	) name9544 (
		_w9573_,
		_w9577_,
		_w9578_
	);
	LUT3 #(
		.INIT('h82)
	) name9545 (
		_w3710_,
		_w7075_,
		_w7077_,
		_w9579_
	);
	LUT3 #(
		.INIT('h82)
	) name9546 (
		_w3886_,
		_w6929_,
		_w6931_,
		_w9580_
	);
	LUT2 #(
		.INIT('h8)
	) name9547 (
		_w3709_,
		_w7056_,
		_w9581_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9548 (
		_w3877_,
		_w6645_,
		_w6926_,
		_w6928_,
		_w9582_
	);
	LUT2 #(
		.INIT('h1)
	) name9549 (
		_w9581_,
		_w9582_,
		_w9583_
	);
	LUT2 #(
		.INIT('h4)
	) name9550 (
		_w9580_,
		_w9583_,
		_w9584_
	);
	LUT2 #(
		.INIT('h9)
	) name9551 (
		_w9375_,
		_w9377_,
		_w9585_
	);
	LUT4 #(
		.INIT('h6500)
	) name9552 (
		\a[17] ,
		_w9579_,
		_w9584_,
		_w9585_,
		_w9586_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9553 (
		_w3710_,
		_w7058_,
		_w7073_,
		_w7074_,
		_w9587_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9554 (
		_w3886_,
		_w6645_,
		_w6926_,
		_w6928_,
		_w9588_
	);
	LUT3 #(
		.INIT('h82)
	) name9555 (
		_w3709_,
		_w6922_,
		_w6924_,
		_w9589_
	);
	LUT3 #(
		.INIT('h07)
	) name9556 (
		_w3877_,
		_w7056_,
		_w9589_,
		_w9590_
	);
	LUT2 #(
		.INIT('h4)
	) name9557 (
		_w9588_,
		_w9590_,
		_w9591_
	);
	LUT4 #(
		.INIT('h9a65)
	) name9558 (
		\a[20] ,
		_w9368_,
		_w9372_,
		_w9373_,
		_w9592_
	);
	LUT4 #(
		.INIT('h6500)
	) name9559 (
		\a[17] ,
		_w9587_,
		_w9591_,
		_w9592_,
		_w9593_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9560 (
		_w3709_,
		_w6669_,
		_w6919_,
		_w6921_,
		_w9594_
	);
	LUT4 #(
		.INIT('h007d)
	) name9561 (
		_w3877_,
		_w6922_,
		_w6924_,
		_w9594_,
		_w9595_
	);
	LUT3 #(
		.INIT('h70)
	) name9562 (
		_w3886_,
		_w7056_,
		_w9595_,
		_w9596_
	);
	LUT4 #(
		.INIT('h95aa)
	) name9563 (
		\a[17] ,
		_w3710_,
		_w8298_,
		_w9596_,
		_w9597_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name9564 (
		\a[20] ,
		_w9360_,
		_w9357_,
		_w9359_,
		_w9598_
	);
	LUT3 #(
		.INIT('h4b)
	) name9565 (
		_w9363_,
		_w9366_,
		_w9598_,
		_w9599_
	);
	LUT2 #(
		.INIT('h4)
	) name9566 (
		_w9597_,
		_w9599_,
		_w9600_
	);
	LUT3 #(
		.INIT('h82)
	) name9567 (
		_w3710_,
		_w7069_,
		_w7071_,
		_w9601_
	);
	LUT3 #(
		.INIT('h82)
	) name9568 (
		_w3886_,
		_w6922_,
		_w6924_,
		_w9602_
	);
	LUT2 #(
		.INIT('h8)
	) name9569 (
		_w3709_,
		_w7062_,
		_w9603_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9570 (
		_w3877_,
		_w6669_,
		_w6919_,
		_w6921_,
		_w9604_
	);
	LUT2 #(
		.INIT('h1)
	) name9571 (
		_w9603_,
		_w9604_,
		_w9605_
	);
	LUT2 #(
		.INIT('h4)
	) name9572 (
		_w9602_,
		_w9605_,
		_w9606_
	);
	LUT2 #(
		.INIT('h8)
	) name9573 (
		\a[20] ,
		_w9360_,
		_w9607_
	);
	LUT3 #(
		.INIT('h4b)
	) name9574 (
		_w9357_,
		_w9359_,
		_w9607_,
		_w9608_
	);
	LUT4 #(
		.INIT('h6500)
	) name9575 (
		\a[17] ,
		_w9601_,
		_w9606_,
		_w9608_,
		_w9609_
	);
	LUT4 #(
		.INIT('h2882)
	) name9576 (
		_w3710_,
		_w6914_,
		_w6916_,
		_w7067_,
		_w9610_
	);
	LUT4 #(
		.INIT('ha802)
	) name9577 (
		_w3877_,
		_w6689_,
		_w6911_,
		_w6913_,
		_w9611_
	);
	LUT4 #(
		.INIT('h007d)
	) name9578 (
		_w3886_,
		_w6914_,
		_w6916_,
		_w9611_,
		_w9612_
	);
	LUT4 #(
		.INIT('h5401)
	) name9579 (
		_w3708_,
		_w6689_,
		_w6911_,
		_w6913_,
		_w9613_
	);
	LUT2 #(
		.INIT('h2)
	) name9580 (
		\a[17] ,
		_w9613_,
		_w9614_
	);
	LUT3 #(
		.INIT('h40)
	) name9581 (
		_w9610_,
		_w9612_,
		_w9614_,
		_w9615_
	);
	LUT3 #(
		.INIT('h28)
	) name9582 (
		_w3710_,
		_w7062_,
		_w8358_,
		_w9616_
	);
	LUT4 #(
		.INIT('ha802)
	) name9583 (
		_w3709_,
		_w6689_,
		_w6911_,
		_w6913_,
		_w9617_
	);
	LUT4 #(
		.INIT('h007d)
	) name9584 (
		_w3877_,
		_w6914_,
		_w6916_,
		_w9617_,
		_w9618_
	);
	LUT3 #(
		.INIT('h70)
	) name9585 (
		_w3886_,
		_w7062_,
		_w9618_,
		_w9619_
	);
	LUT4 #(
		.INIT('h0800)
	) name9586 (
		_w9360_,
		_w9615_,
		_w9616_,
		_w9619_,
		_w9620_
	);
	LUT3 #(
		.INIT('h28)
	) name9587 (
		_w3710_,
		_w7065_,
		_w7068_,
		_w9621_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9588 (
		_w3886_,
		_w6669_,
		_w6919_,
		_w6921_,
		_w9622_
	);
	LUT3 #(
		.INIT('h82)
	) name9589 (
		_w3709_,
		_w6914_,
		_w6916_,
		_w9623_
	);
	LUT3 #(
		.INIT('h07)
	) name9590 (
		_w3877_,
		_w7062_,
		_w9623_,
		_w9624_
	);
	LUT2 #(
		.INIT('h4)
	) name9591 (
		_w9622_,
		_w9624_,
		_w9625_
	);
	LUT4 #(
		.INIT('ha6aa)
	) name9592 (
		_w9360_,
		_w9615_,
		_w9616_,
		_w9619_,
		_w9626_
	);
	LUT4 #(
		.INIT('h6500)
	) name9593 (
		\a[17] ,
		_w9621_,
		_w9625_,
		_w9626_,
		_w9627_
	);
	LUT2 #(
		.INIT('h1)
	) name9594 (
		_w9620_,
		_w9627_,
		_w9628_
	);
	LUT4 #(
		.INIT('h009a)
	) name9595 (
		\a[17] ,
		_w9601_,
		_w9606_,
		_w9608_,
		_w9629_
	);
	LUT4 #(
		.INIT('h9a65)
	) name9596 (
		\a[17] ,
		_w9601_,
		_w9606_,
		_w9608_,
		_w9630_
	);
	LUT3 #(
		.INIT('h54)
	) name9597 (
		_w9609_,
		_w9628_,
		_w9629_,
		_w9631_
	);
	LUT2 #(
		.INIT('h2)
	) name9598 (
		_w9597_,
		_w9599_,
		_w9632_
	);
	LUT2 #(
		.INIT('h9)
	) name9599 (
		_w9597_,
		_w9599_,
		_w9633_
	);
	LUT4 #(
		.INIT('h9a65)
	) name9600 (
		\a[17] ,
		_w9587_,
		_w9591_,
		_w9592_,
		_w9634_
	);
	LUT4 #(
		.INIT('h4d00)
	) name9601 (
		_w9597_,
		_w9599_,
		_w9631_,
		_w9634_,
		_w9635_
	);
	LUT4 #(
		.INIT('h9a65)
	) name9602 (
		\a[17] ,
		_w9579_,
		_w9584_,
		_w9585_,
		_w9636_
	);
	LUT4 #(
		.INIT('h0155)
	) name9603 (
		_w9586_,
		_w9593_,
		_w9635_,
		_w9636_,
		_w9637_
	);
	LUT2 #(
		.INIT('h4)
	) name9604 (
		_w9573_,
		_w9577_,
		_w9638_
	);
	LUT2 #(
		.INIT('h9)
	) name9605 (
		_w9573_,
		_w9577_,
		_w9639_
	);
	LUT4 #(
		.INIT('h9699)
	) name9606 (
		\a[17] ,
		_w9566_,
		_w9567_,
		_w9571_,
		_w9640_
	);
	LUT4 #(
		.INIT('h2b00)
	) name9607 (
		_w9573_,
		_w9577_,
		_w9637_,
		_w9640_,
		_w9641_
	);
	LUT4 #(
		.INIT('h9699)
	) name9608 (
		\a[17] ,
		_w9558_,
		_w9559_,
		_w9564_,
		_w9642_
	);
	LUT4 #(
		.INIT('h0155)
	) name9609 (
		_w9565_,
		_w9572_,
		_w9641_,
		_w9642_,
		_w9643_
	);
	LUT2 #(
		.INIT('h2)
	) name9610 (
		_w9555_,
		_w9556_,
		_w9644_
	);
	LUT2 #(
		.INIT('h9)
	) name9611 (
		_w9555_,
		_w9556_,
		_w9645_
	);
	LUT4 #(
		.INIT('h9a65)
	) name9612 (
		\a[17] ,
		_w9545_,
		_w9549_,
		_w9550_,
		_w9646_
	);
	LUT4 #(
		.INIT('h4d00)
	) name9613 (
		_w9555_,
		_w9556_,
		_w9643_,
		_w9646_,
		_w9647_
	);
	LUT4 #(
		.INIT('h9a65)
	) name9614 (
		\a[17] ,
		_w9537_,
		_w9542_,
		_w9543_,
		_w9648_
	);
	LUT4 #(
		.INIT('h0155)
	) name9615 (
		_w9544_,
		_w9551_,
		_w9647_,
		_w9648_,
		_w9649_
	);
	LUT2 #(
		.INIT('h4)
	) name9616 (
		_w9531_,
		_w9535_,
		_w9650_
	);
	LUT2 #(
		.INIT('h9)
	) name9617 (
		_w9531_,
		_w9535_,
		_w9651_
	);
	LUT4 #(
		.INIT('h9699)
	) name9618 (
		\a[17] ,
		_w9524_,
		_w9525_,
		_w9529_,
		_w9652_
	);
	LUT4 #(
		.INIT('h2b00)
	) name9619 (
		_w9531_,
		_w9535_,
		_w9649_,
		_w9652_,
		_w9653_
	);
	LUT4 #(
		.INIT('h9a65)
	) name9620 (
		\a[17] ,
		_w9516_,
		_w9521_,
		_w9522_,
		_w9654_
	);
	LUT4 #(
		.INIT('h0155)
	) name9621 (
		_w9523_,
		_w9530_,
		_w9653_,
		_w9654_,
		_w9655_
	);
	LUT2 #(
		.INIT('h2)
	) name9622 (
		_w9513_,
		_w9514_,
		_w9656_
	);
	LUT2 #(
		.INIT('h9)
	) name9623 (
		_w9513_,
		_w9514_,
		_w9657_
	);
	LUT4 #(
		.INIT('h9a65)
	) name9624 (
		\a[17] ,
		_w9503_,
		_w9507_,
		_w9508_,
		_w9658_
	);
	LUT4 #(
		.INIT('h4d00)
	) name9625 (
		_w9513_,
		_w9514_,
		_w9655_,
		_w9658_,
		_w9659_
	);
	LUT4 #(
		.INIT('h9a65)
	) name9626 (
		\a[17] ,
		_w9495_,
		_w9500_,
		_w9501_,
		_w9660_
	);
	LUT4 #(
		.INIT('h0155)
	) name9627 (
		_w9502_,
		_w9509_,
		_w9659_,
		_w9660_,
		_w9661_
	);
	LUT2 #(
		.INIT('h2)
	) name9628 (
		_w9492_,
		_w9493_,
		_w9662_
	);
	LUT2 #(
		.INIT('h9)
	) name9629 (
		_w9492_,
		_w9493_,
		_w9663_
	);
	LUT4 #(
		.INIT('h9a65)
	) name9630 (
		\a[17] ,
		_w9482_,
		_w9486_,
		_w9487_,
		_w9664_
	);
	LUT4 #(
		.INIT('h4d00)
	) name9631 (
		_w9492_,
		_w9493_,
		_w9661_,
		_w9664_,
		_w9665_
	);
	LUT4 #(
		.INIT('h9a65)
	) name9632 (
		\a[17] ,
		_w9474_,
		_w9479_,
		_w9480_,
		_w9666_
	);
	LUT4 #(
		.INIT('h0155)
	) name9633 (
		_w9481_,
		_w9488_,
		_w9665_,
		_w9666_,
		_w9667_
	);
	LUT2 #(
		.INIT('h2)
	) name9634 (
		_w9471_,
		_w9472_,
		_w9668_
	);
	LUT2 #(
		.INIT('h9)
	) name9635 (
		_w9471_,
		_w9472_,
		_w9669_
	);
	LUT4 #(
		.INIT('h9a65)
	) name9636 (
		\a[17] ,
		_w9461_,
		_w9465_,
		_w9466_,
		_w9670_
	);
	LUT4 #(
		.INIT('h4d00)
	) name9637 (
		_w9471_,
		_w9472_,
		_w9667_,
		_w9670_,
		_w9671_
	);
	LUT4 #(
		.INIT('h9a65)
	) name9638 (
		\a[17] ,
		_w9453_,
		_w9458_,
		_w9459_,
		_w9672_
	);
	LUT4 #(
		.INIT('h0155)
	) name9639 (
		_w9460_,
		_w9467_,
		_w9671_,
		_w9672_,
		_w9673_
	);
	LUT4 #(
		.INIT('h6996)
	) name9640 (
		_w9181_,
		_w9414_,
		_w9415_,
		_w9419_,
		_w9674_
	);
	LUT4 #(
		.INIT('h04c8)
	) name9641 (
		_w3257_,
		_w4033_,
		_w6964_,
		_w6966_,
		_w9675_
	);
	LUT4 #(
		.INIT('h007d)
	) name9642 (
		_w4367_,
		_w6967_,
		_w6969_,
		_w9675_,
		_w9676_
	);
	LUT3 #(
		.INIT('h70)
	) name9643 (
		_w4382_,
		_w7008_,
		_w9676_,
		_w9677_
	);
	LUT4 #(
		.INIT('h95aa)
	) name9644 (
		\a[14] ,
		_w4034_,
		_w7403_,
		_w9677_,
		_w9678_
	);
	LUT3 #(
		.INIT('he8)
	) name9645 (
		_w9673_,
		_w9674_,
		_w9678_,
		_w9679_
	);
	LUT4 #(
		.INIT('h0096)
	) name9646 (
		_w9220_,
		_w9420_,
		_w9426_,
		_w9679_,
		_w9680_
	);
	LUT4 #(
		.INIT('h6900)
	) name9647 (
		_w9220_,
		_w9420_,
		_w9426_,
		_w9679_,
		_w9681_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9648 (
		_w4459_,
		_w7004_,
		_w7127_,
		_w7128_,
		_w9682_
	);
	LUT4 #(
		.INIT('h04c8)
	) name9649 (
		_w2622_,
		_w4700_,
		_w6978_,
		_w6980_,
		_w9683_
	);
	LUT3 #(
		.INIT('h84)
	) name9650 (
		_w2872_,
		_w4458_,
		_w6975_,
		_w9684_
	);
	LUT3 #(
		.INIT('h07)
	) name9651 (
		_w4684_,
		_w7002_,
		_w9684_,
		_w9685_
	);
	LUT2 #(
		.INIT('h4)
	) name9652 (
		_w9683_,
		_w9685_,
		_w9686_
	);
	LUT3 #(
		.INIT('h9a)
	) name9653 (
		\a[11] ,
		_w9682_,
		_w9686_,
		_w9687_
	);
	LUT3 #(
		.INIT('h54)
	) name9654 (
		_w9680_,
		_w9681_,
		_w9687_,
		_w9688_
	);
	LUT3 #(
		.INIT('h82)
	) name9655 (
		_w4876_,
		_w7135_,
		_w7172_,
		_w9689_
	);
	LUT3 #(
		.INIT('h28)
	) name9656 (
		_w5286_,
		_w7136_,
		_w7168_,
		_w9690_
	);
	LUT2 #(
		.INIT('h8)
	) name9657 (
		_w4875_,
		_w6996_,
		_w9691_
	);
	LUT4 #(
		.INIT('h04c8)
	) name9658 (
		_w2411_,
		_w5271_,
		_w6983_,
		_w6993_,
		_w9692_
	);
	LUT2 #(
		.INIT('h1)
	) name9659 (
		_w9691_,
		_w9692_,
		_w9693_
	);
	LUT2 #(
		.INIT('h4)
	) name9660 (
		_w9690_,
		_w9693_,
		_w9694_
	);
	LUT3 #(
		.INIT('h9a)
	) name9661 (
		\a[8] ,
		_w9689_,
		_w9694_,
		_w9695_
	);
	LUT4 #(
		.INIT('h0445)
	) name9662 (
		_w9451_,
		_w9452_,
		_w9688_,
		_w9695_,
		_w9696_
	);
	LUT4 #(
		.INIT('h9669)
	) name9663 (
		_w9007_,
		_w9199_,
		_w9218_,
		_w9435_,
		_w9697_
	);
	LUT4 #(
		.INIT('ha220)
	) name9664 (
		_w9451_,
		_w9452_,
		_w9688_,
		_w9695_,
		_w9698_
	);
	LUT4 #(
		.INIT('h599a)
	) name9665 (
		_w9451_,
		_w9452_,
		_w9688_,
		_w9695_,
		_w9699_
	);
	LUT3 #(
		.INIT('h51)
	) name9666 (
		_w9696_,
		_w9697_,
		_w9698_,
		_w9700_
	);
	LUT4 #(
		.INIT('h9669)
	) name9667 (
		_w9200_,
		_w9201_,
		_w9207_,
		_w9436_,
		_w9701_
	);
	LUT3 #(
		.INIT('h21)
	) name9668 (
		_w9443_,
		_w9700_,
		_w9701_,
		_w9702_
	);
	LUT2 #(
		.INIT('h6)
	) name9669 (
		_w9697_,
		_w9699_,
		_w9703_
	);
	LUT4 #(
		.INIT('h028a)
	) name9670 (
		_w5523_,
		_w7136_,
		_w7166_,
		_w7167_,
		_w9704_
	);
	LUT3 #(
		.INIT('h0b)
	) name9671 (
		_w7136_,
		_w7166_,
		_w7866_,
		_w9705_
	);
	LUT2 #(
		.INIT('h1)
	) name9672 (
		_w9704_,
		_w9705_,
		_w9706_
	);
	LUT4 #(
		.INIT('h5700)
	) name9673 (
		_w35_,
		_w7418_,
		_w7419_,
		_w9706_,
		_w9707_
	);
	LUT2 #(
		.INIT('h6)
	) name9674 (
		\a[5] ,
		_w9707_,
		_w9708_
	);
	LUT4 #(
		.INIT('h9669)
	) name9675 (
		_w9220_,
		_w9420_,
		_w9426_,
		_w9679_,
		_w9709_
	);
	LUT3 #(
		.INIT('h1e)
	) name9676 (
		_w9467_,
		_w9671_,
		_w9672_,
		_w9710_
	);
	LUT3 #(
		.INIT('h82)
	) name9677 (
		_w4034_,
		_w7117_,
		_w7119_,
		_w9711_
	);
	LUT3 #(
		.INIT('h82)
	) name9678 (
		_w4382_,
		_w6967_,
		_w6969_,
		_w9712_
	);
	LUT2 #(
		.INIT('h8)
	) name9679 (
		_w4033_,
		_w7014_,
		_w9713_
	);
	LUT4 #(
		.INIT('h04c8)
	) name9680 (
		_w3257_,
		_w4367_,
		_w6964_,
		_w6966_,
		_w9714_
	);
	LUT2 #(
		.INIT('h1)
	) name9681 (
		_w9713_,
		_w9714_,
		_w9715_
	);
	LUT2 #(
		.INIT('h4)
	) name9682 (
		_w9712_,
		_w9715_,
		_w9716_
	);
	LUT4 #(
		.INIT('h4844)
	) name9683 (
		\a[14] ,
		_w9710_,
		_w9711_,
		_w9716_,
		_w9717_
	);
	LUT4 #(
		.INIT('h54ab)
	) name9684 (
		_w9473_,
		_w9667_,
		_w9668_,
		_w9670_,
		_w9718_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9685 (
		_w4034_,
		_w7016_,
		_w7115_,
		_w7116_,
		_w9719_
	);
	LUT4 #(
		.INIT('h04c8)
	) name9686 (
		_w3257_,
		_w4382_,
		_w6964_,
		_w6966_,
		_w9720_
	);
	LUT3 #(
		.INIT('h82)
	) name9687 (
		_w4033_,
		_w6960_,
		_w6962_,
		_w9721_
	);
	LUT3 #(
		.INIT('h07)
	) name9688 (
		_w4367_,
		_w7014_,
		_w9721_,
		_w9722_
	);
	LUT2 #(
		.INIT('h4)
	) name9689 (
		_w9720_,
		_w9722_,
		_w9723_
	);
	LUT4 #(
		.INIT('h4844)
	) name9690 (
		\a[14] ,
		_w9718_,
		_w9719_,
		_w9723_,
		_w9724_
	);
	LUT2 #(
		.INIT('h9)
	) name9691 (
		_w9667_,
		_w9669_,
		_w9725_
	);
	LUT4 #(
		.INIT('h5060)
	) name9692 (
		_w3409_,
		_w3650_,
		_w4033_,
		_w6959_,
		_w9726_
	);
	LUT4 #(
		.INIT('h007d)
	) name9693 (
		_w4367_,
		_w6960_,
		_w6962_,
		_w9726_,
		_w9727_
	);
	LUT3 #(
		.INIT('h70)
	) name9694 (
		_w4382_,
		_w7014_,
		_w9727_,
		_w9728_
	);
	LUT4 #(
		.INIT('h95aa)
	) name9695 (
		\a[14] ,
		_w4034_,
		_w7291_,
		_w9728_,
		_w9729_
	);
	LUT2 #(
		.INIT('h2)
	) name9696 (
		_w9725_,
		_w9729_,
		_w9730_
	);
	LUT3 #(
		.INIT('h1e)
	) name9697 (
		_w9488_,
		_w9665_,
		_w9666_,
		_w9731_
	);
	LUT3 #(
		.INIT('h82)
	) name9698 (
		_w4034_,
		_w7111_,
		_w7113_,
		_w9732_
	);
	LUT3 #(
		.INIT('h82)
	) name9699 (
		_w4382_,
		_w6960_,
		_w6962_,
		_w9733_
	);
	LUT2 #(
		.INIT('h8)
	) name9700 (
		_w4033_,
		_w7020_,
		_w9734_
	);
	LUT4 #(
		.INIT('h5060)
	) name9701 (
		_w3409_,
		_w3650_,
		_w4367_,
		_w6959_,
		_w9735_
	);
	LUT2 #(
		.INIT('h1)
	) name9702 (
		_w9734_,
		_w9735_,
		_w9736_
	);
	LUT2 #(
		.INIT('h4)
	) name9703 (
		_w9733_,
		_w9736_,
		_w9737_
	);
	LUT4 #(
		.INIT('h4844)
	) name9704 (
		\a[14] ,
		_w9731_,
		_w9732_,
		_w9737_,
		_w9738_
	);
	LUT4 #(
		.INIT('h54ab)
	) name9705 (
		_w9494_,
		_w9661_,
		_w9662_,
		_w9664_,
		_w9739_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9706 (
		_w4034_,
		_w7022_,
		_w7109_,
		_w7110_,
		_w9740_
	);
	LUT4 #(
		.INIT('h5060)
	) name9707 (
		_w3409_,
		_w3650_,
		_w4382_,
		_w6959_,
		_w9741_
	);
	LUT3 #(
		.INIT('h84)
	) name9708 (
		_w3706_,
		_w4033_,
		_w6957_,
		_w9742_
	);
	LUT3 #(
		.INIT('h07)
	) name9709 (
		_w4367_,
		_w7020_,
		_w9742_,
		_w9743_
	);
	LUT2 #(
		.INIT('h4)
	) name9710 (
		_w9741_,
		_w9743_,
		_w9744_
	);
	LUT4 #(
		.INIT('h4844)
	) name9711 (
		\a[14] ,
		_w9739_,
		_w9740_,
		_w9744_,
		_w9745_
	);
	LUT2 #(
		.INIT('h9)
	) name9712 (
		_w9661_,
		_w9663_,
		_w9746_
	);
	LUT4 #(
		.INIT('h04c8)
	) name9713 (
		_w3882_,
		_w4033_,
		_w6954_,
		_w6956_,
		_w9747_
	);
	LUT4 #(
		.INIT('h007b)
	) name9714 (
		_w3706_,
		_w4367_,
		_w6957_,
		_w9747_,
		_w9748_
	);
	LUT3 #(
		.INIT('h70)
	) name9715 (
		_w4382_,
		_w7020_,
		_w9748_,
		_w9749_
	);
	LUT4 #(
		.INIT('h95aa)
	) name9716 (
		\a[14] ,
		_w4034_,
		_w7465_,
		_w9749_,
		_w9750_
	);
	LUT2 #(
		.INIT('h2)
	) name9717 (
		_w9746_,
		_w9750_,
		_w9751_
	);
	LUT3 #(
		.INIT('h1e)
	) name9718 (
		_w9509_,
		_w9659_,
		_w9660_,
		_w9752_
	);
	LUT3 #(
		.INIT('h82)
	) name9719 (
		_w4034_,
		_w7105_,
		_w7107_,
		_w9753_
	);
	LUT3 #(
		.INIT('h84)
	) name9720 (
		_w3706_,
		_w4382_,
		_w6957_,
		_w9754_
	);
	LUT2 #(
		.INIT('h8)
	) name9721 (
		_w4033_,
		_w7026_,
		_w9755_
	);
	LUT4 #(
		.INIT('h04c8)
	) name9722 (
		_w3882_,
		_w4367_,
		_w6954_,
		_w6956_,
		_w9756_
	);
	LUT2 #(
		.INIT('h1)
	) name9723 (
		_w9755_,
		_w9756_,
		_w9757_
	);
	LUT2 #(
		.INIT('h4)
	) name9724 (
		_w9754_,
		_w9757_,
		_w9758_
	);
	LUT4 #(
		.INIT('h4844)
	) name9725 (
		\a[14] ,
		_w9752_,
		_w9753_,
		_w9758_,
		_w9759_
	);
	LUT4 #(
		.INIT('h54ab)
	) name9726 (
		_w9515_,
		_w9655_,
		_w9656_,
		_w9658_,
		_w9760_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9727 (
		_w4034_,
		_w7028_,
		_w7103_,
		_w7104_,
		_w9761_
	);
	LUT4 #(
		.INIT('h04c8)
	) name9728 (
		_w3882_,
		_w4382_,
		_w6954_,
		_w6956_,
		_w9762_
	);
	LUT3 #(
		.INIT('h84)
	) name9729 (
		_w4030_,
		_w4033_,
		_w6952_,
		_w9763_
	);
	LUT3 #(
		.INIT('h07)
	) name9730 (
		_w4367_,
		_w7026_,
		_w9763_,
		_w9764_
	);
	LUT2 #(
		.INIT('h4)
	) name9731 (
		_w9762_,
		_w9764_,
		_w9765_
	);
	LUT4 #(
		.INIT('h4844)
	) name9732 (
		\a[14] ,
		_w9760_,
		_w9761_,
		_w9765_,
		_w9766_
	);
	LUT2 #(
		.INIT('h9)
	) name9733 (
		_w9655_,
		_w9657_,
		_w9767_
	);
	LUT4 #(
		.INIT('h2228)
	) name9734 (
		_w4033_,
		_w4099_,
		_w4378_,
		_w6951_,
		_w9768_
	);
	LUT4 #(
		.INIT('h007b)
	) name9735 (
		_w4030_,
		_w4367_,
		_w6952_,
		_w9768_,
		_w9769_
	);
	LUT3 #(
		.INIT('h70)
	) name9736 (
		_w4382_,
		_w7026_,
		_w9769_,
		_w9770_
	);
	LUT4 #(
		.INIT('h95aa)
	) name9737 (
		\a[14] ,
		_w4034_,
		_w7562_,
		_w9770_,
		_w9771_
	);
	LUT2 #(
		.INIT('h2)
	) name9738 (
		_w9767_,
		_w9771_,
		_w9772_
	);
	LUT3 #(
		.INIT('h1e)
	) name9739 (
		_w9530_,
		_w9653_,
		_w9654_,
		_w9773_
	);
	LUT3 #(
		.INIT('h82)
	) name9740 (
		_w4034_,
		_w7099_,
		_w7101_,
		_w9774_
	);
	LUT3 #(
		.INIT('h84)
	) name9741 (
		_w4030_,
		_w4382_,
		_w6952_,
		_w9775_
	);
	LUT2 #(
		.INIT('h8)
	) name9742 (
		_w4033_,
		_w7032_,
		_w9776_
	);
	LUT4 #(
		.INIT('h4448)
	) name9743 (
		_w4099_,
		_w4367_,
		_w4378_,
		_w6951_,
		_w9777_
	);
	LUT2 #(
		.INIT('h1)
	) name9744 (
		_w9776_,
		_w9777_,
		_w9778_
	);
	LUT2 #(
		.INIT('h4)
	) name9745 (
		_w9775_,
		_w9778_,
		_w9779_
	);
	LUT4 #(
		.INIT('h4844)
	) name9746 (
		\a[14] ,
		_w9773_,
		_w9774_,
		_w9779_,
		_w9780_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9747 (
		_w4034_,
		_w7034_,
		_w7097_,
		_w7098_,
		_w9781_
	);
	LUT4 #(
		.INIT('h5060)
	) name9748 (
		_w4099_,
		_w4378_,
		_w4382_,
		_w6951_,
		_w9782_
	);
	LUT3 #(
		.INIT('h82)
	) name9749 (
		_w4033_,
		_w6947_,
		_w6949_,
		_w9783_
	);
	LUT3 #(
		.INIT('h07)
	) name9750 (
		_w4367_,
		_w7032_,
		_w9783_,
		_w9784_
	);
	LUT2 #(
		.INIT('h4)
	) name9751 (
		_w9782_,
		_w9784_,
		_w9785_
	);
	LUT4 #(
		.INIT('h54ab)
	) name9752 (
		_w9536_,
		_w9649_,
		_w9650_,
		_w9652_,
		_w9786_
	);
	LUT4 #(
		.INIT('h6500)
	) name9753 (
		\a[14] ,
		_w9781_,
		_w9785_,
		_w9786_,
		_w9787_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9754 (
		_w4033_,
		_w4695_,
		_w6944_,
		_w6946_,
		_w9788_
	);
	LUT4 #(
		.INIT('h007d)
	) name9755 (
		_w4367_,
		_w6947_,
		_w6949_,
		_w9788_,
		_w9789_
	);
	LUT3 #(
		.INIT('h70)
	) name9756 (
		_w4382_,
		_w7032_,
		_w9789_,
		_w9790_
	);
	LUT4 #(
		.INIT('h95aa)
	) name9757 (
		\a[14] ,
		_w4034_,
		_w7882_,
		_w9790_,
		_w9791_
	);
	LUT2 #(
		.INIT('h9)
	) name9758 (
		_w9649_,
		_w9651_,
		_w9792_
	);
	LUT2 #(
		.INIT('h4)
	) name9759 (
		_w9791_,
		_w9792_,
		_w9793_
	);
	LUT3 #(
		.INIT('h1e)
	) name9760 (
		_w9551_,
		_w9647_,
		_w9648_,
		_w9794_
	);
	LUT3 #(
		.INIT('h82)
	) name9761 (
		_w4034_,
		_w7093_,
		_w7095_,
		_w9795_
	);
	LUT3 #(
		.INIT('h82)
	) name9762 (
		_w4382_,
		_w6947_,
		_w6949_,
		_w9796_
	);
	LUT2 #(
		.INIT('h8)
	) name9763 (
		_w4033_,
		_w7038_,
		_w9797_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9764 (
		_w4367_,
		_w4695_,
		_w6944_,
		_w6946_,
		_w9798_
	);
	LUT2 #(
		.INIT('h1)
	) name9765 (
		_w9797_,
		_w9798_,
		_w9799_
	);
	LUT2 #(
		.INIT('h4)
	) name9766 (
		_w9796_,
		_w9799_,
		_w9800_
	);
	LUT4 #(
		.INIT('h4844)
	) name9767 (
		\a[14] ,
		_w9794_,
		_w9795_,
		_w9800_,
		_w9801_
	);
	LUT4 #(
		.INIT('h54ab)
	) name9768 (
		_w9557_,
		_w9643_,
		_w9644_,
		_w9646_,
		_w9802_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9769 (
		_w4034_,
		_w7040_,
		_w7091_,
		_w7092_,
		_w9803_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9770 (
		_w4382_,
		_w4695_,
		_w6944_,
		_w6946_,
		_w9804_
	);
	LUT3 #(
		.INIT('h82)
	) name9771 (
		_w4033_,
		_w6940_,
		_w6942_,
		_w9805_
	);
	LUT3 #(
		.INIT('h07)
	) name9772 (
		_w4367_,
		_w7038_,
		_w9805_,
		_w9806_
	);
	LUT2 #(
		.INIT('h4)
	) name9773 (
		_w9804_,
		_w9806_,
		_w9807_
	);
	LUT4 #(
		.INIT('h4844)
	) name9774 (
		\a[14] ,
		_w9802_,
		_w9803_,
		_w9807_,
		_w9808_
	);
	LUT2 #(
		.INIT('h9)
	) name9775 (
		_w9643_,
		_w9645_,
		_w9809_
	);
	LUT4 #(
		.INIT('h2228)
	) name9776 (
		_w4033_,
		_w5067_,
		_w5282_,
		_w6939_,
		_w9810_
	);
	LUT4 #(
		.INIT('h007d)
	) name9777 (
		_w4367_,
		_w6940_,
		_w6942_,
		_w9810_,
		_w9811_
	);
	LUT3 #(
		.INIT('h70)
	) name9778 (
		_w4382_,
		_w7038_,
		_w9811_,
		_w9812_
	);
	LUT4 #(
		.INIT('h95aa)
	) name9779 (
		\a[14] ,
		_w4034_,
		_w8018_,
		_w9812_,
		_w9813_
	);
	LUT2 #(
		.INIT('h2)
	) name9780 (
		_w9809_,
		_w9813_,
		_w9814_
	);
	LUT3 #(
		.INIT('h82)
	) name9781 (
		_w4034_,
		_w7087_,
		_w7089_,
		_w9815_
	);
	LUT3 #(
		.INIT('h82)
	) name9782 (
		_w4382_,
		_w6940_,
		_w6942_,
		_w9816_
	);
	LUT2 #(
		.INIT('h8)
	) name9783 (
		_w4033_,
		_w7044_,
		_w9817_
	);
	LUT4 #(
		.INIT('h2228)
	) name9784 (
		_w4367_,
		_w5067_,
		_w5282_,
		_w6939_,
		_w9818_
	);
	LUT2 #(
		.INIT('h1)
	) name9785 (
		_w9817_,
		_w9818_,
		_w9819_
	);
	LUT2 #(
		.INIT('h4)
	) name9786 (
		_w9816_,
		_w9819_,
		_w9820_
	);
	LUT3 #(
		.INIT('h1e)
	) name9787 (
		_w9572_,
		_w9641_,
		_w9642_,
		_w9821_
	);
	LUT4 #(
		.INIT('h6500)
	) name9788 (
		\a[14] ,
		_w9815_,
		_w9820_,
		_w9821_,
		_w9822_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9789 (
		_w4034_,
		_w7046_,
		_w7085_,
		_w7086_,
		_w9823_
	);
	LUT4 #(
		.INIT('h2228)
	) name9790 (
		_w4382_,
		_w5067_,
		_w5282_,
		_w6939_,
		_w9824_
	);
	LUT3 #(
		.INIT('h82)
	) name9791 (
		_w4033_,
		_w6935_,
		_w6937_,
		_w9825_
	);
	LUT3 #(
		.INIT('h07)
	) name9792 (
		_w4367_,
		_w7044_,
		_w9825_,
		_w9826_
	);
	LUT2 #(
		.INIT('h4)
	) name9793 (
		_w9824_,
		_w9826_,
		_w9827_
	);
	LUT4 #(
		.INIT('h54ab)
	) name9794 (
		_w9578_,
		_w9637_,
		_w9638_,
		_w9640_,
		_w9828_
	);
	LUT4 #(
		.INIT('h6500)
	) name9795 (
		\a[14] ,
		_w9823_,
		_w9827_,
		_w9828_,
		_w9829_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9796 (
		_w4033_,
		_w6043_,
		_w6933_,
		_w6934_,
		_w9830_
	);
	LUT4 #(
		.INIT('h007d)
	) name9797 (
		_w4367_,
		_w6935_,
		_w6937_,
		_w9830_,
		_w9831_
	);
	LUT3 #(
		.INIT('h70)
	) name9798 (
		_w4382_,
		_w7044_,
		_w9831_,
		_w9832_
	);
	LUT4 #(
		.INIT('h95aa)
	) name9799 (
		\a[14] ,
		_w4034_,
		_w8005_,
		_w9832_,
		_w9833_
	);
	LUT2 #(
		.INIT('h9)
	) name9800 (
		_w9637_,
		_w9639_,
		_w9834_
	);
	LUT2 #(
		.INIT('h4)
	) name9801 (
		_w9833_,
		_w9834_,
		_w9835_
	);
	LUT3 #(
		.INIT('h1e)
	) name9802 (
		_w9593_,
		_w9635_,
		_w9636_,
		_w9836_
	);
	LUT3 #(
		.INIT('h82)
	) name9803 (
		_w4034_,
		_w7081_,
		_w7083_,
		_w9837_
	);
	LUT3 #(
		.INIT('h82)
	) name9804 (
		_w4382_,
		_w6935_,
		_w6937_,
		_w9838_
	);
	LUT2 #(
		.INIT('h8)
	) name9805 (
		_w4033_,
		_w7050_,
		_w9839_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9806 (
		_w4367_,
		_w6043_,
		_w6933_,
		_w6934_,
		_w9840_
	);
	LUT2 #(
		.INIT('h1)
	) name9807 (
		_w9839_,
		_w9840_,
		_w9841_
	);
	LUT2 #(
		.INIT('h4)
	) name9808 (
		_w9838_,
		_w9841_,
		_w9842_
	);
	LUT4 #(
		.INIT('h4844)
	) name9809 (
		\a[14] ,
		_w9836_,
		_w9837_,
		_w9842_,
		_w9843_
	);
	LUT4 #(
		.INIT('h54ab)
	) name9810 (
		_w9600_,
		_w9631_,
		_w9632_,
		_w9634_,
		_w9844_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9811 (
		_w4034_,
		_w7052_,
		_w7079_,
		_w7080_,
		_w9845_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9812 (
		_w4382_,
		_w6043_,
		_w6933_,
		_w6934_,
		_w9846_
	);
	LUT3 #(
		.INIT('h82)
	) name9813 (
		_w4033_,
		_w6929_,
		_w6931_,
		_w9847_
	);
	LUT3 #(
		.INIT('h07)
	) name9814 (
		_w4367_,
		_w7050_,
		_w9847_,
		_w9848_
	);
	LUT2 #(
		.INIT('h4)
	) name9815 (
		_w9846_,
		_w9848_,
		_w9849_
	);
	LUT4 #(
		.INIT('h4844)
	) name9816 (
		\a[14] ,
		_w9844_,
		_w9845_,
		_w9849_,
		_w9850_
	);
	LUT2 #(
		.INIT('h9)
	) name9817 (
		_w9631_,
		_w9633_,
		_w9851_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9818 (
		_w4033_,
		_w6645_,
		_w6926_,
		_w6928_,
		_w9852_
	);
	LUT4 #(
		.INIT('h007d)
	) name9819 (
		_w4367_,
		_w6929_,
		_w6931_,
		_w9852_,
		_w9853_
	);
	LUT3 #(
		.INIT('h70)
	) name9820 (
		_w4382_,
		_w7050_,
		_w9853_,
		_w9854_
	);
	LUT4 #(
		.INIT('h95aa)
	) name9821 (
		\a[14] ,
		_w4034_,
		_w8227_,
		_w9854_,
		_w9855_
	);
	LUT2 #(
		.INIT('h2)
	) name9822 (
		_w9851_,
		_w9855_,
		_w9856_
	);
	LUT3 #(
		.INIT('h82)
	) name9823 (
		_w4034_,
		_w7075_,
		_w7077_,
		_w9857_
	);
	LUT3 #(
		.INIT('h82)
	) name9824 (
		_w4382_,
		_w6929_,
		_w6931_,
		_w9858_
	);
	LUT2 #(
		.INIT('h8)
	) name9825 (
		_w4033_,
		_w7056_,
		_w9859_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9826 (
		_w4367_,
		_w6645_,
		_w6926_,
		_w6928_,
		_w9860_
	);
	LUT2 #(
		.INIT('h1)
	) name9827 (
		_w9859_,
		_w9860_,
		_w9861_
	);
	LUT2 #(
		.INIT('h4)
	) name9828 (
		_w9858_,
		_w9861_,
		_w9862_
	);
	LUT2 #(
		.INIT('h9)
	) name9829 (
		_w9628_,
		_w9630_,
		_w9863_
	);
	LUT4 #(
		.INIT('h6500)
	) name9830 (
		\a[14] ,
		_w9857_,
		_w9862_,
		_w9863_,
		_w9864_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9831 (
		_w4034_,
		_w7058_,
		_w7073_,
		_w7074_,
		_w9865_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9832 (
		_w4382_,
		_w6645_,
		_w6926_,
		_w6928_,
		_w9866_
	);
	LUT3 #(
		.INIT('h82)
	) name9833 (
		_w4033_,
		_w6922_,
		_w6924_,
		_w9867_
	);
	LUT3 #(
		.INIT('h07)
	) name9834 (
		_w4367_,
		_w7056_,
		_w9867_,
		_w9868_
	);
	LUT2 #(
		.INIT('h4)
	) name9835 (
		_w9866_,
		_w9868_,
		_w9869_
	);
	LUT4 #(
		.INIT('h9a65)
	) name9836 (
		\a[17] ,
		_w9621_,
		_w9625_,
		_w9626_,
		_w9870_
	);
	LUT4 #(
		.INIT('h6500)
	) name9837 (
		\a[14] ,
		_w9865_,
		_w9869_,
		_w9870_,
		_w9871_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9838 (
		_w4033_,
		_w6669_,
		_w6919_,
		_w6921_,
		_w9872_
	);
	LUT4 #(
		.INIT('h007d)
	) name9839 (
		_w4367_,
		_w6922_,
		_w6924_,
		_w9872_,
		_w9873_
	);
	LUT3 #(
		.INIT('h70)
	) name9840 (
		_w4382_,
		_w7056_,
		_w9873_,
		_w9874_
	);
	LUT4 #(
		.INIT('h95aa)
	) name9841 (
		\a[14] ,
		_w4034_,
		_w8298_,
		_w9874_,
		_w9875_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name9842 (
		\a[17] ,
		_w9613_,
		_w9610_,
		_w9612_,
		_w9876_
	);
	LUT3 #(
		.INIT('h4b)
	) name9843 (
		_w9616_,
		_w9619_,
		_w9876_,
		_w9877_
	);
	LUT2 #(
		.INIT('h4)
	) name9844 (
		_w9875_,
		_w9877_,
		_w9878_
	);
	LUT3 #(
		.INIT('h82)
	) name9845 (
		_w4034_,
		_w7069_,
		_w7071_,
		_w9879_
	);
	LUT3 #(
		.INIT('h82)
	) name9846 (
		_w4382_,
		_w6922_,
		_w6924_,
		_w9880_
	);
	LUT2 #(
		.INIT('h8)
	) name9847 (
		_w4033_,
		_w7062_,
		_w9881_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9848 (
		_w4367_,
		_w6669_,
		_w6919_,
		_w6921_,
		_w9882_
	);
	LUT2 #(
		.INIT('h1)
	) name9849 (
		_w9881_,
		_w9882_,
		_w9883_
	);
	LUT2 #(
		.INIT('h4)
	) name9850 (
		_w9880_,
		_w9883_,
		_w9884_
	);
	LUT2 #(
		.INIT('h8)
	) name9851 (
		\a[17] ,
		_w9613_,
		_w9885_
	);
	LUT3 #(
		.INIT('h4b)
	) name9852 (
		_w9610_,
		_w9612_,
		_w9885_,
		_w9886_
	);
	LUT4 #(
		.INIT('h6500)
	) name9853 (
		\a[14] ,
		_w9879_,
		_w9884_,
		_w9886_,
		_w9887_
	);
	LUT4 #(
		.INIT('h2882)
	) name9854 (
		_w4034_,
		_w6914_,
		_w6916_,
		_w7067_,
		_w9888_
	);
	LUT4 #(
		.INIT('ha802)
	) name9855 (
		_w4367_,
		_w6689_,
		_w6911_,
		_w6913_,
		_w9889_
	);
	LUT4 #(
		.INIT('h007d)
	) name9856 (
		_w4382_,
		_w6914_,
		_w6916_,
		_w9889_,
		_w9890_
	);
	LUT4 #(
		.INIT('h5401)
	) name9857 (
		_w4032_,
		_w6689_,
		_w6911_,
		_w6913_,
		_w9891_
	);
	LUT2 #(
		.INIT('h2)
	) name9858 (
		\a[14] ,
		_w9891_,
		_w9892_
	);
	LUT3 #(
		.INIT('h40)
	) name9859 (
		_w9888_,
		_w9890_,
		_w9892_,
		_w9893_
	);
	LUT3 #(
		.INIT('h28)
	) name9860 (
		_w4034_,
		_w7062_,
		_w8358_,
		_w9894_
	);
	LUT4 #(
		.INIT('ha802)
	) name9861 (
		_w4033_,
		_w6689_,
		_w6911_,
		_w6913_,
		_w9895_
	);
	LUT4 #(
		.INIT('h007d)
	) name9862 (
		_w4367_,
		_w6914_,
		_w6916_,
		_w9895_,
		_w9896_
	);
	LUT3 #(
		.INIT('h70)
	) name9863 (
		_w4382_,
		_w7062_,
		_w9896_,
		_w9897_
	);
	LUT4 #(
		.INIT('h0800)
	) name9864 (
		_w9613_,
		_w9893_,
		_w9894_,
		_w9897_,
		_w9898_
	);
	LUT3 #(
		.INIT('h28)
	) name9865 (
		_w4034_,
		_w7065_,
		_w7068_,
		_w9899_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9866 (
		_w4382_,
		_w6669_,
		_w6919_,
		_w6921_,
		_w9900_
	);
	LUT3 #(
		.INIT('h82)
	) name9867 (
		_w4033_,
		_w6914_,
		_w6916_,
		_w9901_
	);
	LUT3 #(
		.INIT('h07)
	) name9868 (
		_w4367_,
		_w7062_,
		_w9901_,
		_w9902_
	);
	LUT2 #(
		.INIT('h4)
	) name9869 (
		_w9900_,
		_w9902_,
		_w9903_
	);
	LUT4 #(
		.INIT('ha6aa)
	) name9870 (
		_w9613_,
		_w9893_,
		_w9894_,
		_w9897_,
		_w9904_
	);
	LUT4 #(
		.INIT('h6500)
	) name9871 (
		\a[14] ,
		_w9899_,
		_w9903_,
		_w9904_,
		_w9905_
	);
	LUT2 #(
		.INIT('h1)
	) name9872 (
		_w9898_,
		_w9905_,
		_w9906_
	);
	LUT4 #(
		.INIT('h009a)
	) name9873 (
		\a[14] ,
		_w9879_,
		_w9884_,
		_w9886_,
		_w9907_
	);
	LUT4 #(
		.INIT('h9a65)
	) name9874 (
		\a[14] ,
		_w9879_,
		_w9884_,
		_w9886_,
		_w9908_
	);
	LUT3 #(
		.INIT('h54)
	) name9875 (
		_w9887_,
		_w9906_,
		_w9907_,
		_w9909_
	);
	LUT2 #(
		.INIT('h2)
	) name9876 (
		_w9875_,
		_w9877_,
		_w9910_
	);
	LUT2 #(
		.INIT('h9)
	) name9877 (
		_w9875_,
		_w9877_,
		_w9911_
	);
	LUT4 #(
		.INIT('h9a65)
	) name9878 (
		\a[14] ,
		_w9865_,
		_w9869_,
		_w9870_,
		_w9912_
	);
	LUT4 #(
		.INIT('h4d00)
	) name9879 (
		_w9875_,
		_w9877_,
		_w9909_,
		_w9912_,
		_w9913_
	);
	LUT4 #(
		.INIT('h9a65)
	) name9880 (
		\a[14] ,
		_w9857_,
		_w9862_,
		_w9863_,
		_w9914_
	);
	LUT4 #(
		.INIT('h0155)
	) name9881 (
		_w9864_,
		_w9871_,
		_w9913_,
		_w9914_,
		_w9915_
	);
	LUT2 #(
		.INIT('h4)
	) name9882 (
		_w9851_,
		_w9855_,
		_w9916_
	);
	LUT2 #(
		.INIT('h9)
	) name9883 (
		_w9851_,
		_w9855_,
		_w9917_
	);
	LUT4 #(
		.INIT('h9699)
	) name9884 (
		\a[14] ,
		_w9844_,
		_w9845_,
		_w9849_,
		_w9918_
	);
	LUT4 #(
		.INIT('h2b00)
	) name9885 (
		_w9851_,
		_w9855_,
		_w9915_,
		_w9918_,
		_w9919_
	);
	LUT4 #(
		.INIT('h9699)
	) name9886 (
		\a[14] ,
		_w9836_,
		_w9837_,
		_w9842_,
		_w9920_
	);
	LUT4 #(
		.INIT('h0155)
	) name9887 (
		_w9843_,
		_w9850_,
		_w9919_,
		_w9920_,
		_w9921_
	);
	LUT2 #(
		.INIT('h2)
	) name9888 (
		_w9833_,
		_w9834_,
		_w9922_
	);
	LUT2 #(
		.INIT('h9)
	) name9889 (
		_w9833_,
		_w9834_,
		_w9923_
	);
	LUT4 #(
		.INIT('h9a65)
	) name9890 (
		\a[14] ,
		_w9823_,
		_w9827_,
		_w9828_,
		_w9924_
	);
	LUT4 #(
		.INIT('h4d00)
	) name9891 (
		_w9833_,
		_w9834_,
		_w9921_,
		_w9924_,
		_w9925_
	);
	LUT4 #(
		.INIT('h9a65)
	) name9892 (
		\a[14] ,
		_w9815_,
		_w9820_,
		_w9821_,
		_w9926_
	);
	LUT4 #(
		.INIT('h0155)
	) name9893 (
		_w9822_,
		_w9829_,
		_w9925_,
		_w9926_,
		_w9927_
	);
	LUT2 #(
		.INIT('h4)
	) name9894 (
		_w9809_,
		_w9813_,
		_w9928_
	);
	LUT2 #(
		.INIT('h9)
	) name9895 (
		_w9809_,
		_w9813_,
		_w9929_
	);
	LUT4 #(
		.INIT('h9699)
	) name9896 (
		\a[14] ,
		_w9802_,
		_w9803_,
		_w9807_,
		_w9930_
	);
	LUT4 #(
		.INIT('h2b00)
	) name9897 (
		_w9809_,
		_w9813_,
		_w9927_,
		_w9930_,
		_w9931_
	);
	LUT4 #(
		.INIT('h9699)
	) name9898 (
		\a[14] ,
		_w9794_,
		_w9795_,
		_w9800_,
		_w9932_
	);
	LUT4 #(
		.INIT('h0155)
	) name9899 (
		_w9801_,
		_w9808_,
		_w9931_,
		_w9932_,
		_w9933_
	);
	LUT2 #(
		.INIT('h2)
	) name9900 (
		_w9791_,
		_w9792_,
		_w9934_
	);
	LUT2 #(
		.INIT('h9)
	) name9901 (
		_w9791_,
		_w9792_,
		_w9935_
	);
	LUT4 #(
		.INIT('h9a65)
	) name9902 (
		\a[14] ,
		_w9781_,
		_w9785_,
		_w9786_,
		_w9936_
	);
	LUT4 #(
		.INIT('h4d00)
	) name9903 (
		_w9791_,
		_w9792_,
		_w9933_,
		_w9936_,
		_w9937_
	);
	LUT4 #(
		.INIT('h9699)
	) name9904 (
		\a[14] ,
		_w9773_,
		_w9774_,
		_w9779_,
		_w9938_
	);
	LUT4 #(
		.INIT('h0155)
	) name9905 (
		_w9780_,
		_w9787_,
		_w9937_,
		_w9938_,
		_w9939_
	);
	LUT2 #(
		.INIT('h4)
	) name9906 (
		_w9767_,
		_w9771_,
		_w9940_
	);
	LUT2 #(
		.INIT('h9)
	) name9907 (
		_w9767_,
		_w9771_,
		_w9941_
	);
	LUT4 #(
		.INIT('h9699)
	) name9908 (
		\a[14] ,
		_w9760_,
		_w9761_,
		_w9765_,
		_w9942_
	);
	LUT4 #(
		.INIT('h2b00)
	) name9909 (
		_w9767_,
		_w9771_,
		_w9939_,
		_w9942_,
		_w9943_
	);
	LUT4 #(
		.INIT('h9699)
	) name9910 (
		\a[14] ,
		_w9752_,
		_w9753_,
		_w9758_,
		_w9944_
	);
	LUT4 #(
		.INIT('h0155)
	) name9911 (
		_w9759_,
		_w9766_,
		_w9943_,
		_w9944_,
		_w9945_
	);
	LUT2 #(
		.INIT('h4)
	) name9912 (
		_w9746_,
		_w9750_,
		_w9946_
	);
	LUT2 #(
		.INIT('h9)
	) name9913 (
		_w9746_,
		_w9750_,
		_w9947_
	);
	LUT4 #(
		.INIT('h9699)
	) name9914 (
		\a[14] ,
		_w9739_,
		_w9740_,
		_w9744_,
		_w9948_
	);
	LUT4 #(
		.INIT('h2b00)
	) name9915 (
		_w9746_,
		_w9750_,
		_w9945_,
		_w9948_,
		_w9949_
	);
	LUT4 #(
		.INIT('h9699)
	) name9916 (
		\a[14] ,
		_w9731_,
		_w9732_,
		_w9737_,
		_w9950_
	);
	LUT4 #(
		.INIT('h0155)
	) name9917 (
		_w9738_,
		_w9745_,
		_w9949_,
		_w9950_,
		_w9951_
	);
	LUT2 #(
		.INIT('h4)
	) name9918 (
		_w9725_,
		_w9729_,
		_w9952_
	);
	LUT2 #(
		.INIT('h9)
	) name9919 (
		_w9725_,
		_w9729_,
		_w9953_
	);
	LUT4 #(
		.INIT('h9699)
	) name9920 (
		\a[14] ,
		_w9718_,
		_w9719_,
		_w9723_,
		_w9954_
	);
	LUT4 #(
		.INIT('h2b00)
	) name9921 (
		_w9725_,
		_w9729_,
		_w9951_,
		_w9954_,
		_w9955_
	);
	LUT4 #(
		.INIT('h9699)
	) name9922 (
		\a[14] ,
		_w9710_,
		_w9711_,
		_w9716_,
		_w9956_
	);
	LUT4 #(
		.INIT('h0155)
	) name9923 (
		_w9717_,
		_w9724_,
		_w9955_,
		_w9956_,
		_w9957_
	);
	LUT4 #(
		.INIT('h0069)
	) name9924 (
		_w9673_,
		_w9674_,
		_w9678_,
		_w9957_,
		_w9958_
	);
	LUT4 #(
		.INIT('h9600)
	) name9925 (
		_w9673_,
		_w9674_,
		_w9678_,
		_w9957_,
		_w9959_
	);
	LUT4 #(
		.INIT('h04c8)
	) name9926 (
		_w2983_,
		_w4458_,
		_w6972_,
		_w6974_,
		_w9960_
	);
	LUT4 #(
		.INIT('h007b)
	) name9927 (
		_w2872_,
		_w4684_,
		_w6975_,
		_w9960_,
		_w9961_
	);
	LUT3 #(
		.INIT('h70)
	) name9928 (
		_w4700_,
		_w7002_,
		_w9961_,
		_w9962_
	);
	LUT4 #(
		.INIT('h95aa)
	) name9929 (
		\a[11] ,
		_w4459_,
		_w7426_,
		_w9962_,
		_w9963_
	);
	LUT3 #(
		.INIT('h54)
	) name9930 (
		_w9958_,
		_w9959_,
		_w9963_,
		_w9964_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9931 (
		_w4876_,
		_w6998_,
		_w7133_,
		_w7134_,
		_w9965_
	);
	LUT4 #(
		.INIT('h04c8)
	) name9932 (
		_w2411_,
		_w5286_,
		_w6983_,
		_w6993_,
		_w9966_
	);
	LUT3 #(
		.INIT('h84)
	) name9933 (
		_w2546_,
		_w4875_,
		_w6981_,
		_w9967_
	);
	LUT3 #(
		.INIT('h07)
	) name9934 (
		_w5271_,
		_w6996_,
		_w9967_,
		_w9968_
	);
	LUT2 #(
		.INIT('h4)
	) name9935 (
		_w9966_,
		_w9968_,
		_w9969_
	);
	LUT3 #(
		.INIT('h9a)
	) name9936 (
		\a[8] ,
		_w9965_,
		_w9969_,
		_w9970_
	);
	LUT4 #(
		.INIT('hf660)
	) name9937 (
		_w9687_,
		_w9709_,
		_w9964_,
		_w9970_,
		_w9971_
	);
	LUT2 #(
		.INIT('h1)
	) name9938 (
		_w9708_,
		_w9971_,
		_w9972_
	);
	LUT2 #(
		.INIT('h8)
	) name9939 (
		_w9708_,
		_w9971_,
		_w9973_
	);
	LUT3 #(
		.INIT('h96)
	) name9940 (
		_w9452_,
		_w9688_,
		_w9695_,
		_w9974_
	);
	LUT3 #(
		.INIT('h45)
	) name9941 (
		_w9972_,
		_w9973_,
		_w9974_,
		_w9975_
	);
	LUT2 #(
		.INIT('h2)
	) name9942 (
		_w9703_,
		_w9975_,
		_w9976_
	);
	LUT2 #(
		.INIT('h6)
	) name9943 (
		_w9708_,
		_w9971_,
		_w9977_
	);
	LUT4 #(
		.INIT('h9669)
	) name9944 (
		_w9687_,
		_w9709_,
		_w9964_,
		_w9970_,
		_w9978_
	);
	LUT3 #(
		.INIT('h82)
	) name9945 (
		_w4459_,
		_w7123_,
		_w7125_,
		_w9979_
	);
	LUT3 #(
		.INIT('h84)
	) name9946 (
		_w2872_,
		_w4700_,
		_w6975_,
		_w9980_
	);
	LUT2 #(
		.INIT('h8)
	) name9947 (
		_w4458_,
		_w7008_,
		_w9981_
	);
	LUT4 #(
		.INIT('h04c8)
	) name9948 (
		_w2983_,
		_w4684_,
		_w6972_,
		_w6974_,
		_w9982_
	);
	LUT2 #(
		.INIT('h1)
	) name9949 (
		_w9981_,
		_w9982_,
		_w9983_
	);
	LUT2 #(
		.INIT('h4)
	) name9950 (
		_w9980_,
		_w9983_,
		_w9984_
	);
	LUT3 #(
		.INIT('h1e)
	) name9951 (
		_w9724_,
		_w9955_,
		_w9956_,
		_w9985_
	);
	LUT4 #(
		.INIT('h6500)
	) name9952 (
		\a[11] ,
		_w9979_,
		_w9984_,
		_w9985_,
		_w9986_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9953 (
		_w4459_,
		_w7010_,
		_w7121_,
		_w7122_,
		_w9987_
	);
	LUT4 #(
		.INIT('h04c8)
	) name9954 (
		_w2983_,
		_w4700_,
		_w6972_,
		_w6974_,
		_w9988_
	);
	LUT3 #(
		.INIT('h82)
	) name9955 (
		_w4458_,
		_w6967_,
		_w6969_,
		_w9989_
	);
	LUT3 #(
		.INIT('h07)
	) name9956 (
		_w4684_,
		_w7008_,
		_w9989_,
		_w9990_
	);
	LUT2 #(
		.INIT('h4)
	) name9957 (
		_w9988_,
		_w9990_,
		_w9991_
	);
	LUT4 #(
		.INIT('h54ab)
	) name9958 (
		_w9730_,
		_w9951_,
		_w9952_,
		_w9954_,
		_w9992_
	);
	LUT4 #(
		.INIT('h6500)
	) name9959 (
		\a[11] ,
		_w9987_,
		_w9991_,
		_w9992_,
		_w9993_
	);
	LUT4 #(
		.INIT('h04c8)
	) name9960 (
		_w3257_,
		_w4458_,
		_w6964_,
		_w6966_,
		_w9994_
	);
	LUT4 #(
		.INIT('h007d)
	) name9961 (
		_w4684_,
		_w6967_,
		_w6969_,
		_w9994_,
		_w9995_
	);
	LUT3 #(
		.INIT('h70)
	) name9962 (
		_w4700_,
		_w7008_,
		_w9995_,
		_w9996_
	);
	LUT4 #(
		.INIT('h95aa)
	) name9963 (
		\a[11] ,
		_w4459_,
		_w7403_,
		_w9996_,
		_w9997_
	);
	LUT2 #(
		.INIT('h9)
	) name9964 (
		_w9951_,
		_w9953_,
		_w9998_
	);
	LUT2 #(
		.INIT('h4)
	) name9965 (
		_w9997_,
		_w9998_,
		_w9999_
	);
	LUT3 #(
		.INIT('h82)
	) name9966 (
		_w4459_,
		_w7117_,
		_w7119_,
		_w10000_
	);
	LUT3 #(
		.INIT('h82)
	) name9967 (
		_w4700_,
		_w6967_,
		_w6969_,
		_w10001_
	);
	LUT2 #(
		.INIT('h8)
	) name9968 (
		_w4458_,
		_w7014_,
		_w10002_
	);
	LUT4 #(
		.INIT('h04c8)
	) name9969 (
		_w3257_,
		_w4684_,
		_w6964_,
		_w6966_,
		_w10003_
	);
	LUT2 #(
		.INIT('h1)
	) name9970 (
		_w10002_,
		_w10003_,
		_w10004_
	);
	LUT2 #(
		.INIT('h4)
	) name9971 (
		_w10001_,
		_w10004_,
		_w10005_
	);
	LUT3 #(
		.INIT('h1e)
	) name9972 (
		_w9745_,
		_w9949_,
		_w9950_,
		_w10006_
	);
	LUT4 #(
		.INIT('h6500)
	) name9973 (
		\a[11] ,
		_w10000_,
		_w10005_,
		_w10006_,
		_w10007_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9974 (
		_w4459_,
		_w7016_,
		_w7115_,
		_w7116_,
		_w10008_
	);
	LUT4 #(
		.INIT('h04c8)
	) name9975 (
		_w3257_,
		_w4700_,
		_w6964_,
		_w6966_,
		_w10009_
	);
	LUT3 #(
		.INIT('h82)
	) name9976 (
		_w4458_,
		_w6960_,
		_w6962_,
		_w10010_
	);
	LUT3 #(
		.INIT('h07)
	) name9977 (
		_w4684_,
		_w7014_,
		_w10010_,
		_w10011_
	);
	LUT2 #(
		.INIT('h4)
	) name9978 (
		_w10009_,
		_w10011_,
		_w10012_
	);
	LUT4 #(
		.INIT('h54ab)
	) name9979 (
		_w9751_,
		_w9945_,
		_w9946_,
		_w9948_,
		_w10013_
	);
	LUT4 #(
		.INIT('h6500)
	) name9980 (
		\a[11] ,
		_w10008_,
		_w10012_,
		_w10013_,
		_w10014_
	);
	LUT4 #(
		.INIT('h5060)
	) name9981 (
		_w3409_,
		_w3650_,
		_w4458_,
		_w6959_,
		_w10015_
	);
	LUT4 #(
		.INIT('h007d)
	) name9982 (
		_w4684_,
		_w6960_,
		_w6962_,
		_w10015_,
		_w10016_
	);
	LUT3 #(
		.INIT('h70)
	) name9983 (
		_w4700_,
		_w7014_,
		_w10016_,
		_w10017_
	);
	LUT4 #(
		.INIT('h95aa)
	) name9984 (
		\a[11] ,
		_w4459_,
		_w7291_,
		_w10017_,
		_w10018_
	);
	LUT2 #(
		.INIT('h9)
	) name9985 (
		_w9945_,
		_w9947_,
		_w10019_
	);
	LUT2 #(
		.INIT('h4)
	) name9986 (
		_w10018_,
		_w10019_,
		_w10020_
	);
	LUT3 #(
		.INIT('h82)
	) name9987 (
		_w4459_,
		_w7111_,
		_w7113_,
		_w10021_
	);
	LUT3 #(
		.INIT('h82)
	) name9988 (
		_w4700_,
		_w6960_,
		_w6962_,
		_w10022_
	);
	LUT2 #(
		.INIT('h8)
	) name9989 (
		_w4458_,
		_w7020_,
		_w10023_
	);
	LUT4 #(
		.INIT('h5060)
	) name9990 (
		_w3409_,
		_w3650_,
		_w4684_,
		_w6959_,
		_w10024_
	);
	LUT2 #(
		.INIT('h1)
	) name9991 (
		_w10023_,
		_w10024_,
		_w10025_
	);
	LUT2 #(
		.INIT('h4)
	) name9992 (
		_w10022_,
		_w10025_,
		_w10026_
	);
	LUT3 #(
		.INIT('h1e)
	) name9993 (
		_w9766_,
		_w9943_,
		_w9944_,
		_w10027_
	);
	LUT4 #(
		.INIT('h6500)
	) name9994 (
		\a[11] ,
		_w10021_,
		_w10026_,
		_w10027_,
		_w10028_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9995 (
		_w4459_,
		_w7022_,
		_w7109_,
		_w7110_,
		_w10029_
	);
	LUT4 #(
		.INIT('h5060)
	) name9996 (
		_w3409_,
		_w3650_,
		_w4700_,
		_w6959_,
		_w10030_
	);
	LUT3 #(
		.INIT('h84)
	) name9997 (
		_w3706_,
		_w4458_,
		_w6957_,
		_w10031_
	);
	LUT3 #(
		.INIT('h07)
	) name9998 (
		_w4684_,
		_w7020_,
		_w10031_,
		_w10032_
	);
	LUT2 #(
		.INIT('h4)
	) name9999 (
		_w10030_,
		_w10032_,
		_w10033_
	);
	LUT4 #(
		.INIT('h54ab)
	) name10000 (
		_w9772_,
		_w9939_,
		_w9940_,
		_w9942_,
		_w10034_
	);
	LUT4 #(
		.INIT('h6500)
	) name10001 (
		\a[11] ,
		_w10029_,
		_w10033_,
		_w10034_,
		_w10035_
	);
	LUT4 #(
		.INIT('h04c8)
	) name10002 (
		_w3882_,
		_w4458_,
		_w6954_,
		_w6956_,
		_w10036_
	);
	LUT4 #(
		.INIT('h007b)
	) name10003 (
		_w3706_,
		_w4684_,
		_w6957_,
		_w10036_,
		_w10037_
	);
	LUT3 #(
		.INIT('h70)
	) name10004 (
		_w4700_,
		_w7020_,
		_w10037_,
		_w10038_
	);
	LUT4 #(
		.INIT('h95aa)
	) name10005 (
		\a[11] ,
		_w4459_,
		_w7465_,
		_w10038_,
		_w10039_
	);
	LUT2 #(
		.INIT('h9)
	) name10006 (
		_w9939_,
		_w9941_,
		_w10040_
	);
	LUT2 #(
		.INIT('h4)
	) name10007 (
		_w10039_,
		_w10040_,
		_w10041_
	);
	LUT3 #(
		.INIT('h82)
	) name10008 (
		_w4459_,
		_w7105_,
		_w7107_,
		_w10042_
	);
	LUT3 #(
		.INIT('h84)
	) name10009 (
		_w3706_,
		_w4700_,
		_w6957_,
		_w10043_
	);
	LUT2 #(
		.INIT('h8)
	) name10010 (
		_w4458_,
		_w7026_,
		_w10044_
	);
	LUT4 #(
		.INIT('h04c8)
	) name10011 (
		_w3882_,
		_w4684_,
		_w6954_,
		_w6956_,
		_w10045_
	);
	LUT2 #(
		.INIT('h1)
	) name10012 (
		_w10044_,
		_w10045_,
		_w10046_
	);
	LUT2 #(
		.INIT('h4)
	) name10013 (
		_w10043_,
		_w10046_,
		_w10047_
	);
	LUT3 #(
		.INIT('h1e)
	) name10014 (
		_w9787_,
		_w9937_,
		_w9938_,
		_w10048_
	);
	LUT4 #(
		.INIT('h6500)
	) name10015 (
		\a[11] ,
		_w10042_,
		_w10047_,
		_w10048_,
		_w10049_
	);
	LUT4 #(
		.INIT('h54ab)
	) name10016 (
		_w9793_,
		_w9933_,
		_w9934_,
		_w9936_,
		_w10050_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10017 (
		_w4459_,
		_w7028_,
		_w7103_,
		_w7104_,
		_w10051_
	);
	LUT4 #(
		.INIT('h04c8)
	) name10018 (
		_w3882_,
		_w4700_,
		_w6954_,
		_w6956_,
		_w10052_
	);
	LUT3 #(
		.INIT('h84)
	) name10019 (
		_w4030_,
		_w4458_,
		_w6952_,
		_w10053_
	);
	LUT3 #(
		.INIT('h07)
	) name10020 (
		_w4684_,
		_w7026_,
		_w10053_,
		_w10054_
	);
	LUT2 #(
		.INIT('h4)
	) name10021 (
		_w10052_,
		_w10054_,
		_w10055_
	);
	LUT4 #(
		.INIT('h4844)
	) name10022 (
		\a[11] ,
		_w10050_,
		_w10051_,
		_w10055_,
		_w10056_
	);
	LUT2 #(
		.INIT('h9)
	) name10023 (
		_w9933_,
		_w9935_,
		_w10057_
	);
	LUT4 #(
		.INIT('h5060)
	) name10024 (
		_w4099_,
		_w4378_,
		_w4458_,
		_w6951_,
		_w10058_
	);
	LUT4 #(
		.INIT('h007b)
	) name10025 (
		_w4030_,
		_w4684_,
		_w6952_,
		_w10058_,
		_w10059_
	);
	LUT3 #(
		.INIT('h70)
	) name10026 (
		_w4700_,
		_w7026_,
		_w10059_,
		_w10060_
	);
	LUT4 #(
		.INIT('h95aa)
	) name10027 (
		\a[11] ,
		_w4459_,
		_w7562_,
		_w10060_,
		_w10061_
	);
	LUT2 #(
		.INIT('h2)
	) name10028 (
		_w10057_,
		_w10061_,
		_w10062_
	);
	LUT3 #(
		.INIT('h82)
	) name10029 (
		_w4459_,
		_w7099_,
		_w7101_,
		_w10063_
	);
	LUT3 #(
		.INIT('h84)
	) name10030 (
		_w4030_,
		_w4700_,
		_w6952_,
		_w10064_
	);
	LUT2 #(
		.INIT('h8)
	) name10031 (
		_w4458_,
		_w7032_,
		_w10065_
	);
	LUT4 #(
		.INIT('h5060)
	) name10032 (
		_w4099_,
		_w4378_,
		_w4684_,
		_w6951_,
		_w10066_
	);
	LUT2 #(
		.INIT('h1)
	) name10033 (
		_w10065_,
		_w10066_,
		_w10067_
	);
	LUT2 #(
		.INIT('h4)
	) name10034 (
		_w10064_,
		_w10067_,
		_w10068_
	);
	LUT3 #(
		.INIT('h1e)
	) name10035 (
		_w9808_,
		_w9931_,
		_w9932_,
		_w10069_
	);
	LUT4 #(
		.INIT('h6500)
	) name10036 (
		\a[11] ,
		_w10063_,
		_w10068_,
		_w10069_,
		_w10070_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10037 (
		_w4459_,
		_w7034_,
		_w7097_,
		_w7098_,
		_w10071_
	);
	LUT4 #(
		.INIT('h5060)
	) name10038 (
		_w4099_,
		_w4378_,
		_w4700_,
		_w6951_,
		_w10072_
	);
	LUT3 #(
		.INIT('h82)
	) name10039 (
		_w4458_,
		_w6947_,
		_w6949_,
		_w10073_
	);
	LUT3 #(
		.INIT('h07)
	) name10040 (
		_w4684_,
		_w7032_,
		_w10073_,
		_w10074_
	);
	LUT2 #(
		.INIT('h4)
	) name10041 (
		_w10072_,
		_w10074_,
		_w10075_
	);
	LUT4 #(
		.INIT('h54ab)
	) name10042 (
		_w9814_,
		_w9927_,
		_w9928_,
		_w9930_,
		_w10076_
	);
	LUT4 #(
		.INIT('h6500)
	) name10043 (
		\a[11] ,
		_w10071_,
		_w10075_,
		_w10076_,
		_w10077_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10044 (
		_w4458_,
		_w4695_,
		_w6944_,
		_w6946_,
		_w10078_
	);
	LUT4 #(
		.INIT('h007d)
	) name10045 (
		_w4684_,
		_w6947_,
		_w6949_,
		_w10078_,
		_w10079_
	);
	LUT3 #(
		.INIT('h70)
	) name10046 (
		_w4700_,
		_w7032_,
		_w10079_,
		_w10080_
	);
	LUT4 #(
		.INIT('h95aa)
	) name10047 (
		\a[11] ,
		_w4459_,
		_w7882_,
		_w10080_,
		_w10081_
	);
	LUT2 #(
		.INIT('h9)
	) name10048 (
		_w9927_,
		_w9929_,
		_w10082_
	);
	LUT2 #(
		.INIT('h4)
	) name10049 (
		_w10081_,
		_w10082_,
		_w10083_
	);
	LUT3 #(
		.INIT('h1e)
	) name10050 (
		_w9829_,
		_w9925_,
		_w9926_,
		_w10084_
	);
	LUT3 #(
		.INIT('h82)
	) name10051 (
		_w4459_,
		_w7093_,
		_w7095_,
		_w10085_
	);
	LUT3 #(
		.INIT('h82)
	) name10052 (
		_w4700_,
		_w6947_,
		_w6949_,
		_w10086_
	);
	LUT2 #(
		.INIT('h8)
	) name10053 (
		_w4458_,
		_w7038_,
		_w10087_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10054 (
		_w4684_,
		_w4695_,
		_w6944_,
		_w6946_,
		_w10088_
	);
	LUT2 #(
		.INIT('h1)
	) name10055 (
		_w10087_,
		_w10088_,
		_w10089_
	);
	LUT2 #(
		.INIT('h4)
	) name10056 (
		_w10086_,
		_w10089_,
		_w10090_
	);
	LUT4 #(
		.INIT('h4844)
	) name10057 (
		\a[11] ,
		_w10084_,
		_w10085_,
		_w10090_,
		_w10091_
	);
	LUT4 #(
		.INIT('h54ab)
	) name10058 (
		_w9835_,
		_w9921_,
		_w9922_,
		_w9924_,
		_w10092_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10059 (
		_w4459_,
		_w7040_,
		_w7091_,
		_w7092_,
		_w10093_
	);
	LUT4 #(
		.INIT('h04c8)
	) name10060 (
		_w4695_,
		_w4700_,
		_w6944_,
		_w6946_,
		_w10094_
	);
	LUT3 #(
		.INIT('h82)
	) name10061 (
		_w4458_,
		_w6940_,
		_w6942_,
		_w10095_
	);
	LUT3 #(
		.INIT('h07)
	) name10062 (
		_w4684_,
		_w7038_,
		_w10095_,
		_w10096_
	);
	LUT2 #(
		.INIT('h4)
	) name10063 (
		_w10094_,
		_w10096_,
		_w10097_
	);
	LUT4 #(
		.INIT('h4844)
	) name10064 (
		\a[11] ,
		_w10092_,
		_w10093_,
		_w10097_,
		_w10098_
	);
	LUT2 #(
		.INIT('h9)
	) name10065 (
		_w9921_,
		_w9923_,
		_w10099_
	);
	LUT4 #(
		.INIT('h2228)
	) name10066 (
		_w4458_,
		_w5067_,
		_w5282_,
		_w6939_,
		_w10100_
	);
	LUT4 #(
		.INIT('h007d)
	) name10067 (
		_w4684_,
		_w6940_,
		_w6942_,
		_w10100_,
		_w10101_
	);
	LUT3 #(
		.INIT('h70)
	) name10068 (
		_w4700_,
		_w7038_,
		_w10101_,
		_w10102_
	);
	LUT4 #(
		.INIT('h95aa)
	) name10069 (
		\a[11] ,
		_w4459_,
		_w8018_,
		_w10102_,
		_w10103_
	);
	LUT2 #(
		.INIT('h2)
	) name10070 (
		_w10099_,
		_w10103_,
		_w10104_
	);
	LUT3 #(
		.INIT('h82)
	) name10071 (
		_w4459_,
		_w7087_,
		_w7089_,
		_w10105_
	);
	LUT3 #(
		.INIT('h82)
	) name10072 (
		_w4700_,
		_w6940_,
		_w6942_,
		_w10106_
	);
	LUT2 #(
		.INIT('h8)
	) name10073 (
		_w4458_,
		_w7044_,
		_w10107_
	);
	LUT4 #(
		.INIT('h2228)
	) name10074 (
		_w4684_,
		_w5067_,
		_w5282_,
		_w6939_,
		_w10108_
	);
	LUT2 #(
		.INIT('h1)
	) name10075 (
		_w10107_,
		_w10108_,
		_w10109_
	);
	LUT2 #(
		.INIT('h4)
	) name10076 (
		_w10106_,
		_w10109_,
		_w10110_
	);
	LUT3 #(
		.INIT('h1e)
	) name10077 (
		_w9850_,
		_w9919_,
		_w9920_,
		_w10111_
	);
	LUT4 #(
		.INIT('h6500)
	) name10078 (
		\a[11] ,
		_w10105_,
		_w10110_,
		_w10111_,
		_w10112_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10079 (
		_w4459_,
		_w7046_,
		_w7085_,
		_w7086_,
		_w10113_
	);
	LUT4 #(
		.INIT('h2228)
	) name10080 (
		_w4700_,
		_w5067_,
		_w5282_,
		_w6939_,
		_w10114_
	);
	LUT3 #(
		.INIT('h82)
	) name10081 (
		_w4458_,
		_w6935_,
		_w6937_,
		_w10115_
	);
	LUT3 #(
		.INIT('h07)
	) name10082 (
		_w4684_,
		_w7044_,
		_w10115_,
		_w10116_
	);
	LUT2 #(
		.INIT('h4)
	) name10083 (
		_w10114_,
		_w10116_,
		_w10117_
	);
	LUT4 #(
		.INIT('h54ab)
	) name10084 (
		_w9856_,
		_w9915_,
		_w9916_,
		_w9918_,
		_w10118_
	);
	LUT4 #(
		.INIT('h6500)
	) name10085 (
		\a[11] ,
		_w10113_,
		_w10117_,
		_w10118_,
		_w10119_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10086 (
		_w4458_,
		_w6043_,
		_w6933_,
		_w6934_,
		_w10120_
	);
	LUT4 #(
		.INIT('h007d)
	) name10087 (
		_w4684_,
		_w6935_,
		_w6937_,
		_w10120_,
		_w10121_
	);
	LUT3 #(
		.INIT('h70)
	) name10088 (
		_w4700_,
		_w7044_,
		_w10121_,
		_w10122_
	);
	LUT4 #(
		.INIT('h95aa)
	) name10089 (
		\a[11] ,
		_w4459_,
		_w8005_,
		_w10122_,
		_w10123_
	);
	LUT2 #(
		.INIT('h9)
	) name10090 (
		_w9915_,
		_w9917_,
		_w10124_
	);
	LUT2 #(
		.INIT('h4)
	) name10091 (
		_w10123_,
		_w10124_,
		_w10125_
	);
	LUT3 #(
		.INIT('h1e)
	) name10092 (
		_w9871_,
		_w9913_,
		_w9914_,
		_w10126_
	);
	LUT3 #(
		.INIT('h82)
	) name10093 (
		_w4459_,
		_w7081_,
		_w7083_,
		_w10127_
	);
	LUT3 #(
		.INIT('h82)
	) name10094 (
		_w4700_,
		_w6935_,
		_w6937_,
		_w10128_
	);
	LUT2 #(
		.INIT('h8)
	) name10095 (
		_w4458_,
		_w7050_,
		_w10129_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10096 (
		_w4684_,
		_w6043_,
		_w6933_,
		_w6934_,
		_w10130_
	);
	LUT2 #(
		.INIT('h1)
	) name10097 (
		_w10129_,
		_w10130_,
		_w10131_
	);
	LUT2 #(
		.INIT('h4)
	) name10098 (
		_w10128_,
		_w10131_,
		_w10132_
	);
	LUT4 #(
		.INIT('h4844)
	) name10099 (
		\a[11] ,
		_w10126_,
		_w10127_,
		_w10132_,
		_w10133_
	);
	LUT4 #(
		.INIT('h54ab)
	) name10100 (
		_w9878_,
		_w9909_,
		_w9910_,
		_w9912_,
		_w10134_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10101 (
		_w4459_,
		_w7052_,
		_w7079_,
		_w7080_,
		_w10135_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10102 (
		_w4700_,
		_w6043_,
		_w6933_,
		_w6934_,
		_w10136_
	);
	LUT3 #(
		.INIT('h82)
	) name10103 (
		_w4458_,
		_w6929_,
		_w6931_,
		_w10137_
	);
	LUT3 #(
		.INIT('h07)
	) name10104 (
		_w4684_,
		_w7050_,
		_w10137_,
		_w10138_
	);
	LUT2 #(
		.INIT('h4)
	) name10105 (
		_w10136_,
		_w10138_,
		_w10139_
	);
	LUT4 #(
		.INIT('h4844)
	) name10106 (
		\a[11] ,
		_w10134_,
		_w10135_,
		_w10139_,
		_w10140_
	);
	LUT2 #(
		.INIT('h9)
	) name10107 (
		_w9909_,
		_w9911_,
		_w10141_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10108 (
		_w4458_,
		_w6645_,
		_w6926_,
		_w6928_,
		_w10142_
	);
	LUT4 #(
		.INIT('h007d)
	) name10109 (
		_w4684_,
		_w6929_,
		_w6931_,
		_w10142_,
		_w10143_
	);
	LUT3 #(
		.INIT('h70)
	) name10110 (
		_w4700_,
		_w7050_,
		_w10143_,
		_w10144_
	);
	LUT4 #(
		.INIT('h95aa)
	) name10111 (
		\a[11] ,
		_w4459_,
		_w8227_,
		_w10144_,
		_w10145_
	);
	LUT2 #(
		.INIT('h2)
	) name10112 (
		_w10141_,
		_w10145_,
		_w10146_
	);
	LUT3 #(
		.INIT('h82)
	) name10113 (
		_w4459_,
		_w7075_,
		_w7077_,
		_w10147_
	);
	LUT3 #(
		.INIT('h82)
	) name10114 (
		_w4700_,
		_w6929_,
		_w6931_,
		_w10148_
	);
	LUT2 #(
		.INIT('h8)
	) name10115 (
		_w4458_,
		_w7056_,
		_w10149_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10116 (
		_w4684_,
		_w6645_,
		_w6926_,
		_w6928_,
		_w10150_
	);
	LUT2 #(
		.INIT('h1)
	) name10117 (
		_w10149_,
		_w10150_,
		_w10151_
	);
	LUT2 #(
		.INIT('h4)
	) name10118 (
		_w10148_,
		_w10151_,
		_w10152_
	);
	LUT2 #(
		.INIT('h9)
	) name10119 (
		_w9906_,
		_w9908_,
		_w10153_
	);
	LUT4 #(
		.INIT('h6500)
	) name10120 (
		\a[11] ,
		_w10147_,
		_w10152_,
		_w10153_,
		_w10154_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10121 (
		_w4459_,
		_w7058_,
		_w7073_,
		_w7074_,
		_w10155_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10122 (
		_w4700_,
		_w6645_,
		_w6926_,
		_w6928_,
		_w10156_
	);
	LUT3 #(
		.INIT('h82)
	) name10123 (
		_w4458_,
		_w6922_,
		_w6924_,
		_w10157_
	);
	LUT3 #(
		.INIT('h07)
	) name10124 (
		_w4684_,
		_w7056_,
		_w10157_,
		_w10158_
	);
	LUT2 #(
		.INIT('h4)
	) name10125 (
		_w10156_,
		_w10158_,
		_w10159_
	);
	LUT4 #(
		.INIT('h9a65)
	) name10126 (
		\a[14] ,
		_w9899_,
		_w9903_,
		_w9904_,
		_w10160_
	);
	LUT4 #(
		.INIT('h6500)
	) name10127 (
		\a[11] ,
		_w10155_,
		_w10159_,
		_w10160_,
		_w10161_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10128 (
		_w4458_,
		_w6669_,
		_w6919_,
		_w6921_,
		_w10162_
	);
	LUT4 #(
		.INIT('h007d)
	) name10129 (
		_w4684_,
		_w6922_,
		_w6924_,
		_w10162_,
		_w10163_
	);
	LUT3 #(
		.INIT('h70)
	) name10130 (
		_w4700_,
		_w7056_,
		_w10163_,
		_w10164_
	);
	LUT4 #(
		.INIT('h95aa)
	) name10131 (
		\a[11] ,
		_w4459_,
		_w8298_,
		_w10164_,
		_w10165_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name10132 (
		\a[14] ,
		_w9891_,
		_w9888_,
		_w9890_,
		_w10166_
	);
	LUT3 #(
		.INIT('h4b)
	) name10133 (
		_w9894_,
		_w9897_,
		_w10166_,
		_w10167_
	);
	LUT2 #(
		.INIT('h4)
	) name10134 (
		_w10165_,
		_w10167_,
		_w10168_
	);
	LUT3 #(
		.INIT('h82)
	) name10135 (
		_w4459_,
		_w7069_,
		_w7071_,
		_w10169_
	);
	LUT3 #(
		.INIT('h82)
	) name10136 (
		_w4700_,
		_w6922_,
		_w6924_,
		_w10170_
	);
	LUT2 #(
		.INIT('h8)
	) name10137 (
		_w4458_,
		_w7062_,
		_w10171_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10138 (
		_w4684_,
		_w6669_,
		_w6919_,
		_w6921_,
		_w10172_
	);
	LUT2 #(
		.INIT('h1)
	) name10139 (
		_w10171_,
		_w10172_,
		_w10173_
	);
	LUT2 #(
		.INIT('h4)
	) name10140 (
		_w10170_,
		_w10173_,
		_w10174_
	);
	LUT2 #(
		.INIT('h8)
	) name10141 (
		\a[14] ,
		_w9891_,
		_w10175_
	);
	LUT3 #(
		.INIT('h4b)
	) name10142 (
		_w9888_,
		_w9890_,
		_w10175_,
		_w10176_
	);
	LUT4 #(
		.INIT('h6500)
	) name10143 (
		\a[11] ,
		_w10169_,
		_w10174_,
		_w10176_,
		_w10177_
	);
	LUT4 #(
		.INIT('h2882)
	) name10144 (
		_w4459_,
		_w6914_,
		_w6916_,
		_w7067_,
		_w10178_
	);
	LUT4 #(
		.INIT('ha802)
	) name10145 (
		_w4684_,
		_w6689_,
		_w6911_,
		_w6913_,
		_w10179_
	);
	LUT4 #(
		.INIT('h007d)
	) name10146 (
		_w4700_,
		_w6914_,
		_w6916_,
		_w10179_,
		_w10180_
	);
	LUT4 #(
		.INIT('h5401)
	) name10147 (
		_w4457_,
		_w6689_,
		_w6911_,
		_w6913_,
		_w10181_
	);
	LUT2 #(
		.INIT('h2)
	) name10148 (
		\a[11] ,
		_w10181_,
		_w10182_
	);
	LUT3 #(
		.INIT('h40)
	) name10149 (
		_w10178_,
		_w10180_,
		_w10182_,
		_w10183_
	);
	LUT3 #(
		.INIT('h28)
	) name10150 (
		_w4459_,
		_w7062_,
		_w8358_,
		_w10184_
	);
	LUT4 #(
		.INIT('ha802)
	) name10151 (
		_w4458_,
		_w6689_,
		_w6911_,
		_w6913_,
		_w10185_
	);
	LUT4 #(
		.INIT('h007d)
	) name10152 (
		_w4684_,
		_w6914_,
		_w6916_,
		_w10185_,
		_w10186_
	);
	LUT3 #(
		.INIT('h70)
	) name10153 (
		_w4700_,
		_w7062_,
		_w10186_,
		_w10187_
	);
	LUT4 #(
		.INIT('h0800)
	) name10154 (
		_w9891_,
		_w10183_,
		_w10184_,
		_w10187_,
		_w10188_
	);
	LUT3 #(
		.INIT('h28)
	) name10155 (
		_w4459_,
		_w7065_,
		_w7068_,
		_w10189_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10156 (
		_w4700_,
		_w6669_,
		_w6919_,
		_w6921_,
		_w10190_
	);
	LUT3 #(
		.INIT('h82)
	) name10157 (
		_w4458_,
		_w6914_,
		_w6916_,
		_w10191_
	);
	LUT3 #(
		.INIT('h07)
	) name10158 (
		_w4684_,
		_w7062_,
		_w10191_,
		_w10192_
	);
	LUT2 #(
		.INIT('h4)
	) name10159 (
		_w10190_,
		_w10192_,
		_w10193_
	);
	LUT4 #(
		.INIT('ha6aa)
	) name10160 (
		_w9891_,
		_w10183_,
		_w10184_,
		_w10187_,
		_w10194_
	);
	LUT4 #(
		.INIT('h6500)
	) name10161 (
		\a[11] ,
		_w10189_,
		_w10193_,
		_w10194_,
		_w10195_
	);
	LUT2 #(
		.INIT('h1)
	) name10162 (
		_w10188_,
		_w10195_,
		_w10196_
	);
	LUT4 #(
		.INIT('h009a)
	) name10163 (
		\a[11] ,
		_w10169_,
		_w10174_,
		_w10176_,
		_w10197_
	);
	LUT4 #(
		.INIT('h9a65)
	) name10164 (
		\a[11] ,
		_w10169_,
		_w10174_,
		_w10176_,
		_w10198_
	);
	LUT3 #(
		.INIT('h54)
	) name10165 (
		_w10177_,
		_w10196_,
		_w10197_,
		_w10199_
	);
	LUT2 #(
		.INIT('h2)
	) name10166 (
		_w10165_,
		_w10167_,
		_w10200_
	);
	LUT2 #(
		.INIT('h9)
	) name10167 (
		_w10165_,
		_w10167_,
		_w10201_
	);
	LUT4 #(
		.INIT('h9a65)
	) name10168 (
		\a[11] ,
		_w10155_,
		_w10159_,
		_w10160_,
		_w10202_
	);
	LUT4 #(
		.INIT('h4d00)
	) name10169 (
		_w10165_,
		_w10167_,
		_w10199_,
		_w10202_,
		_w10203_
	);
	LUT4 #(
		.INIT('h9a65)
	) name10170 (
		\a[11] ,
		_w10147_,
		_w10152_,
		_w10153_,
		_w10204_
	);
	LUT4 #(
		.INIT('h0155)
	) name10171 (
		_w10154_,
		_w10161_,
		_w10203_,
		_w10204_,
		_w10205_
	);
	LUT2 #(
		.INIT('h4)
	) name10172 (
		_w10141_,
		_w10145_,
		_w10206_
	);
	LUT2 #(
		.INIT('h9)
	) name10173 (
		_w10141_,
		_w10145_,
		_w10207_
	);
	LUT4 #(
		.INIT('h9699)
	) name10174 (
		\a[11] ,
		_w10134_,
		_w10135_,
		_w10139_,
		_w10208_
	);
	LUT4 #(
		.INIT('h2b00)
	) name10175 (
		_w10141_,
		_w10145_,
		_w10205_,
		_w10208_,
		_w10209_
	);
	LUT4 #(
		.INIT('h9699)
	) name10176 (
		\a[11] ,
		_w10126_,
		_w10127_,
		_w10132_,
		_w10210_
	);
	LUT4 #(
		.INIT('h0155)
	) name10177 (
		_w10133_,
		_w10140_,
		_w10209_,
		_w10210_,
		_w10211_
	);
	LUT2 #(
		.INIT('h2)
	) name10178 (
		_w10123_,
		_w10124_,
		_w10212_
	);
	LUT2 #(
		.INIT('h9)
	) name10179 (
		_w10123_,
		_w10124_,
		_w10213_
	);
	LUT4 #(
		.INIT('h9a65)
	) name10180 (
		\a[11] ,
		_w10113_,
		_w10117_,
		_w10118_,
		_w10214_
	);
	LUT4 #(
		.INIT('h4d00)
	) name10181 (
		_w10123_,
		_w10124_,
		_w10211_,
		_w10214_,
		_w10215_
	);
	LUT4 #(
		.INIT('h9a65)
	) name10182 (
		\a[11] ,
		_w10105_,
		_w10110_,
		_w10111_,
		_w10216_
	);
	LUT4 #(
		.INIT('h0155)
	) name10183 (
		_w10112_,
		_w10119_,
		_w10215_,
		_w10216_,
		_w10217_
	);
	LUT2 #(
		.INIT('h4)
	) name10184 (
		_w10099_,
		_w10103_,
		_w10218_
	);
	LUT2 #(
		.INIT('h9)
	) name10185 (
		_w10099_,
		_w10103_,
		_w10219_
	);
	LUT4 #(
		.INIT('h9699)
	) name10186 (
		\a[11] ,
		_w10092_,
		_w10093_,
		_w10097_,
		_w10220_
	);
	LUT4 #(
		.INIT('h2b00)
	) name10187 (
		_w10099_,
		_w10103_,
		_w10217_,
		_w10220_,
		_w10221_
	);
	LUT4 #(
		.INIT('h9699)
	) name10188 (
		\a[11] ,
		_w10084_,
		_w10085_,
		_w10090_,
		_w10222_
	);
	LUT4 #(
		.INIT('h0155)
	) name10189 (
		_w10091_,
		_w10098_,
		_w10221_,
		_w10222_,
		_w10223_
	);
	LUT2 #(
		.INIT('h2)
	) name10190 (
		_w10081_,
		_w10082_,
		_w10224_
	);
	LUT2 #(
		.INIT('h9)
	) name10191 (
		_w10081_,
		_w10082_,
		_w10225_
	);
	LUT4 #(
		.INIT('h9a65)
	) name10192 (
		\a[11] ,
		_w10071_,
		_w10075_,
		_w10076_,
		_w10226_
	);
	LUT4 #(
		.INIT('h4d00)
	) name10193 (
		_w10081_,
		_w10082_,
		_w10223_,
		_w10226_,
		_w10227_
	);
	LUT4 #(
		.INIT('h9a65)
	) name10194 (
		\a[11] ,
		_w10063_,
		_w10068_,
		_w10069_,
		_w10228_
	);
	LUT4 #(
		.INIT('h0155)
	) name10195 (
		_w10070_,
		_w10077_,
		_w10227_,
		_w10228_,
		_w10229_
	);
	LUT2 #(
		.INIT('h4)
	) name10196 (
		_w10057_,
		_w10061_,
		_w10230_
	);
	LUT2 #(
		.INIT('h9)
	) name10197 (
		_w10057_,
		_w10061_,
		_w10231_
	);
	LUT4 #(
		.INIT('h9699)
	) name10198 (
		\a[11] ,
		_w10050_,
		_w10051_,
		_w10055_,
		_w10232_
	);
	LUT4 #(
		.INIT('h2b00)
	) name10199 (
		_w10057_,
		_w10061_,
		_w10229_,
		_w10232_,
		_w10233_
	);
	LUT4 #(
		.INIT('h9a65)
	) name10200 (
		\a[11] ,
		_w10042_,
		_w10047_,
		_w10048_,
		_w10234_
	);
	LUT4 #(
		.INIT('h0155)
	) name10201 (
		_w10049_,
		_w10056_,
		_w10233_,
		_w10234_,
		_w10235_
	);
	LUT2 #(
		.INIT('h2)
	) name10202 (
		_w10039_,
		_w10040_,
		_w10236_
	);
	LUT2 #(
		.INIT('h9)
	) name10203 (
		_w10039_,
		_w10040_,
		_w10237_
	);
	LUT4 #(
		.INIT('h9a65)
	) name10204 (
		\a[11] ,
		_w10029_,
		_w10033_,
		_w10034_,
		_w10238_
	);
	LUT4 #(
		.INIT('h4d00)
	) name10205 (
		_w10039_,
		_w10040_,
		_w10235_,
		_w10238_,
		_w10239_
	);
	LUT4 #(
		.INIT('h9a65)
	) name10206 (
		\a[11] ,
		_w10021_,
		_w10026_,
		_w10027_,
		_w10240_
	);
	LUT4 #(
		.INIT('h0155)
	) name10207 (
		_w10028_,
		_w10035_,
		_w10239_,
		_w10240_,
		_w10241_
	);
	LUT2 #(
		.INIT('h2)
	) name10208 (
		_w10018_,
		_w10019_,
		_w10242_
	);
	LUT2 #(
		.INIT('h9)
	) name10209 (
		_w10018_,
		_w10019_,
		_w10243_
	);
	LUT4 #(
		.INIT('h9a65)
	) name10210 (
		\a[11] ,
		_w10008_,
		_w10012_,
		_w10013_,
		_w10244_
	);
	LUT4 #(
		.INIT('h4d00)
	) name10211 (
		_w10018_,
		_w10019_,
		_w10241_,
		_w10244_,
		_w10245_
	);
	LUT4 #(
		.INIT('h9a65)
	) name10212 (
		\a[11] ,
		_w10000_,
		_w10005_,
		_w10006_,
		_w10246_
	);
	LUT4 #(
		.INIT('h0155)
	) name10213 (
		_w10007_,
		_w10014_,
		_w10245_,
		_w10246_,
		_w10247_
	);
	LUT2 #(
		.INIT('h2)
	) name10214 (
		_w9997_,
		_w9998_,
		_w10248_
	);
	LUT2 #(
		.INIT('h9)
	) name10215 (
		_w9997_,
		_w9998_,
		_w10249_
	);
	LUT4 #(
		.INIT('h9a65)
	) name10216 (
		\a[11] ,
		_w9987_,
		_w9991_,
		_w9992_,
		_w10250_
	);
	LUT4 #(
		.INIT('h4d00)
	) name10217 (
		_w9997_,
		_w9998_,
		_w10247_,
		_w10250_,
		_w10251_
	);
	LUT4 #(
		.INIT('h9a65)
	) name10218 (
		\a[11] ,
		_w9979_,
		_w9984_,
		_w9985_,
		_w10252_
	);
	LUT4 #(
		.INIT('h0155)
	) name10219 (
		_w9986_,
		_w9993_,
		_w10251_,
		_w10252_,
		_w10253_
	);
	LUT4 #(
		.INIT('h6996)
	) name10220 (
		_w9673_,
		_w9674_,
		_w9678_,
		_w9957_,
		_w10254_
	);
	LUT4 #(
		.INIT('h04c8)
	) name10221 (
		_w2622_,
		_w4875_,
		_w6978_,
		_w6980_,
		_w10255_
	);
	LUT4 #(
		.INIT('h007b)
	) name10222 (
		_w2546_,
		_w5271_,
		_w6981_,
		_w10255_,
		_w10256_
	);
	LUT3 #(
		.INIT('h70)
	) name10223 (
		_w5286_,
		_w6996_,
		_w10256_,
		_w10257_
	);
	LUT4 #(
		.INIT('h95aa)
	) name10224 (
		\a[8] ,
		_w4876_,
		_w7500_,
		_w10257_,
		_w10258_
	);
	LUT4 #(
		.INIT('hde48)
	) name10225 (
		_w9963_,
		_w10253_,
		_w10254_,
		_w10258_,
		_w10259_
	);
	LUT4 #(
		.INIT('h0a02)
	) name10226 (
		_w35_,
		_w7169_,
		_w7419_,
		_w7686_,
		_w10260_
	);
	LUT3 #(
		.INIT('h28)
	) name10227 (
		_w5524_,
		_w7136_,
		_w7168_,
		_w10261_
	);
	LUT3 #(
		.INIT('h40)
	) name10228 (
		_w6324_,
		_w7136_,
		_w7167_,
		_w10262_
	);
	LUT3 #(
		.INIT('h31)
	) name10229 (
		_w9705_,
		_w10261_,
		_w10262_,
		_w10263_
	);
	LUT3 #(
		.INIT('h9a)
	) name10230 (
		\a[5] ,
		_w10260_,
		_w10263_,
		_w10264_
	);
	LUT3 #(
		.INIT('hd4)
	) name10231 (
		_w9978_,
		_w10259_,
		_w10264_,
		_w10265_
	);
	LUT3 #(
		.INIT('h06)
	) name10232 (
		_w9974_,
		_w9977_,
		_w10265_,
		_w10266_
	);
	LUT3 #(
		.INIT('h90)
	) name10233 (
		_w9974_,
		_w9977_,
		_w10265_,
		_w10267_
	);
	LUT3 #(
		.INIT('h69)
	) name10234 (
		_w9974_,
		_w9977_,
		_w10265_,
		_w10268_
	);
	LUT3 #(
		.INIT('h1e)
	) name10235 (
		_w9993_,
		_w10251_,
		_w10252_,
		_w10269_
	);
	LUT3 #(
		.INIT('h82)
	) name10236 (
		_w4876_,
		_w7129_,
		_w7131_,
		_w10270_
	);
	LUT3 #(
		.INIT('h84)
	) name10237 (
		_w2546_,
		_w5286_,
		_w6981_,
		_w10271_
	);
	LUT2 #(
		.INIT('h8)
	) name10238 (
		_w4875_,
		_w7002_,
		_w10272_
	);
	LUT4 #(
		.INIT('h04c8)
	) name10239 (
		_w2622_,
		_w5271_,
		_w6978_,
		_w6980_,
		_w10273_
	);
	LUT2 #(
		.INIT('h1)
	) name10240 (
		_w10272_,
		_w10273_,
		_w10274_
	);
	LUT2 #(
		.INIT('h4)
	) name10241 (
		_w10271_,
		_w10274_,
		_w10275_
	);
	LUT4 #(
		.INIT('h4844)
	) name10242 (
		\a[8] ,
		_w10269_,
		_w10270_,
		_w10275_,
		_w10276_
	);
	LUT4 #(
		.INIT('h54ab)
	) name10243 (
		_w9999_,
		_w10247_,
		_w10248_,
		_w10250_,
		_w10277_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10244 (
		_w4876_,
		_w7004_,
		_w7127_,
		_w7128_,
		_w10278_
	);
	LUT4 #(
		.INIT('h04c8)
	) name10245 (
		_w2622_,
		_w5286_,
		_w6978_,
		_w6980_,
		_w10279_
	);
	LUT3 #(
		.INIT('h84)
	) name10246 (
		_w2872_,
		_w4875_,
		_w6975_,
		_w10280_
	);
	LUT3 #(
		.INIT('h07)
	) name10247 (
		_w5271_,
		_w7002_,
		_w10280_,
		_w10281_
	);
	LUT2 #(
		.INIT('h4)
	) name10248 (
		_w10279_,
		_w10281_,
		_w10282_
	);
	LUT4 #(
		.INIT('h4844)
	) name10249 (
		\a[8] ,
		_w10277_,
		_w10278_,
		_w10282_,
		_w10283_
	);
	LUT2 #(
		.INIT('h9)
	) name10250 (
		_w10247_,
		_w10249_,
		_w10284_
	);
	LUT4 #(
		.INIT('h04c8)
	) name10251 (
		_w2983_,
		_w4875_,
		_w6972_,
		_w6974_,
		_w10285_
	);
	LUT4 #(
		.INIT('h007b)
	) name10252 (
		_w2872_,
		_w5271_,
		_w6975_,
		_w10285_,
		_w10286_
	);
	LUT3 #(
		.INIT('h70)
	) name10253 (
		_w5286_,
		_w7002_,
		_w10286_,
		_w10287_
	);
	LUT4 #(
		.INIT('h95aa)
	) name10254 (
		\a[8] ,
		_w4876_,
		_w7426_,
		_w10287_,
		_w10288_
	);
	LUT2 #(
		.INIT('h2)
	) name10255 (
		_w10284_,
		_w10288_,
		_w10289_
	);
	LUT3 #(
		.INIT('h1e)
	) name10256 (
		_w10014_,
		_w10245_,
		_w10246_,
		_w10290_
	);
	LUT3 #(
		.INIT('h82)
	) name10257 (
		_w4876_,
		_w7123_,
		_w7125_,
		_w10291_
	);
	LUT3 #(
		.INIT('h84)
	) name10258 (
		_w2872_,
		_w5286_,
		_w6975_,
		_w10292_
	);
	LUT2 #(
		.INIT('h8)
	) name10259 (
		_w4875_,
		_w7008_,
		_w10293_
	);
	LUT4 #(
		.INIT('h04c8)
	) name10260 (
		_w2983_,
		_w5271_,
		_w6972_,
		_w6974_,
		_w10294_
	);
	LUT2 #(
		.INIT('h1)
	) name10261 (
		_w10293_,
		_w10294_,
		_w10295_
	);
	LUT2 #(
		.INIT('h4)
	) name10262 (
		_w10292_,
		_w10295_,
		_w10296_
	);
	LUT4 #(
		.INIT('h4844)
	) name10263 (
		\a[8] ,
		_w10290_,
		_w10291_,
		_w10296_,
		_w10297_
	);
	LUT4 #(
		.INIT('h54ab)
	) name10264 (
		_w10020_,
		_w10241_,
		_w10242_,
		_w10244_,
		_w10298_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10265 (
		_w4876_,
		_w7010_,
		_w7121_,
		_w7122_,
		_w10299_
	);
	LUT4 #(
		.INIT('h04c8)
	) name10266 (
		_w2983_,
		_w5286_,
		_w6972_,
		_w6974_,
		_w10300_
	);
	LUT3 #(
		.INIT('h82)
	) name10267 (
		_w4875_,
		_w6967_,
		_w6969_,
		_w10301_
	);
	LUT3 #(
		.INIT('h07)
	) name10268 (
		_w5271_,
		_w7008_,
		_w10301_,
		_w10302_
	);
	LUT2 #(
		.INIT('h4)
	) name10269 (
		_w10300_,
		_w10302_,
		_w10303_
	);
	LUT4 #(
		.INIT('h4844)
	) name10270 (
		\a[8] ,
		_w10298_,
		_w10299_,
		_w10303_,
		_w10304_
	);
	LUT2 #(
		.INIT('h9)
	) name10271 (
		_w10241_,
		_w10243_,
		_w10305_
	);
	LUT4 #(
		.INIT('h04c8)
	) name10272 (
		_w3257_,
		_w4875_,
		_w6964_,
		_w6966_,
		_w10306_
	);
	LUT4 #(
		.INIT('h007d)
	) name10273 (
		_w5271_,
		_w6967_,
		_w6969_,
		_w10306_,
		_w10307_
	);
	LUT3 #(
		.INIT('h70)
	) name10274 (
		_w5286_,
		_w7008_,
		_w10307_,
		_w10308_
	);
	LUT4 #(
		.INIT('h95aa)
	) name10275 (
		\a[8] ,
		_w4876_,
		_w7403_,
		_w10308_,
		_w10309_
	);
	LUT2 #(
		.INIT('h2)
	) name10276 (
		_w10305_,
		_w10309_,
		_w10310_
	);
	LUT3 #(
		.INIT('h1e)
	) name10277 (
		_w10035_,
		_w10239_,
		_w10240_,
		_w10311_
	);
	LUT3 #(
		.INIT('h82)
	) name10278 (
		_w4876_,
		_w7117_,
		_w7119_,
		_w10312_
	);
	LUT3 #(
		.INIT('h82)
	) name10279 (
		_w5286_,
		_w6967_,
		_w6969_,
		_w10313_
	);
	LUT2 #(
		.INIT('h8)
	) name10280 (
		_w4875_,
		_w7014_,
		_w10314_
	);
	LUT4 #(
		.INIT('h04c8)
	) name10281 (
		_w3257_,
		_w5271_,
		_w6964_,
		_w6966_,
		_w10315_
	);
	LUT2 #(
		.INIT('h1)
	) name10282 (
		_w10314_,
		_w10315_,
		_w10316_
	);
	LUT2 #(
		.INIT('h4)
	) name10283 (
		_w10313_,
		_w10316_,
		_w10317_
	);
	LUT4 #(
		.INIT('h4844)
	) name10284 (
		\a[8] ,
		_w10311_,
		_w10312_,
		_w10317_,
		_w10318_
	);
	LUT4 #(
		.INIT('h54ab)
	) name10285 (
		_w10041_,
		_w10235_,
		_w10236_,
		_w10238_,
		_w10319_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10286 (
		_w4876_,
		_w7016_,
		_w7115_,
		_w7116_,
		_w10320_
	);
	LUT4 #(
		.INIT('h04c8)
	) name10287 (
		_w3257_,
		_w5286_,
		_w6964_,
		_w6966_,
		_w10321_
	);
	LUT3 #(
		.INIT('h82)
	) name10288 (
		_w4875_,
		_w6960_,
		_w6962_,
		_w10322_
	);
	LUT3 #(
		.INIT('h07)
	) name10289 (
		_w5271_,
		_w7014_,
		_w10322_,
		_w10323_
	);
	LUT2 #(
		.INIT('h4)
	) name10290 (
		_w10321_,
		_w10323_,
		_w10324_
	);
	LUT4 #(
		.INIT('h4844)
	) name10291 (
		\a[8] ,
		_w10319_,
		_w10320_,
		_w10324_,
		_w10325_
	);
	LUT2 #(
		.INIT('h9)
	) name10292 (
		_w10235_,
		_w10237_,
		_w10326_
	);
	LUT4 #(
		.INIT('h5060)
	) name10293 (
		_w3409_,
		_w3650_,
		_w4875_,
		_w6959_,
		_w10327_
	);
	LUT4 #(
		.INIT('h007d)
	) name10294 (
		_w5271_,
		_w6960_,
		_w6962_,
		_w10327_,
		_w10328_
	);
	LUT3 #(
		.INIT('h70)
	) name10295 (
		_w5286_,
		_w7014_,
		_w10328_,
		_w10329_
	);
	LUT4 #(
		.INIT('h95aa)
	) name10296 (
		\a[8] ,
		_w4876_,
		_w7291_,
		_w10329_,
		_w10330_
	);
	LUT2 #(
		.INIT('h2)
	) name10297 (
		_w10326_,
		_w10330_,
		_w10331_
	);
	LUT3 #(
		.INIT('h1e)
	) name10298 (
		_w10056_,
		_w10233_,
		_w10234_,
		_w10332_
	);
	LUT3 #(
		.INIT('h82)
	) name10299 (
		_w4876_,
		_w7111_,
		_w7113_,
		_w10333_
	);
	LUT3 #(
		.INIT('h82)
	) name10300 (
		_w5286_,
		_w6960_,
		_w6962_,
		_w10334_
	);
	LUT2 #(
		.INIT('h8)
	) name10301 (
		_w4875_,
		_w7020_,
		_w10335_
	);
	LUT4 #(
		.INIT('h5060)
	) name10302 (
		_w3409_,
		_w3650_,
		_w5271_,
		_w6959_,
		_w10336_
	);
	LUT2 #(
		.INIT('h1)
	) name10303 (
		_w10335_,
		_w10336_,
		_w10337_
	);
	LUT2 #(
		.INIT('h4)
	) name10304 (
		_w10334_,
		_w10337_,
		_w10338_
	);
	LUT4 #(
		.INIT('h4844)
	) name10305 (
		\a[8] ,
		_w10332_,
		_w10333_,
		_w10338_,
		_w10339_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10306 (
		_w4876_,
		_w7022_,
		_w7109_,
		_w7110_,
		_w10340_
	);
	LUT4 #(
		.INIT('h5060)
	) name10307 (
		_w3409_,
		_w3650_,
		_w5286_,
		_w6959_,
		_w10341_
	);
	LUT3 #(
		.INIT('h84)
	) name10308 (
		_w3706_,
		_w4875_,
		_w6957_,
		_w10342_
	);
	LUT3 #(
		.INIT('h07)
	) name10309 (
		_w5271_,
		_w7020_,
		_w10342_,
		_w10343_
	);
	LUT2 #(
		.INIT('h4)
	) name10310 (
		_w10341_,
		_w10343_,
		_w10344_
	);
	LUT4 #(
		.INIT('h54ab)
	) name10311 (
		_w10062_,
		_w10229_,
		_w10230_,
		_w10232_,
		_w10345_
	);
	LUT4 #(
		.INIT('h6500)
	) name10312 (
		\a[8] ,
		_w10340_,
		_w10344_,
		_w10345_,
		_w10346_
	);
	LUT4 #(
		.INIT('h04c8)
	) name10313 (
		_w3882_,
		_w4875_,
		_w6954_,
		_w6956_,
		_w10347_
	);
	LUT4 #(
		.INIT('h007b)
	) name10314 (
		_w3706_,
		_w5271_,
		_w6957_,
		_w10347_,
		_w10348_
	);
	LUT3 #(
		.INIT('h70)
	) name10315 (
		_w5286_,
		_w7020_,
		_w10348_,
		_w10349_
	);
	LUT4 #(
		.INIT('h95aa)
	) name10316 (
		\a[8] ,
		_w4876_,
		_w7465_,
		_w10349_,
		_w10350_
	);
	LUT2 #(
		.INIT('h9)
	) name10317 (
		_w10229_,
		_w10231_,
		_w10351_
	);
	LUT2 #(
		.INIT('h4)
	) name10318 (
		_w10350_,
		_w10351_,
		_w10352_
	);
	LUT3 #(
		.INIT('h1e)
	) name10319 (
		_w10077_,
		_w10227_,
		_w10228_,
		_w10353_
	);
	LUT3 #(
		.INIT('h82)
	) name10320 (
		_w4876_,
		_w7105_,
		_w7107_,
		_w10354_
	);
	LUT3 #(
		.INIT('h84)
	) name10321 (
		_w3706_,
		_w5286_,
		_w6957_,
		_w10355_
	);
	LUT2 #(
		.INIT('h8)
	) name10322 (
		_w4875_,
		_w7026_,
		_w10356_
	);
	LUT4 #(
		.INIT('h04c8)
	) name10323 (
		_w3882_,
		_w5271_,
		_w6954_,
		_w6956_,
		_w10357_
	);
	LUT2 #(
		.INIT('h1)
	) name10324 (
		_w10356_,
		_w10357_,
		_w10358_
	);
	LUT2 #(
		.INIT('h4)
	) name10325 (
		_w10355_,
		_w10358_,
		_w10359_
	);
	LUT4 #(
		.INIT('h4844)
	) name10326 (
		\a[8] ,
		_w10353_,
		_w10354_,
		_w10359_,
		_w10360_
	);
	LUT4 #(
		.INIT('h54ab)
	) name10327 (
		_w10083_,
		_w10223_,
		_w10224_,
		_w10226_,
		_w10361_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10328 (
		_w4876_,
		_w7028_,
		_w7103_,
		_w7104_,
		_w10362_
	);
	LUT4 #(
		.INIT('h04c8)
	) name10329 (
		_w3882_,
		_w5286_,
		_w6954_,
		_w6956_,
		_w10363_
	);
	LUT3 #(
		.INIT('h84)
	) name10330 (
		_w4030_,
		_w4875_,
		_w6952_,
		_w10364_
	);
	LUT3 #(
		.INIT('h07)
	) name10331 (
		_w5271_,
		_w7026_,
		_w10364_,
		_w10365_
	);
	LUT2 #(
		.INIT('h4)
	) name10332 (
		_w10363_,
		_w10365_,
		_w10366_
	);
	LUT4 #(
		.INIT('h4844)
	) name10333 (
		\a[8] ,
		_w10361_,
		_w10362_,
		_w10366_,
		_w10367_
	);
	LUT2 #(
		.INIT('h9)
	) name10334 (
		_w10223_,
		_w10225_,
		_w10368_
	);
	LUT4 #(
		.INIT('h5060)
	) name10335 (
		_w4099_,
		_w4378_,
		_w4875_,
		_w6951_,
		_w10369_
	);
	LUT4 #(
		.INIT('h007b)
	) name10336 (
		_w4030_,
		_w5271_,
		_w6952_,
		_w10369_,
		_w10370_
	);
	LUT3 #(
		.INIT('h70)
	) name10337 (
		_w5286_,
		_w7026_,
		_w10370_,
		_w10371_
	);
	LUT4 #(
		.INIT('h95aa)
	) name10338 (
		\a[8] ,
		_w4876_,
		_w7562_,
		_w10371_,
		_w10372_
	);
	LUT2 #(
		.INIT('h2)
	) name10339 (
		_w10368_,
		_w10372_,
		_w10373_
	);
	LUT3 #(
		.INIT('h82)
	) name10340 (
		_w4876_,
		_w7099_,
		_w7101_,
		_w10374_
	);
	LUT3 #(
		.INIT('h84)
	) name10341 (
		_w4030_,
		_w5286_,
		_w6952_,
		_w10375_
	);
	LUT2 #(
		.INIT('h8)
	) name10342 (
		_w4875_,
		_w7032_,
		_w10376_
	);
	LUT4 #(
		.INIT('h5060)
	) name10343 (
		_w4099_,
		_w4378_,
		_w5271_,
		_w6951_,
		_w10377_
	);
	LUT2 #(
		.INIT('h1)
	) name10344 (
		_w10376_,
		_w10377_,
		_w10378_
	);
	LUT2 #(
		.INIT('h4)
	) name10345 (
		_w10375_,
		_w10378_,
		_w10379_
	);
	LUT3 #(
		.INIT('h1e)
	) name10346 (
		_w10098_,
		_w10221_,
		_w10222_,
		_w10380_
	);
	LUT4 #(
		.INIT('h6500)
	) name10347 (
		\a[8] ,
		_w10374_,
		_w10379_,
		_w10380_,
		_w10381_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10348 (
		_w4876_,
		_w7034_,
		_w7097_,
		_w7098_,
		_w10382_
	);
	LUT4 #(
		.INIT('h5060)
	) name10349 (
		_w4099_,
		_w4378_,
		_w5286_,
		_w6951_,
		_w10383_
	);
	LUT3 #(
		.INIT('h82)
	) name10350 (
		_w4875_,
		_w6947_,
		_w6949_,
		_w10384_
	);
	LUT3 #(
		.INIT('h07)
	) name10351 (
		_w5271_,
		_w7032_,
		_w10384_,
		_w10385_
	);
	LUT2 #(
		.INIT('h4)
	) name10352 (
		_w10383_,
		_w10385_,
		_w10386_
	);
	LUT4 #(
		.INIT('h54ab)
	) name10353 (
		_w10104_,
		_w10217_,
		_w10218_,
		_w10220_,
		_w10387_
	);
	LUT4 #(
		.INIT('h6500)
	) name10354 (
		\a[8] ,
		_w10382_,
		_w10386_,
		_w10387_,
		_w10388_
	);
	LUT4 #(
		.INIT('h04c8)
	) name10355 (
		_w4695_,
		_w4875_,
		_w6944_,
		_w6946_,
		_w10389_
	);
	LUT4 #(
		.INIT('h007d)
	) name10356 (
		_w5271_,
		_w6947_,
		_w6949_,
		_w10389_,
		_w10390_
	);
	LUT3 #(
		.INIT('h70)
	) name10357 (
		_w5286_,
		_w7032_,
		_w10390_,
		_w10391_
	);
	LUT4 #(
		.INIT('h95aa)
	) name10358 (
		\a[8] ,
		_w4876_,
		_w7882_,
		_w10391_,
		_w10392_
	);
	LUT2 #(
		.INIT('h9)
	) name10359 (
		_w10217_,
		_w10219_,
		_w10393_
	);
	LUT2 #(
		.INIT('h4)
	) name10360 (
		_w10392_,
		_w10393_,
		_w10394_
	);
	LUT3 #(
		.INIT('h1e)
	) name10361 (
		_w10119_,
		_w10215_,
		_w10216_,
		_w10395_
	);
	LUT3 #(
		.INIT('h82)
	) name10362 (
		_w4876_,
		_w7093_,
		_w7095_,
		_w10396_
	);
	LUT3 #(
		.INIT('h82)
	) name10363 (
		_w5286_,
		_w6947_,
		_w6949_,
		_w10397_
	);
	LUT2 #(
		.INIT('h8)
	) name10364 (
		_w4875_,
		_w7038_,
		_w10398_
	);
	LUT4 #(
		.INIT('h04c8)
	) name10365 (
		_w4695_,
		_w5271_,
		_w6944_,
		_w6946_,
		_w10399_
	);
	LUT2 #(
		.INIT('h1)
	) name10366 (
		_w10398_,
		_w10399_,
		_w10400_
	);
	LUT2 #(
		.INIT('h4)
	) name10367 (
		_w10397_,
		_w10400_,
		_w10401_
	);
	LUT4 #(
		.INIT('h4844)
	) name10368 (
		\a[8] ,
		_w10395_,
		_w10396_,
		_w10401_,
		_w10402_
	);
	LUT4 #(
		.INIT('h54ab)
	) name10369 (
		_w10125_,
		_w10211_,
		_w10212_,
		_w10214_,
		_w10403_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10370 (
		_w4876_,
		_w7040_,
		_w7091_,
		_w7092_,
		_w10404_
	);
	LUT4 #(
		.INIT('h04c8)
	) name10371 (
		_w4695_,
		_w5286_,
		_w6944_,
		_w6946_,
		_w10405_
	);
	LUT3 #(
		.INIT('h82)
	) name10372 (
		_w4875_,
		_w6940_,
		_w6942_,
		_w10406_
	);
	LUT3 #(
		.INIT('h07)
	) name10373 (
		_w5271_,
		_w7038_,
		_w10406_,
		_w10407_
	);
	LUT2 #(
		.INIT('h4)
	) name10374 (
		_w10405_,
		_w10407_,
		_w10408_
	);
	LUT4 #(
		.INIT('h4844)
	) name10375 (
		\a[8] ,
		_w10403_,
		_w10404_,
		_w10408_,
		_w10409_
	);
	LUT2 #(
		.INIT('h9)
	) name10376 (
		_w10211_,
		_w10213_,
		_w10410_
	);
	LUT4 #(
		.INIT('h2228)
	) name10377 (
		_w4875_,
		_w5067_,
		_w5282_,
		_w6939_,
		_w10411_
	);
	LUT4 #(
		.INIT('h007d)
	) name10378 (
		_w5271_,
		_w6940_,
		_w6942_,
		_w10411_,
		_w10412_
	);
	LUT3 #(
		.INIT('h70)
	) name10379 (
		_w5286_,
		_w7038_,
		_w10412_,
		_w10413_
	);
	LUT4 #(
		.INIT('h95aa)
	) name10380 (
		\a[8] ,
		_w4876_,
		_w8018_,
		_w10413_,
		_w10414_
	);
	LUT2 #(
		.INIT('h2)
	) name10381 (
		_w10410_,
		_w10414_,
		_w10415_
	);
	LUT3 #(
		.INIT('h82)
	) name10382 (
		_w4876_,
		_w7087_,
		_w7089_,
		_w10416_
	);
	LUT3 #(
		.INIT('h82)
	) name10383 (
		_w5286_,
		_w6940_,
		_w6942_,
		_w10417_
	);
	LUT2 #(
		.INIT('h8)
	) name10384 (
		_w4875_,
		_w7044_,
		_w10418_
	);
	LUT4 #(
		.INIT('h4448)
	) name10385 (
		_w5067_,
		_w5271_,
		_w5282_,
		_w6939_,
		_w10419_
	);
	LUT2 #(
		.INIT('h1)
	) name10386 (
		_w10418_,
		_w10419_,
		_w10420_
	);
	LUT2 #(
		.INIT('h4)
	) name10387 (
		_w10417_,
		_w10420_,
		_w10421_
	);
	LUT3 #(
		.INIT('h1e)
	) name10388 (
		_w10140_,
		_w10209_,
		_w10210_,
		_w10422_
	);
	LUT4 #(
		.INIT('h6500)
	) name10389 (
		\a[8] ,
		_w10416_,
		_w10421_,
		_w10422_,
		_w10423_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10390 (
		_w4876_,
		_w7046_,
		_w7085_,
		_w7086_,
		_w10424_
	);
	LUT4 #(
		.INIT('h5060)
	) name10391 (
		_w5067_,
		_w5282_,
		_w5286_,
		_w6939_,
		_w10425_
	);
	LUT3 #(
		.INIT('h82)
	) name10392 (
		_w4875_,
		_w6935_,
		_w6937_,
		_w10426_
	);
	LUT3 #(
		.INIT('h07)
	) name10393 (
		_w5271_,
		_w7044_,
		_w10426_,
		_w10427_
	);
	LUT2 #(
		.INIT('h4)
	) name10394 (
		_w10425_,
		_w10427_,
		_w10428_
	);
	LUT4 #(
		.INIT('h54ab)
	) name10395 (
		_w10146_,
		_w10205_,
		_w10206_,
		_w10208_,
		_w10429_
	);
	LUT4 #(
		.INIT('h6500)
	) name10396 (
		\a[8] ,
		_w10424_,
		_w10428_,
		_w10429_,
		_w10430_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10397 (
		_w4875_,
		_w6043_,
		_w6933_,
		_w6934_,
		_w10431_
	);
	LUT4 #(
		.INIT('h007d)
	) name10398 (
		_w5271_,
		_w6935_,
		_w6937_,
		_w10431_,
		_w10432_
	);
	LUT3 #(
		.INIT('h70)
	) name10399 (
		_w5286_,
		_w7044_,
		_w10432_,
		_w10433_
	);
	LUT4 #(
		.INIT('h95aa)
	) name10400 (
		\a[8] ,
		_w4876_,
		_w8005_,
		_w10433_,
		_w10434_
	);
	LUT2 #(
		.INIT('h9)
	) name10401 (
		_w10205_,
		_w10207_,
		_w10435_
	);
	LUT2 #(
		.INIT('h4)
	) name10402 (
		_w10434_,
		_w10435_,
		_w10436_
	);
	LUT3 #(
		.INIT('h1e)
	) name10403 (
		_w10161_,
		_w10203_,
		_w10204_,
		_w10437_
	);
	LUT3 #(
		.INIT('h82)
	) name10404 (
		_w4876_,
		_w7081_,
		_w7083_,
		_w10438_
	);
	LUT3 #(
		.INIT('h82)
	) name10405 (
		_w5286_,
		_w6935_,
		_w6937_,
		_w10439_
	);
	LUT2 #(
		.INIT('h8)
	) name10406 (
		_w4875_,
		_w7050_,
		_w10440_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10407 (
		_w5271_,
		_w6043_,
		_w6933_,
		_w6934_,
		_w10441_
	);
	LUT2 #(
		.INIT('h1)
	) name10408 (
		_w10440_,
		_w10441_,
		_w10442_
	);
	LUT2 #(
		.INIT('h4)
	) name10409 (
		_w10439_,
		_w10442_,
		_w10443_
	);
	LUT4 #(
		.INIT('h4844)
	) name10410 (
		\a[8] ,
		_w10437_,
		_w10438_,
		_w10443_,
		_w10444_
	);
	LUT4 #(
		.INIT('h54ab)
	) name10411 (
		_w10168_,
		_w10199_,
		_w10200_,
		_w10202_,
		_w10445_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10412 (
		_w4876_,
		_w7052_,
		_w7079_,
		_w7080_,
		_w10446_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10413 (
		_w5286_,
		_w6043_,
		_w6933_,
		_w6934_,
		_w10447_
	);
	LUT3 #(
		.INIT('h82)
	) name10414 (
		_w4875_,
		_w6929_,
		_w6931_,
		_w10448_
	);
	LUT3 #(
		.INIT('h07)
	) name10415 (
		_w5271_,
		_w7050_,
		_w10448_,
		_w10449_
	);
	LUT2 #(
		.INIT('h4)
	) name10416 (
		_w10447_,
		_w10449_,
		_w10450_
	);
	LUT4 #(
		.INIT('h4844)
	) name10417 (
		\a[8] ,
		_w10445_,
		_w10446_,
		_w10450_,
		_w10451_
	);
	LUT2 #(
		.INIT('h9)
	) name10418 (
		_w10199_,
		_w10201_,
		_w10452_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10419 (
		_w4875_,
		_w6645_,
		_w6926_,
		_w6928_,
		_w10453_
	);
	LUT4 #(
		.INIT('h007d)
	) name10420 (
		_w5271_,
		_w6929_,
		_w6931_,
		_w10453_,
		_w10454_
	);
	LUT3 #(
		.INIT('h70)
	) name10421 (
		_w5286_,
		_w7050_,
		_w10454_,
		_w10455_
	);
	LUT4 #(
		.INIT('h95aa)
	) name10422 (
		\a[8] ,
		_w4876_,
		_w8227_,
		_w10455_,
		_w10456_
	);
	LUT2 #(
		.INIT('h2)
	) name10423 (
		_w10452_,
		_w10456_,
		_w10457_
	);
	LUT3 #(
		.INIT('h82)
	) name10424 (
		_w4876_,
		_w7075_,
		_w7077_,
		_w10458_
	);
	LUT3 #(
		.INIT('h82)
	) name10425 (
		_w5286_,
		_w6929_,
		_w6931_,
		_w10459_
	);
	LUT2 #(
		.INIT('h8)
	) name10426 (
		_w4875_,
		_w7056_,
		_w10460_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10427 (
		_w5271_,
		_w6645_,
		_w6926_,
		_w6928_,
		_w10461_
	);
	LUT2 #(
		.INIT('h1)
	) name10428 (
		_w10460_,
		_w10461_,
		_w10462_
	);
	LUT2 #(
		.INIT('h4)
	) name10429 (
		_w10459_,
		_w10462_,
		_w10463_
	);
	LUT2 #(
		.INIT('h9)
	) name10430 (
		_w10196_,
		_w10198_,
		_w10464_
	);
	LUT4 #(
		.INIT('h6500)
	) name10431 (
		\a[8] ,
		_w10458_,
		_w10463_,
		_w10464_,
		_w10465_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10432 (
		_w4876_,
		_w7058_,
		_w7073_,
		_w7074_,
		_w10466_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10433 (
		_w5286_,
		_w6645_,
		_w6926_,
		_w6928_,
		_w10467_
	);
	LUT3 #(
		.INIT('h82)
	) name10434 (
		_w4875_,
		_w6922_,
		_w6924_,
		_w10468_
	);
	LUT3 #(
		.INIT('h07)
	) name10435 (
		_w5271_,
		_w7056_,
		_w10468_,
		_w10469_
	);
	LUT2 #(
		.INIT('h4)
	) name10436 (
		_w10467_,
		_w10469_,
		_w10470_
	);
	LUT4 #(
		.INIT('h9a65)
	) name10437 (
		\a[11] ,
		_w10189_,
		_w10193_,
		_w10194_,
		_w10471_
	);
	LUT4 #(
		.INIT('h6500)
	) name10438 (
		\a[8] ,
		_w10466_,
		_w10470_,
		_w10471_,
		_w10472_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10439 (
		_w4875_,
		_w6669_,
		_w6919_,
		_w6921_,
		_w10473_
	);
	LUT4 #(
		.INIT('h007d)
	) name10440 (
		_w5271_,
		_w6922_,
		_w6924_,
		_w10473_,
		_w10474_
	);
	LUT3 #(
		.INIT('h70)
	) name10441 (
		_w5286_,
		_w7056_,
		_w10474_,
		_w10475_
	);
	LUT4 #(
		.INIT('h95aa)
	) name10442 (
		\a[8] ,
		_w4876_,
		_w8298_,
		_w10475_,
		_w10476_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name10443 (
		\a[11] ,
		_w10181_,
		_w10178_,
		_w10180_,
		_w10477_
	);
	LUT3 #(
		.INIT('h4b)
	) name10444 (
		_w10184_,
		_w10187_,
		_w10477_,
		_w10478_
	);
	LUT2 #(
		.INIT('h4)
	) name10445 (
		_w10476_,
		_w10478_,
		_w10479_
	);
	LUT3 #(
		.INIT('h82)
	) name10446 (
		_w4876_,
		_w7069_,
		_w7071_,
		_w10480_
	);
	LUT3 #(
		.INIT('h82)
	) name10447 (
		_w5286_,
		_w6922_,
		_w6924_,
		_w10481_
	);
	LUT2 #(
		.INIT('h8)
	) name10448 (
		_w4875_,
		_w7062_,
		_w10482_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10449 (
		_w5271_,
		_w6669_,
		_w6919_,
		_w6921_,
		_w10483_
	);
	LUT2 #(
		.INIT('h1)
	) name10450 (
		_w10482_,
		_w10483_,
		_w10484_
	);
	LUT2 #(
		.INIT('h4)
	) name10451 (
		_w10481_,
		_w10484_,
		_w10485_
	);
	LUT2 #(
		.INIT('h8)
	) name10452 (
		\a[11] ,
		_w10181_,
		_w10486_
	);
	LUT3 #(
		.INIT('h4b)
	) name10453 (
		_w10178_,
		_w10180_,
		_w10486_,
		_w10487_
	);
	LUT4 #(
		.INIT('h6500)
	) name10454 (
		\a[8] ,
		_w10480_,
		_w10485_,
		_w10487_,
		_w10488_
	);
	LUT4 #(
		.INIT('h2882)
	) name10455 (
		_w4876_,
		_w6914_,
		_w6916_,
		_w7067_,
		_w10489_
	);
	LUT4 #(
		.INIT('ha802)
	) name10456 (
		_w5271_,
		_w6689_,
		_w6911_,
		_w6913_,
		_w10490_
	);
	LUT4 #(
		.INIT('h007d)
	) name10457 (
		_w5286_,
		_w6914_,
		_w6916_,
		_w10490_,
		_w10491_
	);
	LUT4 #(
		.INIT('h5401)
	) name10458 (
		_w4874_,
		_w6689_,
		_w6911_,
		_w6913_,
		_w10492_
	);
	LUT2 #(
		.INIT('h2)
	) name10459 (
		\a[8] ,
		_w10492_,
		_w10493_
	);
	LUT3 #(
		.INIT('h40)
	) name10460 (
		_w10489_,
		_w10491_,
		_w10493_,
		_w10494_
	);
	LUT3 #(
		.INIT('h28)
	) name10461 (
		_w4876_,
		_w7062_,
		_w8358_,
		_w10495_
	);
	LUT4 #(
		.INIT('ha802)
	) name10462 (
		_w4875_,
		_w6689_,
		_w6911_,
		_w6913_,
		_w10496_
	);
	LUT4 #(
		.INIT('h007d)
	) name10463 (
		_w5271_,
		_w6914_,
		_w6916_,
		_w10496_,
		_w10497_
	);
	LUT3 #(
		.INIT('h70)
	) name10464 (
		_w5286_,
		_w7062_,
		_w10497_,
		_w10498_
	);
	LUT4 #(
		.INIT('h0800)
	) name10465 (
		_w10181_,
		_w10494_,
		_w10495_,
		_w10498_,
		_w10499_
	);
	LUT3 #(
		.INIT('h28)
	) name10466 (
		_w4876_,
		_w7065_,
		_w7068_,
		_w10500_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10467 (
		_w5286_,
		_w6669_,
		_w6919_,
		_w6921_,
		_w10501_
	);
	LUT3 #(
		.INIT('h82)
	) name10468 (
		_w4875_,
		_w6914_,
		_w6916_,
		_w10502_
	);
	LUT3 #(
		.INIT('h07)
	) name10469 (
		_w5271_,
		_w7062_,
		_w10502_,
		_w10503_
	);
	LUT2 #(
		.INIT('h4)
	) name10470 (
		_w10501_,
		_w10503_,
		_w10504_
	);
	LUT4 #(
		.INIT('ha6aa)
	) name10471 (
		_w10181_,
		_w10494_,
		_w10495_,
		_w10498_,
		_w10505_
	);
	LUT4 #(
		.INIT('h6500)
	) name10472 (
		\a[8] ,
		_w10500_,
		_w10504_,
		_w10505_,
		_w10506_
	);
	LUT2 #(
		.INIT('h1)
	) name10473 (
		_w10499_,
		_w10506_,
		_w10507_
	);
	LUT4 #(
		.INIT('h009a)
	) name10474 (
		\a[8] ,
		_w10480_,
		_w10485_,
		_w10487_,
		_w10508_
	);
	LUT4 #(
		.INIT('h9a65)
	) name10475 (
		\a[8] ,
		_w10480_,
		_w10485_,
		_w10487_,
		_w10509_
	);
	LUT3 #(
		.INIT('h54)
	) name10476 (
		_w10488_,
		_w10507_,
		_w10508_,
		_w10510_
	);
	LUT2 #(
		.INIT('h2)
	) name10477 (
		_w10476_,
		_w10478_,
		_w10511_
	);
	LUT2 #(
		.INIT('h9)
	) name10478 (
		_w10476_,
		_w10478_,
		_w10512_
	);
	LUT4 #(
		.INIT('h9a65)
	) name10479 (
		\a[8] ,
		_w10466_,
		_w10470_,
		_w10471_,
		_w10513_
	);
	LUT4 #(
		.INIT('h4d00)
	) name10480 (
		_w10476_,
		_w10478_,
		_w10510_,
		_w10513_,
		_w10514_
	);
	LUT4 #(
		.INIT('h9a65)
	) name10481 (
		\a[8] ,
		_w10458_,
		_w10463_,
		_w10464_,
		_w10515_
	);
	LUT4 #(
		.INIT('h0155)
	) name10482 (
		_w10465_,
		_w10472_,
		_w10514_,
		_w10515_,
		_w10516_
	);
	LUT2 #(
		.INIT('h4)
	) name10483 (
		_w10452_,
		_w10456_,
		_w10517_
	);
	LUT2 #(
		.INIT('h9)
	) name10484 (
		_w10452_,
		_w10456_,
		_w10518_
	);
	LUT4 #(
		.INIT('h9699)
	) name10485 (
		\a[8] ,
		_w10445_,
		_w10446_,
		_w10450_,
		_w10519_
	);
	LUT4 #(
		.INIT('h2b00)
	) name10486 (
		_w10452_,
		_w10456_,
		_w10516_,
		_w10519_,
		_w10520_
	);
	LUT4 #(
		.INIT('h9699)
	) name10487 (
		\a[8] ,
		_w10437_,
		_w10438_,
		_w10443_,
		_w10521_
	);
	LUT4 #(
		.INIT('h0155)
	) name10488 (
		_w10444_,
		_w10451_,
		_w10520_,
		_w10521_,
		_w10522_
	);
	LUT2 #(
		.INIT('h2)
	) name10489 (
		_w10434_,
		_w10435_,
		_w10523_
	);
	LUT2 #(
		.INIT('h9)
	) name10490 (
		_w10434_,
		_w10435_,
		_w10524_
	);
	LUT4 #(
		.INIT('h9a65)
	) name10491 (
		\a[8] ,
		_w10424_,
		_w10428_,
		_w10429_,
		_w10525_
	);
	LUT4 #(
		.INIT('h4d00)
	) name10492 (
		_w10434_,
		_w10435_,
		_w10522_,
		_w10525_,
		_w10526_
	);
	LUT4 #(
		.INIT('h9a65)
	) name10493 (
		\a[8] ,
		_w10416_,
		_w10421_,
		_w10422_,
		_w10527_
	);
	LUT4 #(
		.INIT('h0155)
	) name10494 (
		_w10423_,
		_w10430_,
		_w10526_,
		_w10527_,
		_w10528_
	);
	LUT2 #(
		.INIT('h4)
	) name10495 (
		_w10410_,
		_w10414_,
		_w10529_
	);
	LUT2 #(
		.INIT('h9)
	) name10496 (
		_w10410_,
		_w10414_,
		_w10530_
	);
	LUT4 #(
		.INIT('h9699)
	) name10497 (
		\a[8] ,
		_w10403_,
		_w10404_,
		_w10408_,
		_w10531_
	);
	LUT4 #(
		.INIT('h2b00)
	) name10498 (
		_w10410_,
		_w10414_,
		_w10528_,
		_w10531_,
		_w10532_
	);
	LUT4 #(
		.INIT('h9699)
	) name10499 (
		\a[8] ,
		_w10395_,
		_w10396_,
		_w10401_,
		_w10533_
	);
	LUT4 #(
		.INIT('h0155)
	) name10500 (
		_w10402_,
		_w10409_,
		_w10532_,
		_w10533_,
		_w10534_
	);
	LUT2 #(
		.INIT('h2)
	) name10501 (
		_w10392_,
		_w10393_,
		_w10535_
	);
	LUT2 #(
		.INIT('h9)
	) name10502 (
		_w10392_,
		_w10393_,
		_w10536_
	);
	LUT4 #(
		.INIT('h9a65)
	) name10503 (
		\a[8] ,
		_w10382_,
		_w10386_,
		_w10387_,
		_w10537_
	);
	LUT4 #(
		.INIT('h4d00)
	) name10504 (
		_w10392_,
		_w10393_,
		_w10534_,
		_w10537_,
		_w10538_
	);
	LUT4 #(
		.INIT('h9a65)
	) name10505 (
		\a[8] ,
		_w10374_,
		_w10379_,
		_w10380_,
		_w10539_
	);
	LUT4 #(
		.INIT('h0155)
	) name10506 (
		_w10381_,
		_w10388_,
		_w10538_,
		_w10539_,
		_w10540_
	);
	LUT2 #(
		.INIT('h4)
	) name10507 (
		_w10368_,
		_w10372_,
		_w10541_
	);
	LUT2 #(
		.INIT('h9)
	) name10508 (
		_w10368_,
		_w10372_,
		_w10542_
	);
	LUT4 #(
		.INIT('h9699)
	) name10509 (
		\a[8] ,
		_w10361_,
		_w10362_,
		_w10366_,
		_w10543_
	);
	LUT4 #(
		.INIT('h2b00)
	) name10510 (
		_w10368_,
		_w10372_,
		_w10540_,
		_w10543_,
		_w10544_
	);
	LUT4 #(
		.INIT('h9699)
	) name10511 (
		\a[8] ,
		_w10353_,
		_w10354_,
		_w10359_,
		_w10545_
	);
	LUT4 #(
		.INIT('h0155)
	) name10512 (
		_w10360_,
		_w10367_,
		_w10544_,
		_w10545_,
		_w10546_
	);
	LUT2 #(
		.INIT('h2)
	) name10513 (
		_w10350_,
		_w10351_,
		_w10547_
	);
	LUT2 #(
		.INIT('h9)
	) name10514 (
		_w10350_,
		_w10351_,
		_w10548_
	);
	LUT4 #(
		.INIT('h9a65)
	) name10515 (
		\a[8] ,
		_w10340_,
		_w10344_,
		_w10345_,
		_w10549_
	);
	LUT4 #(
		.INIT('h4d00)
	) name10516 (
		_w10350_,
		_w10351_,
		_w10546_,
		_w10549_,
		_w10550_
	);
	LUT4 #(
		.INIT('h9699)
	) name10517 (
		\a[8] ,
		_w10332_,
		_w10333_,
		_w10338_,
		_w10551_
	);
	LUT4 #(
		.INIT('h0155)
	) name10518 (
		_w10339_,
		_w10346_,
		_w10550_,
		_w10551_,
		_w10552_
	);
	LUT2 #(
		.INIT('h4)
	) name10519 (
		_w10326_,
		_w10330_,
		_w10553_
	);
	LUT2 #(
		.INIT('h9)
	) name10520 (
		_w10326_,
		_w10330_,
		_w10554_
	);
	LUT4 #(
		.INIT('h9699)
	) name10521 (
		\a[8] ,
		_w10319_,
		_w10320_,
		_w10324_,
		_w10555_
	);
	LUT4 #(
		.INIT('h2b00)
	) name10522 (
		_w10326_,
		_w10330_,
		_w10552_,
		_w10555_,
		_w10556_
	);
	LUT4 #(
		.INIT('h9699)
	) name10523 (
		\a[8] ,
		_w10311_,
		_w10312_,
		_w10317_,
		_w10557_
	);
	LUT4 #(
		.INIT('h0155)
	) name10524 (
		_w10318_,
		_w10325_,
		_w10556_,
		_w10557_,
		_w10558_
	);
	LUT2 #(
		.INIT('h4)
	) name10525 (
		_w10305_,
		_w10309_,
		_w10559_
	);
	LUT2 #(
		.INIT('h9)
	) name10526 (
		_w10305_,
		_w10309_,
		_w10560_
	);
	LUT4 #(
		.INIT('h9699)
	) name10527 (
		\a[8] ,
		_w10298_,
		_w10299_,
		_w10303_,
		_w10561_
	);
	LUT4 #(
		.INIT('h2b00)
	) name10528 (
		_w10305_,
		_w10309_,
		_w10558_,
		_w10561_,
		_w10562_
	);
	LUT4 #(
		.INIT('h9699)
	) name10529 (
		\a[8] ,
		_w10290_,
		_w10291_,
		_w10296_,
		_w10563_
	);
	LUT4 #(
		.INIT('h0155)
	) name10530 (
		_w10297_,
		_w10304_,
		_w10562_,
		_w10563_,
		_w10564_
	);
	LUT2 #(
		.INIT('h4)
	) name10531 (
		_w10284_,
		_w10288_,
		_w10565_
	);
	LUT2 #(
		.INIT('h9)
	) name10532 (
		_w10284_,
		_w10288_,
		_w10566_
	);
	LUT4 #(
		.INIT('h9699)
	) name10533 (
		\a[8] ,
		_w10277_,
		_w10278_,
		_w10282_,
		_w10567_
	);
	LUT4 #(
		.INIT('h2b00)
	) name10534 (
		_w10284_,
		_w10288_,
		_w10564_,
		_w10567_,
		_w10568_
	);
	LUT4 #(
		.INIT('h9699)
	) name10535 (
		\a[8] ,
		_w10269_,
		_w10270_,
		_w10275_,
		_w10569_
	);
	LUT4 #(
		.INIT('h0155)
	) name10536 (
		_w10276_,
		_w10283_,
		_w10568_,
		_w10569_,
		_w10570_
	);
	LUT4 #(
		.INIT('h9669)
	) name10537 (
		_w9963_,
		_w10253_,
		_w10254_,
		_w10258_,
		_w10571_
	);
	LUT3 #(
		.INIT('h28)
	) name10538 (
		_w6031_,
		_w7136_,
		_w7168_,
		_w10572_
	);
	LUT4 #(
		.INIT('h028a)
	) name10539 (
		_w6324_,
		_w7136_,
		_w7166_,
		_w7167_,
		_w10573_
	);
	LUT4 #(
		.INIT('h04c8)
	) name10540 (
		_w2411_,
		_w5524_,
		_w6983_,
		_w6993_,
		_w10574_
	);
	LUT3 #(
		.INIT('h01)
	) name10541 (
		_w10573_,
		_w10574_,
		_w10572_,
		_w10575_
	);
	LUT4 #(
		.INIT('h95aa)
	) name10542 (
		\a[5] ,
		_w35_,
		_w7696_,
		_w10575_,
		_w10576_
	);
	LUT3 #(
		.INIT('hb2)
	) name10543 (
		_w10570_,
		_w10571_,
		_w10576_,
		_w10577_
	);
	LUT4 #(
		.INIT('h0096)
	) name10544 (
		_w9978_,
		_w10259_,
		_w10264_,
		_w10577_,
		_w10578_
	);
	LUT4 #(
		.INIT('h6900)
	) name10545 (
		_w9978_,
		_w10259_,
		_w10264_,
		_w10577_,
		_w10579_
	);
	LUT4 #(
		.INIT('h9669)
	) name10546 (
		_w9978_,
		_w10259_,
		_w10264_,
		_w10577_,
		_w10580_
	);
	LUT3 #(
		.INIT('h82)
	) name10547 (
		_w35_,
		_w7135_,
		_w7172_,
		_w10581_
	);
	LUT3 #(
		.INIT('h28)
	) name10548 (
		_w6324_,
		_w7136_,
		_w7168_,
		_w10582_
	);
	LUT2 #(
		.INIT('h8)
	) name10549 (
		_w5524_,
		_w6996_,
		_w10583_
	);
	LUT4 #(
		.INIT('h04c8)
	) name10550 (
		_w2411_,
		_w6031_,
		_w6983_,
		_w6993_,
		_w10584_
	);
	LUT2 #(
		.INIT('h1)
	) name10551 (
		_w10583_,
		_w10584_,
		_w10585_
	);
	LUT2 #(
		.INIT('h4)
	) name10552 (
		_w10582_,
		_w10585_,
		_w10586_
	);
	LUT3 #(
		.INIT('h1e)
	) name10553 (
		_w10283_,
		_w10568_,
		_w10569_,
		_w10587_
	);
	LUT4 #(
		.INIT('h6500)
	) name10554 (
		\a[5] ,
		_w10581_,
		_w10586_,
		_w10587_,
		_w10588_
	);
	LUT4 #(
		.INIT('h028a)
	) name10555 (
		_w6334_,
		_w7136_,
		_w7166_,
		_w7167_,
		_w10589_
	);
	LUT3 #(
		.INIT('hc6)
	) name10556 (
		\a[0] ,
		\a[1] ,
		\a[2] ,
		_w10590_
	);
	LUT3 #(
		.INIT('hb0)
	) name10557 (
		_w7136_,
		_w7166_,
		_w10590_,
		_w10591_
	);
	LUT2 #(
		.INIT('h1)
	) name10558 (
		_w10589_,
		_w10591_,
		_w10592_
	);
	LUT4 #(
		.INIT('h5700)
	) name10559 (
		_w6335_,
		_w7418_,
		_w7419_,
		_w10592_,
		_w10593_
	);
	LUT4 #(
		.INIT('h009a)
	) name10560 (
		\a[5] ,
		_w10581_,
		_w10586_,
		_w10587_,
		_w10594_
	);
	LUT4 #(
		.INIT('h9a65)
	) name10561 (
		\a[5] ,
		_w10581_,
		_w10586_,
		_w10587_,
		_w10595_
	);
	LUT4 #(
		.INIT('h3312)
	) name10562 (
		\a[2] ,
		_w10588_,
		_w10593_,
		_w10594_,
		_w10596_
	);
	LUT4 #(
		.INIT('h0096)
	) name10563 (
		_w10570_,
		_w10571_,
		_w10576_,
		_w10596_,
		_w10597_
	);
	LUT4 #(
		.INIT('h6900)
	) name10564 (
		_w10570_,
		_w10571_,
		_w10576_,
		_w10596_,
		_w10598_
	);
	LUT4 #(
		.INIT('h9669)
	) name10565 (
		_w10570_,
		_w10571_,
		_w10576_,
		_w10596_,
		_w10599_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10566 (
		_w35_,
		_w6998_,
		_w7133_,
		_w7134_,
		_w10600_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10567 (
		_w6324_,
		_w2411_,
		_w6983_,
		_w6993_,
		_w10601_
	);
	LUT3 #(
		.INIT('h84)
	) name10568 (
		_w2546_,
		_w5524_,
		_w6981_,
		_w10602_
	);
	LUT3 #(
		.INIT('h07)
	) name10569 (
		_w6031_,
		_w6996_,
		_w10602_,
		_w10603_
	);
	LUT2 #(
		.INIT('h4)
	) name10570 (
		_w10601_,
		_w10603_,
		_w10604_
	);
	LUT4 #(
		.INIT('h54ab)
	) name10571 (
		_w10289_,
		_w10564_,
		_w10565_,
		_w10567_,
		_w10605_
	);
	LUT4 #(
		.INIT('h6500)
	) name10572 (
		\a[5] ,
		_w10600_,
		_w10604_,
		_w10605_,
		_w10606_
	);
	LUT4 #(
		.INIT('h04c8)
	) name10573 (
		_w2622_,
		_w5524_,
		_w6978_,
		_w6980_,
		_w10607_
	);
	LUT4 #(
		.INIT('h007b)
	) name10574 (
		_w2546_,
		_w6031_,
		_w6981_,
		_w10607_,
		_w10608_
	);
	LUT3 #(
		.INIT('h70)
	) name10575 (
		_w6324_,
		_w6996_,
		_w10608_,
		_w10609_
	);
	LUT4 #(
		.INIT('h95aa)
	) name10576 (
		\a[5] ,
		_w35_,
		_w7500_,
		_w10609_,
		_w10610_
	);
	LUT2 #(
		.INIT('h9)
	) name10577 (
		_w10564_,
		_w10566_,
		_w10611_
	);
	LUT2 #(
		.INIT('h4)
	) name10578 (
		_w10610_,
		_w10611_,
		_w10612_
	);
	LUT3 #(
		.INIT('h82)
	) name10579 (
		_w35_,
		_w7129_,
		_w7131_,
		_w10613_
	);
	LUT3 #(
		.INIT('h82)
	) name10580 (
		_w6324_,
		_w2546_,
		_w6981_,
		_w10614_
	);
	LUT2 #(
		.INIT('h8)
	) name10581 (
		_w5524_,
		_w7002_,
		_w10615_
	);
	LUT4 #(
		.INIT('h04c8)
	) name10582 (
		_w2622_,
		_w6031_,
		_w6978_,
		_w6980_,
		_w10616_
	);
	LUT2 #(
		.INIT('h1)
	) name10583 (
		_w10615_,
		_w10616_,
		_w10617_
	);
	LUT2 #(
		.INIT('h4)
	) name10584 (
		_w10614_,
		_w10617_,
		_w10618_
	);
	LUT3 #(
		.INIT('h1e)
	) name10585 (
		_w10304_,
		_w10562_,
		_w10563_,
		_w10619_
	);
	LUT4 #(
		.INIT('h6500)
	) name10586 (
		\a[5] ,
		_w10613_,
		_w10618_,
		_w10619_,
		_w10620_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10587 (
		_w35_,
		_w7004_,
		_w7127_,
		_w7128_,
		_w10621_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10588 (
		_w6324_,
		_w2622_,
		_w6978_,
		_w6980_,
		_w10622_
	);
	LUT3 #(
		.INIT('h84)
	) name10589 (
		_w2872_,
		_w5524_,
		_w6975_,
		_w10623_
	);
	LUT3 #(
		.INIT('h07)
	) name10590 (
		_w6031_,
		_w7002_,
		_w10623_,
		_w10624_
	);
	LUT2 #(
		.INIT('h4)
	) name10591 (
		_w10622_,
		_w10624_,
		_w10625_
	);
	LUT4 #(
		.INIT('h54ab)
	) name10592 (
		_w10310_,
		_w10558_,
		_w10559_,
		_w10561_,
		_w10626_
	);
	LUT4 #(
		.INIT('h6500)
	) name10593 (
		\a[5] ,
		_w10621_,
		_w10625_,
		_w10626_,
		_w10627_
	);
	LUT4 #(
		.INIT('h04c8)
	) name10594 (
		_w2983_,
		_w5524_,
		_w6972_,
		_w6974_,
		_w10628_
	);
	LUT4 #(
		.INIT('h007b)
	) name10595 (
		_w2872_,
		_w6031_,
		_w6975_,
		_w10628_,
		_w10629_
	);
	LUT3 #(
		.INIT('h70)
	) name10596 (
		_w6324_,
		_w7002_,
		_w10629_,
		_w10630_
	);
	LUT4 #(
		.INIT('h95aa)
	) name10597 (
		\a[5] ,
		_w35_,
		_w7426_,
		_w10630_,
		_w10631_
	);
	LUT2 #(
		.INIT('h9)
	) name10598 (
		_w10558_,
		_w10560_,
		_w10632_
	);
	LUT2 #(
		.INIT('h4)
	) name10599 (
		_w10631_,
		_w10632_,
		_w10633_
	);
	LUT3 #(
		.INIT('h82)
	) name10600 (
		_w35_,
		_w7123_,
		_w7125_,
		_w10634_
	);
	LUT3 #(
		.INIT('h82)
	) name10601 (
		_w6324_,
		_w2872_,
		_w6975_,
		_w10635_
	);
	LUT2 #(
		.INIT('h8)
	) name10602 (
		_w5524_,
		_w7008_,
		_w10636_
	);
	LUT4 #(
		.INIT('h04c8)
	) name10603 (
		_w2983_,
		_w6031_,
		_w6972_,
		_w6974_,
		_w10637_
	);
	LUT2 #(
		.INIT('h1)
	) name10604 (
		_w10636_,
		_w10637_,
		_w10638_
	);
	LUT2 #(
		.INIT('h4)
	) name10605 (
		_w10635_,
		_w10638_,
		_w10639_
	);
	LUT3 #(
		.INIT('h1e)
	) name10606 (
		_w10325_,
		_w10556_,
		_w10557_,
		_w10640_
	);
	LUT4 #(
		.INIT('h6500)
	) name10607 (
		\a[5] ,
		_w10634_,
		_w10639_,
		_w10640_,
		_w10641_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10608 (
		_w35_,
		_w7010_,
		_w7121_,
		_w7122_,
		_w10642_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10609 (
		_w6324_,
		_w2983_,
		_w6972_,
		_w6974_,
		_w10643_
	);
	LUT3 #(
		.INIT('h82)
	) name10610 (
		_w5524_,
		_w6967_,
		_w6969_,
		_w10644_
	);
	LUT3 #(
		.INIT('h07)
	) name10611 (
		_w6031_,
		_w7008_,
		_w10644_,
		_w10645_
	);
	LUT2 #(
		.INIT('h4)
	) name10612 (
		_w10643_,
		_w10645_,
		_w10646_
	);
	LUT4 #(
		.INIT('h54ab)
	) name10613 (
		_w10331_,
		_w10552_,
		_w10553_,
		_w10555_,
		_w10647_
	);
	LUT4 #(
		.INIT('h6500)
	) name10614 (
		\a[5] ,
		_w10642_,
		_w10646_,
		_w10647_,
		_w10648_
	);
	LUT4 #(
		.INIT('h04c8)
	) name10615 (
		_w3257_,
		_w5524_,
		_w6964_,
		_w6966_,
		_w10649_
	);
	LUT4 #(
		.INIT('h007d)
	) name10616 (
		_w6031_,
		_w6967_,
		_w6969_,
		_w10649_,
		_w10650_
	);
	LUT3 #(
		.INIT('h70)
	) name10617 (
		_w6324_,
		_w7008_,
		_w10650_,
		_w10651_
	);
	LUT4 #(
		.INIT('h95aa)
	) name10618 (
		\a[5] ,
		_w35_,
		_w7403_,
		_w10651_,
		_w10652_
	);
	LUT2 #(
		.INIT('h9)
	) name10619 (
		_w10552_,
		_w10554_,
		_w10653_
	);
	LUT2 #(
		.INIT('h4)
	) name10620 (
		_w10652_,
		_w10653_,
		_w10654_
	);
	LUT3 #(
		.INIT('h82)
	) name10621 (
		_w35_,
		_w7117_,
		_w7119_,
		_w10655_
	);
	LUT3 #(
		.INIT('h82)
	) name10622 (
		_w6324_,
		_w6967_,
		_w6969_,
		_w10656_
	);
	LUT2 #(
		.INIT('h8)
	) name10623 (
		_w5524_,
		_w7014_,
		_w10657_
	);
	LUT4 #(
		.INIT('h04c8)
	) name10624 (
		_w3257_,
		_w6031_,
		_w6964_,
		_w6966_,
		_w10658_
	);
	LUT2 #(
		.INIT('h1)
	) name10625 (
		_w10657_,
		_w10658_,
		_w10659_
	);
	LUT2 #(
		.INIT('h4)
	) name10626 (
		_w10656_,
		_w10659_,
		_w10660_
	);
	LUT3 #(
		.INIT('h1e)
	) name10627 (
		_w10346_,
		_w10550_,
		_w10551_,
		_w10661_
	);
	LUT4 #(
		.INIT('h6500)
	) name10628 (
		\a[5] ,
		_w10655_,
		_w10660_,
		_w10661_,
		_w10662_
	);
	LUT4 #(
		.INIT('h54ab)
	) name10629 (
		_w10352_,
		_w10546_,
		_w10547_,
		_w10549_,
		_w10663_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10630 (
		_w35_,
		_w7016_,
		_w7115_,
		_w7116_,
		_w10664_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10631 (
		_w6324_,
		_w3257_,
		_w6964_,
		_w6966_,
		_w10665_
	);
	LUT3 #(
		.INIT('h82)
	) name10632 (
		_w5524_,
		_w6960_,
		_w6962_,
		_w10666_
	);
	LUT3 #(
		.INIT('h07)
	) name10633 (
		_w6031_,
		_w7014_,
		_w10666_,
		_w10667_
	);
	LUT2 #(
		.INIT('h4)
	) name10634 (
		_w10665_,
		_w10667_,
		_w10668_
	);
	LUT4 #(
		.INIT('h4844)
	) name10635 (
		\a[5] ,
		_w10663_,
		_w10664_,
		_w10668_,
		_w10669_
	);
	LUT2 #(
		.INIT('h9)
	) name10636 (
		_w10546_,
		_w10548_,
		_w10670_
	);
	LUT4 #(
		.INIT('h5060)
	) name10637 (
		_w3409_,
		_w3650_,
		_w5524_,
		_w6959_,
		_w10671_
	);
	LUT4 #(
		.INIT('h007d)
	) name10638 (
		_w6031_,
		_w6960_,
		_w6962_,
		_w10671_,
		_w10672_
	);
	LUT3 #(
		.INIT('h70)
	) name10639 (
		_w6324_,
		_w7014_,
		_w10672_,
		_w10673_
	);
	LUT4 #(
		.INIT('h95aa)
	) name10640 (
		\a[5] ,
		_w35_,
		_w7291_,
		_w10673_,
		_w10674_
	);
	LUT2 #(
		.INIT('h2)
	) name10641 (
		_w10670_,
		_w10674_,
		_w10675_
	);
	LUT3 #(
		.INIT('h82)
	) name10642 (
		_w35_,
		_w7111_,
		_w7113_,
		_w10676_
	);
	LUT3 #(
		.INIT('h82)
	) name10643 (
		_w6324_,
		_w6960_,
		_w6962_,
		_w10677_
	);
	LUT2 #(
		.INIT('h8)
	) name10644 (
		_w5524_,
		_w7020_,
		_w10678_
	);
	LUT4 #(
		.INIT('h5060)
	) name10645 (
		_w3409_,
		_w3650_,
		_w6031_,
		_w6959_,
		_w10679_
	);
	LUT2 #(
		.INIT('h1)
	) name10646 (
		_w10678_,
		_w10679_,
		_w10680_
	);
	LUT2 #(
		.INIT('h4)
	) name10647 (
		_w10677_,
		_w10680_,
		_w10681_
	);
	LUT3 #(
		.INIT('h1e)
	) name10648 (
		_w10367_,
		_w10544_,
		_w10545_,
		_w10682_
	);
	LUT4 #(
		.INIT('h6500)
	) name10649 (
		\a[5] ,
		_w10676_,
		_w10681_,
		_w10682_,
		_w10683_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10650 (
		_w35_,
		_w7022_,
		_w7109_,
		_w7110_,
		_w10684_
	);
	LUT4 #(
		.INIT('h2228)
	) name10651 (
		_w6324_,
		_w3409_,
		_w3650_,
		_w6959_,
		_w10685_
	);
	LUT3 #(
		.INIT('h84)
	) name10652 (
		_w3706_,
		_w5524_,
		_w6957_,
		_w10686_
	);
	LUT3 #(
		.INIT('h07)
	) name10653 (
		_w6031_,
		_w7020_,
		_w10686_,
		_w10687_
	);
	LUT2 #(
		.INIT('h4)
	) name10654 (
		_w10685_,
		_w10687_,
		_w10688_
	);
	LUT4 #(
		.INIT('h54ab)
	) name10655 (
		_w10373_,
		_w10540_,
		_w10541_,
		_w10543_,
		_w10689_
	);
	LUT4 #(
		.INIT('h6500)
	) name10656 (
		\a[5] ,
		_w10684_,
		_w10688_,
		_w10689_,
		_w10690_
	);
	LUT4 #(
		.INIT('h04c8)
	) name10657 (
		_w3882_,
		_w5524_,
		_w6954_,
		_w6956_,
		_w10691_
	);
	LUT4 #(
		.INIT('h007b)
	) name10658 (
		_w3706_,
		_w6031_,
		_w6957_,
		_w10691_,
		_w10692_
	);
	LUT3 #(
		.INIT('h70)
	) name10659 (
		_w6324_,
		_w7020_,
		_w10692_,
		_w10693_
	);
	LUT4 #(
		.INIT('h95aa)
	) name10660 (
		\a[5] ,
		_w35_,
		_w7465_,
		_w10693_,
		_w10694_
	);
	LUT2 #(
		.INIT('h9)
	) name10661 (
		_w10540_,
		_w10542_,
		_w10695_
	);
	LUT2 #(
		.INIT('h4)
	) name10662 (
		_w10694_,
		_w10695_,
		_w10696_
	);
	LUT3 #(
		.INIT('h1e)
	) name10663 (
		_w10388_,
		_w10538_,
		_w10539_,
		_w10697_
	);
	LUT3 #(
		.INIT('h82)
	) name10664 (
		_w35_,
		_w7105_,
		_w7107_,
		_w10698_
	);
	LUT3 #(
		.INIT('h82)
	) name10665 (
		_w6324_,
		_w3706_,
		_w6957_,
		_w10699_
	);
	LUT2 #(
		.INIT('h8)
	) name10666 (
		_w5524_,
		_w7026_,
		_w10700_
	);
	LUT4 #(
		.INIT('h04c8)
	) name10667 (
		_w3882_,
		_w6031_,
		_w6954_,
		_w6956_,
		_w10701_
	);
	LUT2 #(
		.INIT('h1)
	) name10668 (
		_w10700_,
		_w10701_,
		_w10702_
	);
	LUT2 #(
		.INIT('h4)
	) name10669 (
		_w10699_,
		_w10702_,
		_w10703_
	);
	LUT4 #(
		.INIT('h4844)
	) name10670 (
		\a[5] ,
		_w10697_,
		_w10698_,
		_w10703_,
		_w10704_
	);
	LUT4 #(
		.INIT('h54ab)
	) name10671 (
		_w10394_,
		_w10534_,
		_w10535_,
		_w10537_,
		_w10705_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10672 (
		_w35_,
		_w7028_,
		_w7103_,
		_w7104_,
		_w10706_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10673 (
		_w6324_,
		_w3882_,
		_w6954_,
		_w6956_,
		_w10707_
	);
	LUT3 #(
		.INIT('h84)
	) name10674 (
		_w4030_,
		_w5524_,
		_w6952_,
		_w10708_
	);
	LUT3 #(
		.INIT('h07)
	) name10675 (
		_w6031_,
		_w7026_,
		_w10708_,
		_w10709_
	);
	LUT2 #(
		.INIT('h4)
	) name10676 (
		_w10707_,
		_w10709_,
		_w10710_
	);
	LUT4 #(
		.INIT('h4844)
	) name10677 (
		\a[5] ,
		_w10705_,
		_w10706_,
		_w10710_,
		_w10711_
	);
	LUT2 #(
		.INIT('h9)
	) name10678 (
		_w10534_,
		_w10536_,
		_w10712_
	);
	LUT4 #(
		.INIT('h5060)
	) name10679 (
		_w4099_,
		_w4378_,
		_w5524_,
		_w6951_,
		_w10713_
	);
	LUT4 #(
		.INIT('h007b)
	) name10680 (
		_w4030_,
		_w6031_,
		_w6952_,
		_w10713_,
		_w10714_
	);
	LUT3 #(
		.INIT('h70)
	) name10681 (
		_w6324_,
		_w7026_,
		_w10714_,
		_w10715_
	);
	LUT4 #(
		.INIT('h95aa)
	) name10682 (
		\a[5] ,
		_w35_,
		_w7562_,
		_w10715_,
		_w10716_
	);
	LUT2 #(
		.INIT('h2)
	) name10683 (
		_w10712_,
		_w10716_,
		_w10717_
	);
	LUT3 #(
		.INIT('h82)
	) name10684 (
		_w35_,
		_w7099_,
		_w7101_,
		_w10718_
	);
	LUT3 #(
		.INIT('h82)
	) name10685 (
		_w6324_,
		_w4030_,
		_w6952_,
		_w10719_
	);
	LUT2 #(
		.INIT('h8)
	) name10686 (
		_w5524_,
		_w7032_,
		_w10720_
	);
	LUT4 #(
		.INIT('h5060)
	) name10687 (
		_w4099_,
		_w4378_,
		_w6031_,
		_w6951_,
		_w10721_
	);
	LUT2 #(
		.INIT('h1)
	) name10688 (
		_w10720_,
		_w10721_,
		_w10722_
	);
	LUT2 #(
		.INIT('h4)
	) name10689 (
		_w10719_,
		_w10722_,
		_w10723_
	);
	LUT3 #(
		.INIT('h1e)
	) name10690 (
		_w10409_,
		_w10532_,
		_w10533_,
		_w10724_
	);
	LUT4 #(
		.INIT('h6500)
	) name10691 (
		\a[5] ,
		_w10718_,
		_w10723_,
		_w10724_,
		_w10725_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10692 (
		_w35_,
		_w7034_,
		_w7097_,
		_w7098_,
		_w10726_
	);
	LUT4 #(
		.INIT('h2228)
	) name10693 (
		_w6324_,
		_w4099_,
		_w4378_,
		_w6951_,
		_w10727_
	);
	LUT3 #(
		.INIT('h82)
	) name10694 (
		_w5524_,
		_w6947_,
		_w6949_,
		_w10728_
	);
	LUT3 #(
		.INIT('h07)
	) name10695 (
		_w6031_,
		_w7032_,
		_w10728_,
		_w10729_
	);
	LUT2 #(
		.INIT('h4)
	) name10696 (
		_w10727_,
		_w10729_,
		_w10730_
	);
	LUT4 #(
		.INIT('h54ab)
	) name10697 (
		_w10415_,
		_w10528_,
		_w10529_,
		_w10531_,
		_w10731_
	);
	LUT4 #(
		.INIT('h6500)
	) name10698 (
		\a[5] ,
		_w10726_,
		_w10730_,
		_w10731_,
		_w10732_
	);
	LUT4 #(
		.INIT('h04c8)
	) name10699 (
		_w4695_,
		_w5524_,
		_w6944_,
		_w6946_,
		_w10733_
	);
	LUT4 #(
		.INIT('h007d)
	) name10700 (
		_w6031_,
		_w6947_,
		_w6949_,
		_w10733_,
		_w10734_
	);
	LUT3 #(
		.INIT('h70)
	) name10701 (
		_w6324_,
		_w7032_,
		_w10734_,
		_w10735_
	);
	LUT4 #(
		.INIT('h95aa)
	) name10702 (
		\a[5] ,
		_w35_,
		_w7882_,
		_w10735_,
		_w10736_
	);
	LUT2 #(
		.INIT('h9)
	) name10703 (
		_w10528_,
		_w10530_,
		_w10737_
	);
	LUT2 #(
		.INIT('h4)
	) name10704 (
		_w10736_,
		_w10737_,
		_w10738_
	);
	LUT3 #(
		.INIT('h1e)
	) name10705 (
		_w10430_,
		_w10526_,
		_w10527_,
		_w10739_
	);
	LUT3 #(
		.INIT('h82)
	) name10706 (
		_w35_,
		_w7093_,
		_w7095_,
		_w10740_
	);
	LUT3 #(
		.INIT('h82)
	) name10707 (
		_w6324_,
		_w6947_,
		_w6949_,
		_w10741_
	);
	LUT2 #(
		.INIT('h8)
	) name10708 (
		_w5524_,
		_w7038_,
		_w10742_
	);
	LUT4 #(
		.INIT('h04c8)
	) name10709 (
		_w4695_,
		_w6031_,
		_w6944_,
		_w6946_,
		_w10743_
	);
	LUT2 #(
		.INIT('h1)
	) name10710 (
		_w10742_,
		_w10743_,
		_w10744_
	);
	LUT2 #(
		.INIT('h4)
	) name10711 (
		_w10741_,
		_w10744_,
		_w10745_
	);
	LUT4 #(
		.INIT('h4844)
	) name10712 (
		\a[5] ,
		_w10739_,
		_w10740_,
		_w10745_,
		_w10746_
	);
	LUT4 #(
		.INIT('h54ab)
	) name10713 (
		_w10436_,
		_w10522_,
		_w10523_,
		_w10525_,
		_w10747_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10714 (
		_w35_,
		_w7040_,
		_w7091_,
		_w7092_,
		_w10748_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10715 (
		_w6324_,
		_w4695_,
		_w6944_,
		_w6946_,
		_w10749_
	);
	LUT3 #(
		.INIT('h82)
	) name10716 (
		_w5524_,
		_w6940_,
		_w6942_,
		_w10750_
	);
	LUT3 #(
		.INIT('h07)
	) name10717 (
		_w6031_,
		_w7038_,
		_w10750_,
		_w10751_
	);
	LUT2 #(
		.INIT('h4)
	) name10718 (
		_w10749_,
		_w10751_,
		_w10752_
	);
	LUT4 #(
		.INIT('h4844)
	) name10719 (
		\a[5] ,
		_w10747_,
		_w10748_,
		_w10752_,
		_w10753_
	);
	LUT2 #(
		.INIT('h9)
	) name10720 (
		_w10522_,
		_w10524_,
		_w10754_
	);
	LUT4 #(
		.INIT('h5060)
	) name10721 (
		_w5067_,
		_w5282_,
		_w5524_,
		_w6939_,
		_w10755_
	);
	LUT4 #(
		.INIT('h007d)
	) name10722 (
		_w6031_,
		_w6940_,
		_w6942_,
		_w10755_,
		_w10756_
	);
	LUT3 #(
		.INIT('h70)
	) name10723 (
		_w6324_,
		_w7038_,
		_w10756_,
		_w10757_
	);
	LUT4 #(
		.INIT('h95aa)
	) name10724 (
		\a[5] ,
		_w35_,
		_w8018_,
		_w10757_,
		_w10758_
	);
	LUT2 #(
		.INIT('h2)
	) name10725 (
		_w10754_,
		_w10758_,
		_w10759_
	);
	LUT3 #(
		.INIT('h82)
	) name10726 (
		_w35_,
		_w7087_,
		_w7089_,
		_w10760_
	);
	LUT3 #(
		.INIT('h82)
	) name10727 (
		_w6324_,
		_w6940_,
		_w6942_,
		_w10761_
	);
	LUT2 #(
		.INIT('h8)
	) name10728 (
		_w5524_,
		_w7044_,
		_w10762_
	);
	LUT4 #(
		.INIT('h5060)
	) name10729 (
		_w5067_,
		_w5282_,
		_w6031_,
		_w6939_,
		_w10763_
	);
	LUT2 #(
		.INIT('h1)
	) name10730 (
		_w10762_,
		_w10763_,
		_w10764_
	);
	LUT2 #(
		.INIT('h4)
	) name10731 (
		_w10761_,
		_w10764_,
		_w10765_
	);
	LUT3 #(
		.INIT('h1e)
	) name10732 (
		_w10451_,
		_w10520_,
		_w10521_,
		_w10766_
	);
	LUT4 #(
		.INIT('h6500)
	) name10733 (
		\a[5] ,
		_w10760_,
		_w10765_,
		_w10766_,
		_w10767_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10734 (
		_w35_,
		_w7046_,
		_w7085_,
		_w7086_,
		_w10768_
	);
	LUT4 #(
		.INIT('h2228)
	) name10735 (
		_w6324_,
		_w5067_,
		_w5282_,
		_w6939_,
		_w10769_
	);
	LUT3 #(
		.INIT('h82)
	) name10736 (
		_w5524_,
		_w6935_,
		_w6937_,
		_w10770_
	);
	LUT3 #(
		.INIT('h07)
	) name10737 (
		_w6031_,
		_w7044_,
		_w10770_,
		_w10771_
	);
	LUT2 #(
		.INIT('h4)
	) name10738 (
		_w10769_,
		_w10771_,
		_w10772_
	);
	LUT4 #(
		.INIT('h54ab)
	) name10739 (
		_w10457_,
		_w10516_,
		_w10517_,
		_w10519_,
		_w10773_
	);
	LUT4 #(
		.INIT('h6500)
	) name10740 (
		\a[5] ,
		_w10768_,
		_w10772_,
		_w10773_,
		_w10774_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10741 (
		_w5524_,
		_w6043_,
		_w6933_,
		_w6934_,
		_w10775_
	);
	LUT4 #(
		.INIT('h007d)
	) name10742 (
		_w6031_,
		_w6935_,
		_w6937_,
		_w10775_,
		_w10776_
	);
	LUT3 #(
		.INIT('h70)
	) name10743 (
		_w6324_,
		_w7044_,
		_w10776_,
		_w10777_
	);
	LUT4 #(
		.INIT('h95aa)
	) name10744 (
		\a[5] ,
		_w35_,
		_w8005_,
		_w10777_,
		_w10778_
	);
	LUT2 #(
		.INIT('h9)
	) name10745 (
		_w10516_,
		_w10518_,
		_w10779_
	);
	LUT2 #(
		.INIT('h4)
	) name10746 (
		_w10778_,
		_w10779_,
		_w10780_
	);
	LUT3 #(
		.INIT('h1e)
	) name10747 (
		_w10472_,
		_w10514_,
		_w10515_,
		_w10781_
	);
	LUT3 #(
		.INIT('h82)
	) name10748 (
		_w35_,
		_w7081_,
		_w7083_,
		_w10782_
	);
	LUT3 #(
		.INIT('h82)
	) name10749 (
		_w6324_,
		_w6935_,
		_w6937_,
		_w10783_
	);
	LUT2 #(
		.INIT('h8)
	) name10750 (
		_w5524_,
		_w7050_,
		_w10784_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10751 (
		_w6031_,
		_w6043_,
		_w6933_,
		_w6934_,
		_w10785_
	);
	LUT2 #(
		.INIT('h1)
	) name10752 (
		_w10784_,
		_w10785_,
		_w10786_
	);
	LUT2 #(
		.INIT('h4)
	) name10753 (
		_w10783_,
		_w10786_,
		_w10787_
	);
	LUT4 #(
		.INIT('h4844)
	) name10754 (
		\a[5] ,
		_w10781_,
		_w10782_,
		_w10787_,
		_w10788_
	);
	LUT4 #(
		.INIT('h54ab)
	) name10755 (
		_w10479_,
		_w10510_,
		_w10511_,
		_w10513_,
		_w10789_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10756 (
		_w35_,
		_w7052_,
		_w7079_,
		_w7080_,
		_w10790_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10757 (
		_w6324_,
		_w6043_,
		_w6933_,
		_w6934_,
		_w10791_
	);
	LUT3 #(
		.INIT('h82)
	) name10758 (
		_w5524_,
		_w6929_,
		_w6931_,
		_w10792_
	);
	LUT3 #(
		.INIT('h07)
	) name10759 (
		_w6031_,
		_w7050_,
		_w10792_,
		_w10793_
	);
	LUT2 #(
		.INIT('h4)
	) name10760 (
		_w10791_,
		_w10793_,
		_w10794_
	);
	LUT4 #(
		.INIT('h4844)
	) name10761 (
		\a[5] ,
		_w10789_,
		_w10790_,
		_w10794_,
		_w10795_
	);
	LUT2 #(
		.INIT('h9)
	) name10762 (
		_w10510_,
		_w10512_,
		_w10796_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10763 (
		_w5524_,
		_w6645_,
		_w6926_,
		_w6928_,
		_w10797_
	);
	LUT4 #(
		.INIT('h007d)
	) name10764 (
		_w6031_,
		_w6929_,
		_w6931_,
		_w10797_,
		_w10798_
	);
	LUT3 #(
		.INIT('h70)
	) name10765 (
		_w6324_,
		_w7050_,
		_w10798_,
		_w10799_
	);
	LUT4 #(
		.INIT('h95aa)
	) name10766 (
		\a[5] ,
		_w35_,
		_w8227_,
		_w10799_,
		_w10800_
	);
	LUT2 #(
		.INIT('h2)
	) name10767 (
		_w10796_,
		_w10800_,
		_w10801_
	);
	LUT3 #(
		.INIT('h82)
	) name10768 (
		_w35_,
		_w7075_,
		_w7077_,
		_w10802_
	);
	LUT3 #(
		.INIT('h82)
	) name10769 (
		_w6324_,
		_w6929_,
		_w6931_,
		_w10803_
	);
	LUT2 #(
		.INIT('h8)
	) name10770 (
		_w5524_,
		_w7056_,
		_w10804_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10771 (
		_w6031_,
		_w6645_,
		_w6926_,
		_w6928_,
		_w10805_
	);
	LUT2 #(
		.INIT('h1)
	) name10772 (
		_w10804_,
		_w10805_,
		_w10806_
	);
	LUT2 #(
		.INIT('h4)
	) name10773 (
		_w10803_,
		_w10806_,
		_w10807_
	);
	LUT2 #(
		.INIT('h9)
	) name10774 (
		_w10507_,
		_w10509_,
		_w10808_
	);
	LUT4 #(
		.INIT('h6500)
	) name10775 (
		\a[5] ,
		_w10802_,
		_w10807_,
		_w10808_,
		_w10809_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10776 (
		_w35_,
		_w7058_,
		_w7073_,
		_w7074_,
		_w10810_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10777 (
		_w6324_,
		_w6645_,
		_w6926_,
		_w6928_,
		_w10811_
	);
	LUT3 #(
		.INIT('h82)
	) name10778 (
		_w5524_,
		_w6922_,
		_w6924_,
		_w10812_
	);
	LUT3 #(
		.INIT('h07)
	) name10779 (
		_w6031_,
		_w7056_,
		_w10812_,
		_w10813_
	);
	LUT2 #(
		.INIT('h4)
	) name10780 (
		_w10811_,
		_w10813_,
		_w10814_
	);
	LUT4 #(
		.INIT('h9a65)
	) name10781 (
		\a[8] ,
		_w10500_,
		_w10504_,
		_w10505_,
		_w10815_
	);
	LUT4 #(
		.INIT('h6500)
	) name10782 (
		\a[5] ,
		_w10810_,
		_w10814_,
		_w10815_,
		_w10816_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10783 (
		_w5524_,
		_w6669_,
		_w6919_,
		_w6921_,
		_w10817_
	);
	LUT4 #(
		.INIT('h007d)
	) name10784 (
		_w6031_,
		_w6922_,
		_w6924_,
		_w10817_,
		_w10818_
	);
	LUT3 #(
		.INIT('h70)
	) name10785 (
		_w6324_,
		_w7056_,
		_w10818_,
		_w10819_
	);
	LUT4 #(
		.INIT('h95aa)
	) name10786 (
		\a[5] ,
		_w35_,
		_w8298_,
		_w10819_,
		_w10820_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name10787 (
		\a[8] ,
		_w10492_,
		_w10489_,
		_w10491_,
		_w10821_
	);
	LUT3 #(
		.INIT('h4b)
	) name10788 (
		_w10495_,
		_w10498_,
		_w10821_,
		_w10822_
	);
	LUT2 #(
		.INIT('h4)
	) name10789 (
		_w10820_,
		_w10822_,
		_w10823_
	);
	LUT3 #(
		.INIT('h82)
	) name10790 (
		_w35_,
		_w7069_,
		_w7071_,
		_w10824_
	);
	LUT3 #(
		.INIT('h82)
	) name10791 (
		_w6324_,
		_w6922_,
		_w6924_,
		_w10825_
	);
	LUT2 #(
		.INIT('h8)
	) name10792 (
		_w5524_,
		_w7062_,
		_w10826_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10793 (
		_w6031_,
		_w6669_,
		_w6919_,
		_w6921_,
		_w10827_
	);
	LUT2 #(
		.INIT('h1)
	) name10794 (
		_w10826_,
		_w10827_,
		_w10828_
	);
	LUT2 #(
		.INIT('h4)
	) name10795 (
		_w10825_,
		_w10828_,
		_w10829_
	);
	LUT2 #(
		.INIT('h8)
	) name10796 (
		\a[8] ,
		_w10492_,
		_w10830_
	);
	LUT3 #(
		.INIT('h4b)
	) name10797 (
		_w10489_,
		_w10491_,
		_w10830_,
		_w10831_
	);
	LUT4 #(
		.INIT('h6500)
	) name10798 (
		\a[5] ,
		_w10824_,
		_w10829_,
		_w10831_,
		_w10832_
	);
	LUT4 #(
		.INIT('h2882)
	) name10799 (
		_w35_,
		_w6914_,
		_w6916_,
		_w7067_,
		_w10833_
	);
	LUT4 #(
		.INIT('ha802)
	) name10800 (
		_w6031_,
		_w6689_,
		_w6911_,
		_w6913_,
		_w10834_
	);
	LUT4 #(
		.INIT('h007d)
	) name10801 (
		_w6324_,
		_w6914_,
		_w6916_,
		_w10834_,
		_w10835_
	);
	LUT4 #(
		.INIT('h5401)
	) name10802 (
		_w34_,
		_w6689_,
		_w6911_,
		_w6913_,
		_w10836_
	);
	LUT2 #(
		.INIT('h2)
	) name10803 (
		\a[5] ,
		_w10836_,
		_w10837_
	);
	LUT3 #(
		.INIT('h40)
	) name10804 (
		_w10833_,
		_w10835_,
		_w10837_,
		_w10838_
	);
	LUT3 #(
		.INIT('h28)
	) name10805 (
		_w35_,
		_w7062_,
		_w8358_,
		_w10839_
	);
	LUT4 #(
		.INIT('ha802)
	) name10806 (
		_w5524_,
		_w6689_,
		_w6911_,
		_w6913_,
		_w10840_
	);
	LUT4 #(
		.INIT('h007d)
	) name10807 (
		_w6031_,
		_w6914_,
		_w6916_,
		_w10840_,
		_w10841_
	);
	LUT3 #(
		.INIT('h70)
	) name10808 (
		_w6324_,
		_w7062_,
		_w10841_,
		_w10842_
	);
	LUT4 #(
		.INIT('h0800)
	) name10809 (
		_w10492_,
		_w10838_,
		_w10839_,
		_w10842_,
		_w10843_
	);
	LUT3 #(
		.INIT('h28)
	) name10810 (
		_w35_,
		_w7065_,
		_w7068_,
		_w10844_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10811 (
		_w6324_,
		_w6669_,
		_w6919_,
		_w6921_,
		_w10845_
	);
	LUT3 #(
		.INIT('h82)
	) name10812 (
		_w5524_,
		_w6914_,
		_w6916_,
		_w10846_
	);
	LUT3 #(
		.INIT('h07)
	) name10813 (
		_w6031_,
		_w7062_,
		_w10846_,
		_w10847_
	);
	LUT2 #(
		.INIT('h4)
	) name10814 (
		_w10845_,
		_w10847_,
		_w10848_
	);
	LUT4 #(
		.INIT('ha6aa)
	) name10815 (
		_w10492_,
		_w10838_,
		_w10839_,
		_w10842_,
		_w10849_
	);
	LUT4 #(
		.INIT('h6500)
	) name10816 (
		\a[5] ,
		_w10844_,
		_w10848_,
		_w10849_,
		_w10850_
	);
	LUT2 #(
		.INIT('h1)
	) name10817 (
		_w10843_,
		_w10850_,
		_w10851_
	);
	LUT4 #(
		.INIT('h009a)
	) name10818 (
		\a[5] ,
		_w10824_,
		_w10829_,
		_w10831_,
		_w10852_
	);
	LUT4 #(
		.INIT('h9a65)
	) name10819 (
		\a[5] ,
		_w10824_,
		_w10829_,
		_w10831_,
		_w10853_
	);
	LUT3 #(
		.INIT('h54)
	) name10820 (
		_w10832_,
		_w10851_,
		_w10852_,
		_w10854_
	);
	LUT2 #(
		.INIT('h2)
	) name10821 (
		_w10820_,
		_w10822_,
		_w10855_
	);
	LUT2 #(
		.INIT('h9)
	) name10822 (
		_w10820_,
		_w10822_,
		_w10856_
	);
	LUT4 #(
		.INIT('h9a65)
	) name10823 (
		\a[5] ,
		_w10810_,
		_w10814_,
		_w10815_,
		_w10857_
	);
	LUT4 #(
		.INIT('h4d00)
	) name10824 (
		_w10820_,
		_w10822_,
		_w10854_,
		_w10857_,
		_w10858_
	);
	LUT4 #(
		.INIT('h9a65)
	) name10825 (
		\a[5] ,
		_w10802_,
		_w10807_,
		_w10808_,
		_w10859_
	);
	LUT4 #(
		.INIT('h0155)
	) name10826 (
		_w10809_,
		_w10816_,
		_w10858_,
		_w10859_,
		_w10860_
	);
	LUT2 #(
		.INIT('h4)
	) name10827 (
		_w10796_,
		_w10800_,
		_w10861_
	);
	LUT2 #(
		.INIT('h9)
	) name10828 (
		_w10796_,
		_w10800_,
		_w10862_
	);
	LUT4 #(
		.INIT('h9699)
	) name10829 (
		\a[5] ,
		_w10789_,
		_w10790_,
		_w10794_,
		_w10863_
	);
	LUT4 #(
		.INIT('h2b00)
	) name10830 (
		_w10796_,
		_w10800_,
		_w10860_,
		_w10863_,
		_w10864_
	);
	LUT4 #(
		.INIT('h9699)
	) name10831 (
		\a[5] ,
		_w10781_,
		_w10782_,
		_w10787_,
		_w10865_
	);
	LUT4 #(
		.INIT('h0155)
	) name10832 (
		_w10788_,
		_w10795_,
		_w10864_,
		_w10865_,
		_w10866_
	);
	LUT2 #(
		.INIT('h2)
	) name10833 (
		_w10778_,
		_w10779_,
		_w10867_
	);
	LUT2 #(
		.INIT('h9)
	) name10834 (
		_w10778_,
		_w10779_,
		_w10868_
	);
	LUT4 #(
		.INIT('h9a65)
	) name10835 (
		\a[5] ,
		_w10768_,
		_w10772_,
		_w10773_,
		_w10869_
	);
	LUT4 #(
		.INIT('h4d00)
	) name10836 (
		_w10778_,
		_w10779_,
		_w10866_,
		_w10869_,
		_w10870_
	);
	LUT4 #(
		.INIT('h9a65)
	) name10837 (
		\a[5] ,
		_w10760_,
		_w10765_,
		_w10766_,
		_w10871_
	);
	LUT4 #(
		.INIT('h0155)
	) name10838 (
		_w10767_,
		_w10774_,
		_w10870_,
		_w10871_,
		_w10872_
	);
	LUT2 #(
		.INIT('h4)
	) name10839 (
		_w10754_,
		_w10758_,
		_w10873_
	);
	LUT2 #(
		.INIT('h9)
	) name10840 (
		_w10754_,
		_w10758_,
		_w10874_
	);
	LUT4 #(
		.INIT('h9699)
	) name10841 (
		\a[5] ,
		_w10747_,
		_w10748_,
		_w10752_,
		_w10875_
	);
	LUT4 #(
		.INIT('h2b00)
	) name10842 (
		_w10754_,
		_w10758_,
		_w10872_,
		_w10875_,
		_w10876_
	);
	LUT4 #(
		.INIT('h9699)
	) name10843 (
		\a[5] ,
		_w10739_,
		_w10740_,
		_w10745_,
		_w10877_
	);
	LUT4 #(
		.INIT('h0155)
	) name10844 (
		_w10746_,
		_w10753_,
		_w10876_,
		_w10877_,
		_w10878_
	);
	LUT2 #(
		.INIT('h2)
	) name10845 (
		_w10736_,
		_w10737_,
		_w10879_
	);
	LUT2 #(
		.INIT('h9)
	) name10846 (
		_w10736_,
		_w10737_,
		_w10880_
	);
	LUT4 #(
		.INIT('h9a65)
	) name10847 (
		\a[5] ,
		_w10726_,
		_w10730_,
		_w10731_,
		_w10881_
	);
	LUT4 #(
		.INIT('h4d00)
	) name10848 (
		_w10736_,
		_w10737_,
		_w10878_,
		_w10881_,
		_w10882_
	);
	LUT4 #(
		.INIT('h9a65)
	) name10849 (
		\a[5] ,
		_w10718_,
		_w10723_,
		_w10724_,
		_w10883_
	);
	LUT4 #(
		.INIT('h0155)
	) name10850 (
		_w10725_,
		_w10732_,
		_w10882_,
		_w10883_,
		_w10884_
	);
	LUT2 #(
		.INIT('h4)
	) name10851 (
		_w10712_,
		_w10716_,
		_w10885_
	);
	LUT2 #(
		.INIT('h9)
	) name10852 (
		_w10712_,
		_w10716_,
		_w10886_
	);
	LUT4 #(
		.INIT('h9699)
	) name10853 (
		\a[5] ,
		_w10705_,
		_w10706_,
		_w10710_,
		_w10887_
	);
	LUT4 #(
		.INIT('h2b00)
	) name10854 (
		_w10712_,
		_w10716_,
		_w10884_,
		_w10887_,
		_w10888_
	);
	LUT4 #(
		.INIT('h9699)
	) name10855 (
		\a[5] ,
		_w10697_,
		_w10698_,
		_w10703_,
		_w10889_
	);
	LUT4 #(
		.INIT('h0155)
	) name10856 (
		_w10704_,
		_w10711_,
		_w10888_,
		_w10889_,
		_w10890_
	);
	LUT2 #(
		.INIT('h2)
	) name10857 (
		_w10694_,
		_w10695_,
		_w10891_
	);
	LUT2 #(
		.INIT('h9)
	) name10858 (
		_w10694_,
		_w10695_,
		_w10892_
	);
	LUT4 #(
		.INIT('h9a65)
	) name10859 (
		\a[5] ,
		_w10684_,
		_w10688_,
		_w10689_,
		_w10893_
	);
	LUT4 #(
		.INIT('h4d00)
	) name10860 (
		_w10694_,
		_w10695_,
		_w10890_,
		_w10893_,
		_w10894_
	);
	LUT4 #(
		.INIT('h9a65)
	) name10861 (
		\a[5] ,
		_w10676_,
		_w10681_,
		_w10682_,
		_w10895_
	);
	LUT4 #(
		.INIT('h0155)
	) name10862 (
		_w10683_,
		_w10690_,
		_w10894_,
		_w10895_,
		_w10896_
	);
	LUT2 #(
		.INIT('h4)
	) name10863 (
		_w10670_,
		_w10674_,
		_w10897_
	);
	LUT2 #(
		.INIT('h9)
	) name10864 (
		_w10670_,
		_w10674_,
		_w10898_
	);
	LUT4 #(
		.INIT('h9699)
	) name10865 (
		\a[5] ,
		_w10663_,
		_w10664_,
		_w10668_,
		_w10899_
	);
	LUT4 #(
		.INIT('h2b00)
	) name10866 (
		_w10670_,
		_w10674_,
		_w10896_,
		_w10899_,
		_w10900_
	);
	LUT4 #(
		.INIT('h9a65)
	) name10867 (
		\a[5] ,
		_w10655_,
		_w10660_,
		_w10661_,
		_w10901_
	);
	LUT4 #(
		.INIT('h0155)
	) name10868 (
		_w10662_,
		_w10669_,
		_w10900_,
		_w10901_,
		_w10902_
	);
	LUT2 #(
		.INIT('h2)
	) name10869 (
		_w10652_,
		_w10653_,
		_w10903_
	);
	LUT2 #(
		.INIT('h9)
	) name10870 (
		_w10652_,
		_w10653_,
		_w10904_
	);
	LUT4 #(
		.INIT('h9a65)
	) name10871 (
		\a[5] ,
		_w10642_,
		_w10646_,
		_w10647_,
		_w10905_
	);
	LUT4 #(
		.INIT('h4d00)
	) name10872 (
		_w10652_,
		_w10653_,
		_w10902_,
		_w10905_,
		_w10906_
	);
	LUT4 #(
		.INIT('h9a65)
	) name10873 (
		\a[5] ,
		_w10634_,
		_w10639_,
		_w10640_,
		_w10907_
	);
	LUT4 #(
		.INIT('h0155)
	) name10874 (
		_w10641_,
		_w10648_,
		_w10906_,
		_w10907_,
		_w10908_
	);
	LUT2 #(
		.INIT('h2)
	) name10875 (
		_w10631_,
		_w10632_,
		_w10909_
	);
	LUT2 #(
		.INIT('h9)
	) name10876 (
		_w10631_,
		_w10632_,
		_w10910_
	);
	LUT4 #(
		.INIT('h9a65)
	) name10877 (
		\a[5] ,
		_w10621_,
		_w10625_,
		_w10626_,
		_w10911_
	);
	LUT4 #(
		.INIT('h4d00)
	) name10878 (
		_w10631_,
		_w10632_,
		_w10908_,
		_w10911_,
		_w10912_
	);
	LUT4 #(
		.INIT('h9a65)
	) name10879 (
		\a[5] ,
		_w10613_,
		_w10618_,
		_w10619_,
		_w10913_
	);
	LUT4 #(
		.INIT('h0155)
	) name10880 (
		_w10620_,
		_w10627_,
		_w10912_,
		_w10913_,
		_w10914_
	);
	LUT2 #(
		.INIT('h2)
	) name10881 (
		_w10610_,
		_w10611_,
		_w10915_
	);
	LUT2 #(
		.INIT('h9)
	) name10882 (
		_w10610_,
		_w10611_,
		_w10916_
	);
	LUT4 #(
		.INIT('h9a65)
	) name10883 (
		\a[5] ,
		_w10600_,
		_w10604_,
		_w10605_,
		_w10917_
	);
	LUT4 #(
		.INIT('h4d00)
	) name10884 (
		_w10610_,
		_w10611_,
		_w10914_,
		_w10917_,
		_w10918_
	);
	LUT2 #(
		.INIT('h1)
	) name10885 (
		_w10606_,
		_w10918_,
		_w10919_
	);
	LUT3 #(
		.INIT('h69)
	) name10886 (
		\a[2] ,
		_w10593_,
		_w10595_,
		_w10920_
	);
	LUT2 #(
		.INIT('h4)
	) name10887 (
		_w10919_,
		_w10920_,
		_w10921_
	);
	LUT2 #(
		.INIT('h9)
	) name10888 (
		_w10919_,
		_w10920_,
		_w10922_
	);
	LUT4 #(
		.INIT('h54ab)
	) name10889 (
		_w10612_,
		_w10914_,
		_w10915_,
		_w10917_,
		_w10923_
	);
	LUT4 #(
		.INIT('h0a02)
	) name10890 (
		_w6335_,
		_w7169_,
		_w7419_,
		_w7686_,
		_w10924_
	);
	LUT3 #(
		.INIT('h28)
	) name10891 (
		_w6334_,
		_w7136_,
		_w7168_,
		_w10925_
	);
	LUT3 #(
		.INIT('h40)
	) name10892 (
		_w6657_,
		_w7136_,
		_w7167_,
		_w10926_
	);
	LUT3 #(
		.INIT('h31)
	) name10893 (
		_w10591_,
		_w10925_,
		_w10926_,
		_w10927_
	);
	LUT3 #(
		.INIT('h9a)
	) name10894 (
		\a[2] ,
		_w10924_,
		_w10927_,
		_w10928_
	);
	LUT4 #(
		.INIT('h4844)
	) name10895 (
		\a[2] ,
		_w10923_,
		_w10924_,
		_w10927_,
		_w10929_
	);
	LUT2 #(
		.INIT('h9)
	) name10896 (
		_w10914_,
		_w10916_,
		_w10930_
	);
	LUT3 #(
		.INIT('h28)
	) name10897 (
		_w6650_,
		_w7136_,
		_w7168_,
		_w10931_
	);
	LUT4 #(
		.INIT('h028a)
	) name10898 (
		_w6657_,
		_w7136_,
		_w7166_,
		_w7167_,
		_w10932_
	);
	LUT4 #(
		.INIT('h04c8)
	) name10899 (
		_w2411_,
		_w6334_,
		_w6983_,
		_w6993_,
		_w10933_
	);
	LUT3 #(
		.INIT('h01)
	) name10900 (
		_w10932_,
		_w10933_,
		_w10931_,
		_w10934_
	);
	LUT4 #(
		.INIT('h95aa)
	) name10901 (
		\a[2] ,
		_w6335_,
		_w7696_,
		_w10934_,
		_w10935_
	);
	LUT2 #(
		.INIT('h2)
	) name10902 (
		_w10930_,
		_w10935_,
		_w10936_
	);
	LUT3 #(
		.INIT('h1e)
	) name10903 (
		_w10627_,
		_w10912_,
		_w10913_,
		_w10937_
	);
	LUT3 #(
		.INIT('h82)
	) name10904 (
		_w6335_,
		_w7135_,
		_w7172_,
		_w10938_
	);
	LUT3 #(
		.INIT('h28)
	) name10905 (
		_w6657_,
		_w7136_,
		_w7168_,
		_w10939_
	);
	LUT2 #(
		.INIT('h8)
	) name10906 (
		_w6334_,
		_w6996_,
		_w10940_
	);
	LUT4 #(
		.INIT('h04c8)
	) name10907 (
		_w2411_,
		_w6650_,
		_w6983_,
		_w6993_,
		_w10941_
	);
	LUT2 #(
		.INIT('h1)
	) name10908 (
		_w10940_,
		_w10941_,
		_w10942_
	);
	LUT2 #(
		.INIT('h4)
	) name10909 (
		_w10939_,
		_w10942_,
		_w10943_
	);
	LUT3 #(
		.INIT('h9a)
	) name10910 (
		\a[2] ,
		_w10938_,
		_w10943_,
		_w10944_
	);
	LUT4 #(
		.INIT('h4844)
	) name10911 (
		\a[2] ,
		_w10937_,
		_w10938_,
		_w10943_,
		_w10945_
	);
	LUT4 #(
		.INIT('h54ab)
	) name10912 (
		_w10633_,
		_w10908_,
		_w10909_,
		_w10911_,
		_w10946_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10913 (
		_w6335_,
		_w6998_,
		_w7133_,
		_w7134_,
		_w10947_
	);
	LUT4 #(
		.INIT('h04c8)
	) name10914 (
		_w2411_,
		_w6657_,
		_w6983_,
		_w6993_,
		_w10948_
	);
	LUT3 #(
		.INIT('h84)
	) name10915 (
		_w2546_,
		_w6334_,
		_w6981_,
		_w10949_
	);
	LUT3 #(
		.INIT('h07)
	) name10916 (
		_w6650_,
		_w6996_,
		_w10949_,
		_w10950_
	);
	LUT2 #(
		.INIT('h4)
	) name10917 (
		_w10948_,
		_w10950_,
		_w10951_
	);
	LUT3 #(
		.INIT('h9a)
	) name10918 (
		\a[2] ,
		_w10947_,
		_w10951_,
		_w10952_
	);
	LUT4 #(
		.INIT('h4844)
	) name10919 (
		\a[2] ,
		_w10946_,
		_w10947_,
		_w10951_,
		_w10953_
	);
	LUT2 #(
		.INIT('h9)
	) name10920 (
		_w10908_,
		_w10910_,
		_w10954_
	);
	LUT4 #(
		.INIT('h04c8)
	) name10921 (
		_w2622_,
		_w6334_,
		_w6978_,
		_w6980_,
		_w10955_
	);
	LUT4 #(
		.INIT('h007b)
	) name10922 (
		_w2546_,
		_w6650_,
		_w6981_,
		_w10955_,
		_w10956_
	);
	LUT3 #(
		.INIT('h70)
	) name10923 (
		_w6657_,
		_w6996_,
		_w10956_,
		_w10957_
	);
	LUT4 #(
		.INIT('h95aa)
	) name10924 (
		\a[2] ,
		_w6335_,
		_w7500_,
		_w10957_,
		_w10958_
	);
	LUT2 #(
		.INIT('h2)
	) name10925 (
		_w10954_,
		_w10958_,
		_w10959_
	);
	LUT3 #(
		.INIT('h1e)
	) name10926 (
		_w10648_,
		_w10906_,
		_w10907_,
		_w10960_
	);
	LUT3 #(
		.INIT('h82)
	) name10927 (
		_w6335_,
		_w7129_,
		_w7131_,
		_w10961_
	);
	LUT3 #(
		.INIT('h84)
	) name10928 (
		_w2546_,
		_w6657_,
		_w6981_,
		_w10962_
	);
	LUT2 #(
		.INIT('h8)
	) name10929 (
		_w6334_,
		_w7002_,
		_w10963_
	);
	LUT4 #(
		.INIT('h04c8)
	) name10930 (
		_w2622_,
		_w6650_,
		_w6978_,
		_w6980_,
		_w10964_
	);
	LUT2 #(
		.INIT('h1)
	) name10931 (
		_w10963_,
		_w10964_,
		_w10965_
	);
	LUT2 #(
		.INIT('h4)
	) name10932 (
		_w10962_,
		_w10965_,
		_w10966_
	);
	LUT3 #(
		.INIT('h9a)
	) name10933 (
		\a[2] ,
		_w10961_,
		_w10966_,
		_w10967_
	);
	LUT4 #(
		.INIT('h4844)
	) name10934 (
		\a[2] ,
		_w10960_,
		_w10961_,
		_w10966_,
		_w10968_
	);
	LUT4 #(
		.INIT('h54ab)
	) name10935 (
		_w10654_,
		_w10902_,
		_w10903_,
		_w10905_,
		_w10969_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10936 (
		_w6335_,
		_w7004_,
		_w7127_,
		_w7128_,
		_w10970_
	);
	LUT4 #(
		.INIT('h04c8)
	) name10937 (
		_w2622_,
		_w6657_,
		_w6978_,
		_w6980_,
		_w10971_
	);
	LUT3 #(
		.INIT('h84)
	) name10938 (
		_w2872_,
		_w6334_,
		_w6975_,
		_w10972_
	);
	LUT3 #(
		.INIT('h07)
	) name10939 (
		_w6650_,
		_w7002_,
		_w10972_,
		_w10973_
	);
	LUT2 #(
		.INIT('h4)
	) name10940 (
		_w10971_,
		_w10973_,
		_w10974_
	);
	LUT3 #(
		.INIT('h9a)
	) name10941 (
		\a[2] ,
		_w10970_,
		_w10974_,
		_w10975_
	);
	LUT4 #(
		.INIT('h4844)
	) name10942 (
		\a[2] ,
		_w10969_,
		_w10970_,
		_w10974_,
		_w10976_
	);
	LUT2 #(
		.INIT('h9)
	) name10943 (
		_w10902_,
		_w10904_,
		_w10977_
	);
	LUT4 #(
		.INIT('h04c8)
	) name10944 (
		_w2983_,
		_w6334_,
		_w6972_,
		_w6974_,
		_w10978_
	);
	LUT4 #(
		.INIT('h007b)
	) name10945 (
		_w2872_,
		_w6650_,
		_w6975_,
		_w10978_,
		_w10979_
	);
	LUT3 #(
		.INIT('h70)
	) name10946 (
		_w6657_,
		_w7002_,
		_w10979_,
		_w10980_
	);
	LUT4 #(
		.INIT('h95aa)
	) name10947 (
		\a[2] ,
		_w6335_,
		_w7426_,
		_w10980_,
		_w10981_
	);
	LUT2 #(
		.INIT('h2)
	) name10948 (
		_w10977_,
		_w10981_,
		_w10982_
	);
	LUT3 #(
		.INIT('h1e)
	) name10949 (
		_w10669_,
		_w10900_,
		_w10901_,
		_w10983_
	);
	LUT3 #(
		.INIT('h82)
	) name10950 (
		_w6335_,
		_w7123_,
		_w7125_,
		_w10984_
	);
	LUT3 #(
		.INIT('h84)
	) name10951 (
		_w2872_,
		_w6657_,
		_w6975_,
		_w10985_
	);
	LUT2 #(
		.INIT('h8)
	) name10952 (
		_w6334_,
		_w7008_,
		_w10986_
	);
	LUT4 #(
		.INIT('h04c8)
	) name10953 (
		_w2983_,
		_w6650_,
		_w6972_,
		_w6974_,
		_w10987_
	);
	LUT2 #(
		.INIT('h1)
	) name10954 (
		_w10986_,
		_w10987_,
		_w10988_
	);
	LUT2 #(
		.INIT('h4)
	) name10955 (
		_w10985_,
		_w10988_,
		_w10989_
	);
	LUT3 #(
		.INIT('h9a)
	) name10956 (
		\a[2] ,
		_w10984_,
		_w10989_,
		_w10990_
	);
	LUT4 #(
		.INIT('h4844)
	) name10957 (
		\a[2] ,
		_w10983_,
		_w10984_,
		_w10989_,
		_w10991_
	);
	LUT4 #(
		.INIT('h9699)
	) name10958 (
		\a[2] ,
		_w10983_,
		_w10984_,
		_w10989_,
		_w10992_
	);
	LUT4 #(
		.INIT('h54ab)
	) name10959 (
		_w10675_,
		_w10896_,
		_w10897_,
		_w10899_,
		_w10993_
	);
	LUT2 #(
		.INIT('h9)
	) name10960 (
		_w10896_,
		_w10898_,
		_w10994_
	);
	LUT3 #(
		.INIT('h1e)
	) name10961 (
		_w10690_,
		_w10894_,
		_w10895_,
		_w10995_
	);
	LUT4 #(
		.INIT('h54ab)
	) name10962 (
		_w10696_,
		_w10890_,
		_w10891_,
		_w10893_,
		_w10996_
	);
	LUT4 #(
		.INIT('h5060)
	) name10963 (
		_w3409_,
		_w3650_,
		_w6334_,
		_w6959_,
		_w10997_
	);
	LUT4 #(
		.INIT('h007d)
	) name10964 (
		_w6650_,
		_w6960_,
		_w6962_,
		_w10997_,
		_w10998_
	);
	LUT3 #(
		.INIT('h70)
	) name10965 (
		_w6657_,
		_w7014_,
		_w10998_,
		_w10999_
	);
	LUT4 #(
		.INIT('h95aa)
	) name10966 (
		\a[2] ,
		_w6335_,
		_w7291_,
		_w10999_,
		_w11000_
	);
	LUT2 #(
		.INIT('h9)
	) name10967 (
		_w10890_,
		_w10892_,
		_w11001_
	);
	LUT2 #(
		.INIT('h2)
	) name10968 (
		_w11000_,
		_w11001_,
		_w11002_
	);
	LUT2 #(
		.INIT('h4)
	) name10969 (
		_w11000_,
		_w11001_,
		_w11003_
	);
	LUT3 #(
		.INIT('h1e)
	) name10970 (
		_w10711_,
		_w10888_,
		_w10889_,
		_w11004_
	);
	LUT3 #(
		.INIT('h82)
	) name10971 (
		_w6335_,
		_w7111_,
		_w7113_,
		_w11005_
	);
	LUT3 #(
		.INIT('h82)
	) name10972 (
		_w6657_,
		_w6960_,
		_w6962_,
		_w11006_
	);
	LUT2 #(
		.INIT('h8)
	) name10973 (
		_w6334_,
		_w7020_,
		_w11007_
	);
	LUT4 #(
		.INIT('h5060)
	) name10974 (
		_w3409_,
		_w3650_,
		_w6650_,
		_w6959_,
		_w11008_
	);
	LUT2 #(
		.INIT('h1)
	) name10975 (
		_w11007_,
		_w11008_,
		_w11009_
	);
	LUT2 #(
		.INIT('h4)
	) name10976 (
		_w11006_,
		_w11009_,
		_w11010_
	);
	LUT4 #(
		.INIT('h2122)
	) name10977 (
		\a[2] ,
		_w11004_,
		_w11005_,
		_w11010_,
		_w11011_
	);
	LUT4 #(
		.INIT('h4844)
	) name10978 (
		\a[2] ,
		_w11004_,
		_w11005_,
		_w11010_,
		_w11012_
	);
	LUT4 #(
		.INIT('h54ab)
	) name10979 (
		_w10717_,
		_w10884_,
		_w10885_,
		_w10887_,
		_w11013_
	);
	LUT4 #(
		.INIT('h02a8)
	) name10980 (
		_w6335_,
		_w7022_,
		_w7109_,
		_w7110_,
		_w11014_
	);
	LUT4 #(
		.INIT('h5060)
	) name10981 (
		_w3409_,
		_w3650_,
		_w6657_,
		_w6959_,
		_w11015_
	);
	LUT3 #(
		.INIT('h84)
	) name10982 (
		_w3706_,
		_w6334_,
		_w6957_,
		_w11016_
	);
	LUT3 #(
		.INIT('h07)
	) name10983 (
		_w6650_,
		_w7020_,
		_w11016_,
		_w11017_
	);
	LUT2 #(
		.INIT('h4)
	) name10984 (
		_w11015_,
		_w11017_,
		_w11018_
	);
	LUT4 #(
		.INIT('h2122)
	) name10985 (
		\a[2] ,
		_w11013_,
		_w11014_,
		_w11018_,
		_w11019_
	);
	LUT4 #(
		.INIT('h4844)
	) name10986 (
		\a[2] ,
		_w11013_,
		_w11014_,
		_w11018_,
		_w11020_
	);
	LUT2 #(
		.INIT('h9)
	) name10987 (
		_w10884_,
		_w10886_,
		_w11021_
	);
	LUT4 #(
		.INIT('h04c8)
	) name10988 (
		_w3882_,
		_w6334_,
		_w6954_,
		_w6956_,
		_w11022_
	);
	LUT4 #(
		.INIT('h007b)
	) name10989 (
		_w3706_,
		_w6650_,
		_w6957_,
		_w11022_,
		_w11023_
	);
	LUT3 #(
		.INIT('h70)
	) name10990 (
		_w6657_,
		_w7020_,
		_w11023_,
		_w11024_
	);
	LUT4 #(
		.INIT('h6a55)
	) name10991 (
		\a[2] ,
		_w6335_,
		_w7465_,
		_w11024_,
		_w11025_
	);
	LUT3 #(
		.INIT('h82)
	) name10992 (
		_w6335_,
		_w7105_,
		_w7107_,
		_w11026_
	);
	LUT3 #(
		.INIT('h84)
	) name10993 (
		_w3706_,
		_w6657_,
		_w6957_,
		_w11027_
	);
	LUT2 #(
		.INIT('h8)
	) name10994 (
		_w6334_,
		_w7026_,
		_w11028_
	);
	LUT4 #(
		.INIT('h04c8)
	) name10995 (
		_w3882_,
		_w6650_,
		_w6954_,
		_w6956_,
		_w11029_
	);
	LUT2 #(
		.INIT('h1)
	) name10996 (
		_w11028_,
		_w11029_,
		_w11030_
	);
	LUT2 #(
		.INIT('h4)
	) name10997 (
		_w11027_,
		_w11030_,
		_w11031_
	);
	LUT3 #(
		.INIT('h9a)
	) name10998 (
		\a[2] ,
		_w11026_,
		_w11031_,
		_w11032_
	);
	LUT3 #(
		.INIT('h1e)
	) name10999 (
		_w10732_,
		_w10882_,
		_w10883_,
		_w11033_
	);
	LUT4 #(
		.INIT('h54ab)
	) name11000 (
		_w10738_,
		_w10878_,
		_w10879_,
		_w10881_,
		_w11034_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11001 (
		_w6335_,
		_w7028_,
		_w7103_,
		_w7104_,
		_w11035_
	);
	LUT4 #(
		.INIT('h04c8)
	) name11002 (
		_w3882_,
		_w6657_,
		_w6954_,
		_w6956_,
		_w11036_
	);
	LUT3 #(
		.INIT('h84)
	) name11003 (
		_w4030_,
		_w6334_,
		_w6952_,
		_w11037_
	);
	LUT3 #(
		.INIT('h07)
	) name11004 (
		_w6650_,
		_w7026_,
		_w11037_,
		_w11038_
	);
	LUT2 #(
		.INIT('h4)
	) name11005 (
		_w11036_,
		_w11038_,
		_w11039_
	);
	LUT4 #(
		.INIT('h4844)
	) name11006 (
		\a[2] ,
		_w11034_,
		_w11035_,
		_w11039_,
		_w11040_
	);
	LUT4 #(
		.INIT('h2122)
	) name11007 (
		\a[2] ,
		_w11034_,
		_w11035_,
		_w11039_,
		_w11041_
	);
	LUT2 #(
		.INIT('h9)
	) name11008 (
		_w10878_,
		_w10880_,
		_w11042_
	);
	LUT4 #(
		.INIT('h5060)
	) name11009 (
		_w4099_,
		_w4378_,
		_w6334_,
		_w6951_,
		_w11043_
	);
	LUT4 #(
		.INIT('h007b)
	) name11010 (
		_w4030_,
		_w6650_,
		_w6952_,
		_w11043_,
		_w11044_
	);
	LUT3 #(
		.INIT('h70)
	) name11011 (
		_w6657_,
		_w7026_,
		_w11044_,
		_w11045_
	);
	LUT4 #(
		.INIT('h95aa)
	) name11012 (
		\a[2] ,
		_w6335_,
		_w7562_,
		_w11045_,
		_w11046_
	);
	LUT3 #(
		.INIT('h1e)
	) name11013 (
		_w10753_,
		_w10876_,
		_w10877_,
		_w11047_
	);
	LUT3 #(
		.INIT('h82)
	) name11014 (
		_w6335_,
		_w7099_,
		_w7101_,
		_w11048_
	);
	LUT3 #(
		.INIT('h84)
	) name11015 (
		_w4030_,
		_w6657_,
		_w6952_,
		_w11049_
	);
	LUT2 #(
		.INIT('h8)
	) name11016 (
		_w6334_,
		_w7032_,
		_w11050_
	);
	LUT4 #(
		.INIT('h5060)
	) name11017 (
		_w4099_,
		_w4378_,
		_w6650_,
		_w6951_,
		_w11051_
	);
	LUT2 #(
		.INIT('h1)
	) name11018 (
		_w11050_,
		_w11051_,
		_w11052_
	);
	LUT2 #(
		.INIT('h4)
	) name11019 (
		_w11049_,
		_w11052_,
		_w11053_
	);
	LUT4 #(
		.INIT('h4844)
	) name11020 (
		\a[2] ,
		_w11047_,
		_w11048_,
		_w11053_,
		_w11054_
	);
	LUT4 #(
		.INIT('h2122)
	) name11021 (
		\a[2] ,
		_w11047_,
		_w11048_,
		_w11053_,
		_w11055_
	);
	LUT4 #(
		.INIT('h54ab)
	) name11022 (
		_w10759_,
		_w10872_,
		_w10873_,
		_w10875_,
		_w11056_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11023 (
		_w6335_,
		_w7034_,
		_w7097_,
		_w7098_,
		_w11057_
	);
	LUT4 #(
		.INIT('h5060)
	) name11024 (
		_w4099_,
		_w4378_,
		_w6657_,
		_w6951_,
		_w11058_
	);
	LUT3 #(
		.INIT('h82)
	) name11025 (
		_w6334_,
		_w6947_,
		_w6949_,
		_w11059_
	);
	LUT3 #(
		.INIT('h07)
	) name11026 (
		_w6650_,
		_w7032_,
		_w11059_,
		_w11060_
	);
	LUT2 #(
		.INIT('h4)
	) name11027 (
		_w11058_,
		_w11060_,
		_w11061_
	);
	LUT4 #(
		.INIT('h4844)
	) name11028 (
		\a[2] ,
		_w11056_,
		_w11057_,
		_w11061_,
		_w11062_
	);
	LUT4 #(
		.INIT('h2122)
	) name11029 (
		\a[2] ,
		_w11056_,
		_w11057_,
		_w11061_,
		_w11063_
	);
	LUT2 #(
		.INIT('h9)
	) name11030 (
		_w10872_,
		_w10874_,
		_w11064_
	);
	LUT4 #(
		.INIT('h04c8)
	) name11031 (
		_w4695_,
		_w6334_,
		_w6944_,
		_w6946_,
		_w11065_
	);
	LUT4 #(
		.INIT('h007d)
	) name11032 (
		_w6650_,
		_w6947_,
		_w6949_,
		_w11065_,
		_w11066_
	);
	LUT3 #(
		.INIT('h70)
	) name11033 (
		_w6657_,
		_w7032_,
		_w11066_,
		_w11067_
	);
	LUT4 #(
		.INIT('h6a55)
	) name11034 (
		\a[2] ,
		_w6335_,
		_w7882_,
		_w11067_,
		_w11068_
	);
	LUT3 #(
		.INIT('h82)
	) name11035 (
		_w6335_,
		_w7093_,
		_w7095_,
		_w11069_
	);
	LUT3 #(
		.INIT('h82)
	) name11036 (
		_w6657_,
		_w6947_,
		_w6949_,
		_w11070_
	);
	LUT2 #(
		.INIT('h8)
	) name11037 (
		_w6334_,
		_w7038_,
		_w11071_
	);
	LUT4 #(
		.INIT('h04c8)
	) name11038 (
		_w4695_,
		_w6650_,
		_w6944_,
		_w6946_,
		_w11072_
	);
	LUT2 #(
		.INIT('h1)
	) name11039 (
		_w11071_,
		_w11072_,
		_w11073_
	);
	LUT2 #(
		.INIT('h4)
	) name11040 (
		_w11070_,
		_w11073_,
		_w11074_
	);
	LUT3 #(
		.INIT('h9a)
	) name11041 (
		\a[2] ,
		_w11069_,
		_w11074_,
		_w11075_
	);
	LUT3 #(
		.INIT('h1e)
	) name11042 (
		_w10774_,
		_w10870_,
		_w10871_,
		_w11076_
	);
	LUT4 #(
		.INIT('h54ab)
	) name11043 (
		_w10780_,
		_w10866_,
		_w10867_,
		_w10869_,
		_w11077_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11044 (
		_w6335_,
		_w7040_,
		_w7091_,
		_w7092_,
		_w11078_
	);
	LUT4 #(
		.INIT('h04c8)
	) name11045 (
		_w4695_,
		_w6657_,
		_w6944_,
		_w6946_,
		_w11079_
	);
	LUT3 #(
		.INIT('h82)
	) name11046 (
		_w6334_,
		_w6940_,
		_w6942_,
		_w11080_
	);
	LUT3 #(
		.INIT('h07)
	) name11047 (
		_w6650_,
		_w7038_,
		_w11080_,
		_w11081_
	);
	LUT2 #(
		.INIT('h4)
	) name11048 (
		_w11079_,
		_w11081_,
		_w11082_
	);
	LUT4 #(
		.INIT('h4844)
	) name11049 (
		\a[2] ,
		_w11077_,
		_w11078_,
		_w11082_,
		_w11083_
	);
	LUT4 #(
		.INIT('h2122)
	) name11050 (
		\a[2] ,
		_w11077_,
		_w11078_,
		_w11082_,
		_w11084_
	);
	LUT4 #(
		.INIT('h5060)
	) name11051 (
		_w5067_,
		_w5282_,
		_w6334_,
		_w6939_,
		_w11085_
	);
	LUT4 #(
		.INIT('h007d)
	) name11052 (
		_w6650_,
		_w6940_,
		_w6942_,
		_w11085_,
		_w11086_
	);
	LUT3 #(
		.INIT('h70)
	) name11053 (
		_w6657_,
		_w7038_,
		_w11086_,
		_w11087_
	);
	LUT4 #(
		.INIT('h95aa)
	) name11054 (
		\a[2] ,
		_w6335_,
		_w8018_,
		_w11087_,
		_w11088_
	);
	LUT2 #(
		.INIT('h9)
	) name11055 (
		_w10866_,
		_w10868_,
		_w11089_
	);
	LUT3 #(
		.INIT('h1e)
	) name11056 (
		_w10795_,
		_w10864_,
		_w10865_,
		_w11090_
	);
	LUT3 #(
		.INIT('h82)
	) name11057 (
		_w6335_,
		_w7087_,
		_w7089_,
		_w11091_
	);
	LUT3 #(
		.INIT('h82)
	) name11058 (
		_w6657_,
		_w6940_,
		_w6942_,
		_w11092_
	);
	LUT2 #(
		.INIT('h8)
	) name11059 (
		_w6334_,
		_w7044_,
		_w11093_
	);
	LUT4 #(
		.INIT('h5060)
	) name11060 (
		_w5067_,
		_w5282_,
		_w6650_,
		_w6939_,
		_w11094_
	);
	LUT2 #(
		.INIT('h1)
	) name11061 (
		_w11093_,
		_w11094_,
		_w11095_
	);
	LUT2 #(
		.INIT('h4)
	) name11062 (
		_w11092_,
		_w11095_,
		_w11096_
	);
	LUT4 #(
		.INIT('h4844)
	) name11063 (
		\a[2] ,
		_w11090_,
		_w11091_,
		_w11096_,
		_w11097_
	);
	LUT4 #(
		.INIT('h2122)
	) name11064 (
		\a[2] ,
		_w11090_,
		_w11091_,
		_w11096_,
		_w11098_
	);
	LUT4 #(
		.INIT('h54ab)
	) name11065 (
		_w10801_,
		_w10860_,
		_w10861_,
		_w10863_,
		_w11099_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11066 (
		_w6335_,
		_w7046_,
		_w7085_,
		_w7086_,
		_w11100_
	);
	LUT4 #(
		.INIT('h5060)
	) name11067 (
		_w5067_,
		_w5282_,
		_w6657_,
		_w6939_,
		_w11101_
	);
	LUT3 #(
		.INIT('h82)
	) name11068 (
		_w6334_,
		_w6935_,
		_w6937_,
		_w11102_
	);
	LUT3 #(
		.INIT('h07)
	) name11069 (
		_w6650_,
		_w7044_,
		_w11102_,
		_w11103_
	);
	LUT2 #(
		.INIT('h4)
	) name11070 (
		_w11101_,
		_w11103_,
		_w11104_
	);
	LUT4 #(
		.INIT('h4844)
	) name11071 (
		\a[2] ,
		_w11099_,
		_w11100_,
		_w11104_,
		_w11105_
	);
	LUT4 #(
		.INIT('h2122)
	) name11072 (
		\a[2] ,
		_w11099_,
		_w11100_,
		_w11104_,
		_w11106_
	);
	LUT2 #(
		.INIT('h9)
	) name11073 (
		_w10860_,
		_w10862_,
		_w11107_
	);
	LUT4 #(
		.INIT('h04c8)
	) name11074 (
		_w6043_,
		_w6334_,
		_w6933_,
		_w6934_,
		_w11108_
	);
	LUT4 #(
		.INIT('h007d)
	) name11075 (
		_w6650_,
		_w6935_,
		_w6937_,
		_w11108_,
		_w11109_
	);
	LUT3 #(
		.INIT('h70)
	) name11076 (
		_w6657_,
		_w7044_,
		_w11109_,
		_w11110_
	);
	LUT4 #(
		.INIT('h6a55)
	) name11077 (
		\a[2] ,
		_w6335_,
		_w8005_,
		_w11110_,
		_w11111_
	);
	LUT3 #(
		.INIT('h1e)
	) name11078 (
		_w10816_,
		_w10858_,
		_w10859_,
		_w11112_
	);
	LUT3 #(
		.INIT('h82)
	) name11079 (
		_w6335_,
		_w7081_,
		_w7083_,
		_w11113_
	);
	LUT3 #(
		.INIT('h82)
	) name11080 (
		_w6657_,
		_w6935_,
		_w6937_,
		_w11114_
	);
	LUT2 #(
		.INIT('h8)
	) name11081 (
		_w6334_,
		_w7050_,
		_w11115_
	);
	LUT4 #(
		.INIT('h04c8)
	) name11082 (
		_w6043_,
		_w6650_,
		_w6933_,
		_w6934_,
		_w11116_
	);
	LUT2 #(
		.INIT('h1)
	) name11083 (
		_w11115_,
		_w11116_,
		_w11117_
	);
	LUT2 #(
		.INIT('h4)
	) name11084 (
		_w11114_,
		_w11117_,
		_w11118_
	);
	LUT4 #(
		.INIT('h4844)
	) name11085 (
		\a[2] ,
		_w11112_,
		_w11113_,
		_w11118_,
		_w11119_
	);
	LUT4 #(
		.INIT('h2122)
	) name11086 (
		\a[2] ,
		_w11112_,
		_w11113_,
		_w11118_,
		_w11120_
	);
	LUT4 #(
		.INIT('h54ab)
	) name11087 (
		_w10823_,
		_w10854_,
		_w10855_,
		_w10857_,
		_w11121_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11088 (
		_w6335_,
		_w7052_,
		_w7079_,
		_w7080_,
		_w11122_
	);
	LUT4 #(
		.INIT('h04c8)
	) name11089 (
		_w6043_,
		_w6657_,
		_w6933_,
		_w6934_,
		_w11123_
	);
	LUT3 #(
		.INIT('h82)
	) name11090 (
		_w6334_,
		_w6929_,
		_w6931_,
		_w11124_
	);
	LUT3 #(
		.INIT('h07)
	) name11091 (
		_w6650_,
		_w7050_,
		_w11124_,
		_w11125_
	);
	LUT2 #(
		.INIT('h4)
	) name11092 (
		_w11123_,
		_w11125_,
		_w11126_
	);
	LUT4 #(
		.INIT('h4844)
	) name11093 (
		\a[2] ,
		_w11121_,
		_w11122_,
		_w11126_,
		_w11127_
	);
	LUT4 #(
		.INIT('h2122)
	) name11094 (
		\a[2] ,
		_w11121_,
		_w11122_,
		_w11126_,
		_w11128_
	);
	LUT2 #(
		.INIT('h9)
	) name11095 (
		_w10854_,
		_w10856_,
		_w11129_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11096 (
		_w6334_,
		_w6645_,
		_w6926_,
		_w6928_,
		_w11130_
	);
	LUT4 #(
		.INIT('h007d)
	) name11097 (
		_w6650_,
		_w6929_,
		_w6931_,
		_w11130_,
		_w11131_
	);
	LUT3 #(
		.INIT('h70)
	) name11098 (
		_w6657_,
		_w7050_,
		_w11131_,
		_w11132_
	);
	LUT4 #(
		.INIT('h95aa)
	) name11099 (
		\a[2] ,
		_w6335_,
		_w8227_,
		_w11132_,
		_w11133_
	);
	LUT2 #(
		.INIT('h9)
	) name11100 (
		_w10851_,
		_w10853_,
		_w11134_
	);
	LUT3 #(
		.INIT('h82)
	) name11101 (
		_w6335_,
		_w7075_,
		_w7077_,
		_w11135_
	);
	LUT3 #(
		.INIT('h82)
	) name11102 (
		_w6657_,
		_w6929_,
		_w6931_,
		_w11136_
	);
	LUT2 #(
		.INIT('h8)
	) name11103 (
		_w6334_,
		_w7056_,
		_w11137_
	);
	LUT4 #(
		.INIT('h04c8)
	) name11104 (
		_w6645_,
		_w6650_,
		_w6926_,
		_w6928_,
		_w11138_
	);
	LUT2 #(
		.INIT('h1)
	) name11105 (
		_w11137_,
		_w11138_,
		_w11139_
	);
	LUT2 #(
		.INIT('h4)
	) name11106 (
		_w11136_,
		_w11139_,
		_w11140_
	);
	LUT4 #(
		.INIT('h4844)
	) name11107 (
		\a[2] ,
		_w11134_,
		_w11135_,
		_w11140_,
		_w11141_
	);
	LUT4 #(
		.INIT('h2122)
	) name11108 (
		\a[2] ,
		_w11134_,
		_w11135_,
		_w11140_,
		_w11142_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11109 (
		_w6335_,
		_w7058_,
		_w7073_,
		_w7074_,
		_w11143_
	);
	LUT4 #(
		.INIT('h04c8)
	) name11110 (
		_w6645_,
		_w6657_,
		_w6926_,
		_w6928_,
		_w11144_
	);
	LUT3 #(
		.INIT('h82)
	) name11111 (
		_w6334_,
		_w6922_,
		_w6924_,
		_w11145_
	);
	LUT3 #(
		.INIT('h07)
	) name11112 (
		_w6650_,
		_w7056_,
		_w11145_,
		_w11146_
	);
	LUT2 #(
		.INIT('h4)
	) name11113 (
		_w11144_,
		_w11146_,
		_w11147_
	);
	LUT4 #(
		.INIT('h9a65)
	) name11114 (
		\a[5] ,
		_w10844_,
		_w10848_,
		_w10849_,
		_w11148_
	);
	LUT4 #(
		.INIT('h6500)
	) name11115 (
		\a[2] ,
		_w11143_,
		_w11147_,
		_w11148_,
		_w11149_
	);
	LUT4 #(
		.INIT('h009a)
	) name11116 (
		\a[2] ,
		_w11143_,
		_w11147_,
		_w11148_,
		_w11150_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name11117 (
		\a[5] ,
		_w10836_,
		_w10833_,
		_w10835_,
		_w11151_
	);
	LUT3 #(
		.INIT('h4b)
	) name11118 (
		_w10839_,
		_w10842_,
		_w11151_,
		_w11152_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11119 (
		_w6334_,
		_w6669_,
		_w6919_,
		_w6921_,
		_w11153_
	);
	LUT4 #(
		.INIT('h007d)
	) name11120 (
		_w6650_,
		_w6922_,
		_w6924_,
		_w11153_,
		_w11154_
	);
	LUT3 #(
		.INIT('h70)
	) name11121 (
		_w6657_,
		_w7056_,
		_w11154_,
		_w11155_
	);
	LUT4 #(
		.INIT('h6a55)
	) name11122 (
		\a[2] ,
		_w6335_,
		_w8298_,
		_w11155_,
		_w11156_
	);
	LUT3 #(
		.INIT('h82)
	) name11123 (
		_w6335_,
		_w7069_,
		_w7071_,
		_w11157_
	);
	LUT3 #(
		.INIT('h82)
	) name11124 (
		_w6657_,
		_w6922_,
		_w6924_,
		_w11158_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11125 (
		_w6650_,
		_w6669_,
		_w6919_,
		_w6921_,
		_w11159_
	);
	LUT2 #(
		.INIT('h8)
	) name11126 (
		_w6334_,
		_w7062_,
		_w11160_
	);
	LUT2 #(
		.INIT('h1)
	) name11127 (
		_w11159_,
		_w11160_,
		_w11161_
	);
	LUT2 #(
		.INIT('h4)
	) name11128 (
		_w11158_,
		_w11161_,
		_w11162_
	);
	LUT3 #(
		.INIT('h9a)
	) name11129 (
		\a[2] ,
		_w11157_,
		_w11162_,
		_w11163_
	);
	LUT3 #(
		.INIT('h28)
	) name11130 (
		_w6335_,
		_w7065_,
		_w7068_,
		_w11164_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11131 (
		_w6657_,
		_w6669_,
		_w6919_,
		_w6921_,
		_w11165_
	);
	LUT3 #(
		.INIT('h82)
	) name11132 (
		_w6334_,
		_w6914_,
		_w6916_,
		_w11166_
	);
	LUT3 #(
		.INIT('h07)
	) name11133 (
		_w6650_,
		_w7062_,
		_w11166_,
		_w11167_
	);
	LUT2 #(
		.INIT('h4)
	) name11134 (
		_w11165_,
		_w11167_,
		_w11168_
	);
	LUT4 #(
		.INIT('h5401)
	) name11135 (
		\a[2] ,
		_w6689_,
		_w6911_,
		_w6913_,
		_w11169_
	);
	LUT3 #(
		.INIT('h0b)
	) name11136 (
		_w11164_,
		_w11168_,
		_w11169_,
		_w11170_
	);
	LUT4 #(
		.INIT('h1441)
	) name11137 (
		_w6333_,
		_w6914_,
		_w6916_,
		_w7067_,
		_w11171_
	);
	LUT4 #(
		.INIT('h060f)
	) name11138 (
		_w6914_,
		_w6916_,
		_w7067_,
		_w10590_,
		_w11172_
	);
	LUT4 #(
		.INIT('h5700)
	) name11139 (
		\a[0] ,
		_w7062_,
		_w11171_,
		_w11172_,
		_w11173_
	);
	LUT2 #(
		.INIT('h1)
	) name11140 (
		_w10836_,
		_w11173_,
		_w11174_
	);
	LUT4 #(
		.INIT('h00ef)
	) name11141 (
		\a[2] ,
		_w11164_,
		_w11168_,
		_w11174_,
		_w11175_
	);
	LUT2 #(
		.INIT('h4)
	) name11142 (
		_w11170_,
		_w11175_,
		_w11176_
	);
	LUT2 #(
		.INIT('h8)
	) name11143 (
		\a[5] ,
		_w10836_,
		_w11177_
	);
	LUT3 #(
		.INIT('h4b)
	) name11144 (
		_w10833_,
		_w10835_,
		_w11177_,
		_w11178_
	);
	LUT3 #(
		.INIT('h2b)
	) name11145 (
		_w11163_,
		_w11176_,
		_w11178_,
		_w11179_
	);
	LUT4 #(
		.INIT('h4054)
	) name11146 (
		_w11150_,
		_w11152_,
		_w11156_,
		_w11179_,
		_w11180_
	);
	LUT4 #(
		.INIT('h4445)
	) name11147 (
		_w11141_,
		_w11142_,
		_w11149_,
		_w11180_,
		_w11181_
	);
	LUT4 #(
		.INIT('h0445)
	) name11148 (
		_w11128_,
		_w11129_,
		_w11133_,
		_w11181_,
		_w11182_
	);
	LUT4 #(
		.INIT('h4445)
	) name11149 (
		_w11119_,
		_w11120_,
		_w11127_,
		_w11182_,
		_w11183_
	);
	LUT4 #(
		.INIT('h4054)
	) name11150 (
		_w11106_,
		_w11107_,
		_w11111_,
		_w11183_,
		_w11184_
	);
	LUT4 #(
		.INIT('h4445)
	) name11151 (
		_w11097_,
		_w11098_,
		_w11105_,
		_w11184_,
		_w11185_
	);
	LUT4 #(
		.INIT('h1051)
	) name11152 (
		_w11084_,
		_w11088_,
		_w11089_,
		_w11185_,
		_w11186_
	);
	LUT4 #(
		.INIT('hef0e)
	) name11153 (
		_w11083_,
		_w11186_,
		_w11075_,
		_w11076_,
		_w11187_
	);
	LUT4 #(
		.INIT('h0e08)
	) name11154 (
		_w11064_,
		_w11068_,
		_w11063_,
		_w11187_,
		_w11188_
	);
	LUT4 #(
		.INIT('h4445)
	) name11155 (
		_w11054_,
		_w11055_,
		_w11062_,
		_w11188_,
		_w11189_
	);
	LUT4 #(
		.INIT('h0445)
	) name11156 (
		_w11041_,
		_w11042_,
		_w11046_,
		_w11189_,
		_w11190_
	);
	LUT4 #(
		.INIT('hef0e)
	) name11157 (
		_w11040_,
		_w11190_,
		_w11032_,
		_w11033_,
		_w11191_
	);
	LUT4 #(
		.INIT('h0115)
	) name11158 (
		_w11020_,
		_w11021_,
		_w11025_,
		_w11191_,
		_w11192_
	);
	LUT4 #(
		.INIT('h4445)
	) name11159 (
		_w11011_,
		_w11012_,
		_w11019_,
		_w11192_,
		_w11193_
	);
	LUT3 #(
		.INIT('h54)
	) name11160 (
		_w11002_,
		_w11003_,
		_w11193_,
		_w11194_
	);
	LUT4 #(
		.INIT('h0445)
	) name11161 (
		_w10996_,
		_w11000_,
		_w11001_,
		_w11193_,
		_w11195_
	);
	LUT4 #(
		.INIT('ha220)
	) name11162 (
		_w10996_,
		_w11000_,
		_w11001_,
		_w11193_,
		_w11196_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11163 (
		_w6335_,
		_w7016_,
		_w7115_,
		_w7116_,
		_w11197_
	);
	LUT4 #(
		.INIT('h04c8)
	) name11164 (
		_w3257_,
		_w6657_,
		_w6964_,
		_w6966_,
		_w11198_
	);
	LUT3 #(
		.INIT('h82)
	) name11165 (
		_w6334_,
		_w6960_,
		_w6962_,
		_w11199_
	);
	LUT3 #(
		.INIT('h07)
	) name11166 (
		_w6650_,
		_w7014_,
		_w11199_,
		_w11200_
	);
	LUT2 #(
		.INIT('h4)
	) name11167 (
		_w11198_,
		_w11200_,
		_w11201_
	);
	LUT3 #(
		.INIT('h9a)
	) name11168 (
		\a[2] ,
		_w11197_,
		_w11201_,
		_w11202_
	);
	LUT3 #(
		.INIT('h45)
	) name11169 (
		_w11195_,
		_w11196_,
		_w11202_,
		_w11203_
	);
	LUT4 #(
		.INIT('h1501)
	) name11170 (
		_w10995_,
		_w10996_,
		_w11194_,
		_w11202_,
		_w11204_
	);
	LUT4 #(
		.INIT('h80a8)
	) name11171 (
		_w10995_,
		_w10996_,
		_w11194_,
		_w11202_,
		_w11205_
	);
	LUT3 #(
		.INIT('h82)
	) name11172 (
		_w6335_,
		_w7117_,
		_w7119_,
		_w11206_
	);
	LUT3 #(
		.INIT('h82)
	) name11173 (
		_w6657_,
		_w6967_,
		_w6969_,
		_w11207_
	);
	LUT2 #(
		.INIT('h8)
	) name11174 (
		_w6334_,
		_w7014_,
		_w11208_
	);
	LUT4 #(
		.INIT('h04c8)
	) name11175 (
		_w3257_,
		_w6650_,
		_w6964_,
		_w6966_,
		_w11209_
	);
	LUT2 #(
		.INIT('h1)
	) name11176 (
		_w11208_,
		_w11209_,
		_w11210_
	);
	LUT2 #(
		.INIT('h4)
	) name11177 (
		_w11207_,
		_w11210_,
		_w11211_
	);
	LUT3 #(
		.INIT('h9a)
	) name11178 (
		\a[2] ,
		_w11206_,
		_w11211_,
		_w11212_
	);
	LUT3 #(
		.INIT('h45)
	) name11179 (
		_w11204_,
		_w11205_,
		_w11212_,
		_w11213_
	);
	LUT4 #(
		.INIT('h80a8)
	) name11180 (
		_w10994_,
		_w10995_,
		_w11203_,
		_w11212_,
		_w11214_
	);
	LUT4 #(
		.INIT('h1501)
	) name11181 (
		_w10994_,
		_w10995_,
		_w11203_,
		_w11212_,
		_w11215_
	);
	LUT4 #(
		.INIT('h04c8)
	) name11182 (
		_w3257_,
		_w6334_,
		_w6964_,
		_w6966_,
		_w11216_
	);
	LUT4 #(
		.INIT('h007d)
	) name11183 (
		_w6650_,
		_w6967_,
		_w6969_,
		_w11216_,
		_w11217_
	);
	LUT3 #(
		.INIT('h70)
	) name11184 (
		_w6657_,
		_w7008_,
		_w11217_,
		_w11218_
	);
	LUT4 #(
		.INIT('h6a55)
	) name11185 (
		\a[2] ,
		_w6335_,
		_w7403_,
		_w11218_,
		_w11219_
	);
	LUT3 #(
		.INIT('h45)
	) name11186 (
		_w11214_,
		_w11215_,
		_w11219_,
		_w11220_
	);
	LUT4 #(
		.INIT('ha880)
	) name11187 (
		_w10993_,
		_w10994_,
		_w11213_,
		_w11219_,
		_w11221_
	);
	LUT4 #(
		.INIT('h0115)
	) name11188 (
		_w10993_,
		_w10994_,
		_w11213_,
		_w11219_,
		_w11222_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11189 (
		_w6335_,
		_w7010_,
		_w7121_,
		_w7122_,
		_w11223_
	);
	LUT4 #(
		.INIT('h04c8)
	) name11190 (
		_w2983_,
		_w6657_,
		_w6972_,
		_w6974_,
		_w11224_
	);
	LUT3 #(
		.INIT('h82)
	) name11191 (
		_w6334_,
		_w6967_,
		_w6969_,
		_w11225_
	);
	LUT3 #(
		.INIT('h07)
	) name11192 (
		_w6650_,
		_w7008_,
		_w11225_,
		_w11226_
	);
	LUT2 #(
		.INIT('h4)
	) name11193 (
		_w11224_,
		_w11226_,
		_w11227_
	);
	LUT3 #(
		.INIT('h65)
	) name11194 (
		\a[2] ,
		_w11223_,
		_w11227_,
		_w11228_
	);
	LUT3 #(
		.INIT('h45)
	) name11195 (
		_w11221_,
		_w11222_,
		_w11228_,
		_w11229_
	);
	LUT4 #(
		.INIT('h8a08)
	) name11196 (
		_w10992_,
		_w10993_,
		_w11220_,
		_w11228_,
		_w11230_
	);
	LUT2 #(
		.INIT('h4)
	) name11197 (
		_w10977_,
		_w10981_,
		_w11231_
	);
	LUT2 #(
		.INIT('h9)
	) name11198 (
		_w10977_,
		_w10981_,
		_w11232_
	);
	LUT4 #(
		.INIT('h5501)
	) name11199 (
		_w10982_,
		_w10991_,
		_w11230_,
		_w11231_,
		_w11233_
	);
	LUT4 #(
		.INIT('h2122)
	) name11200 (
		\a[2] ,
		_w10969_,
		_w10970_,
		_w10974_,
		_w11234_
	);
	LUT4 #(
		.INIT('h9699)
	) name11201 (
		\a[2] ,
		_w10969_,
		_w10970_,
		_w10974_,
		_w11235_
	);
	LUT3 #(
		.INIT('h54)
	) name11202 (
		_w10976_,
		_w11233_,
		_w11234_,
		_w11236_
	);
	LUT4 #(
		.INIT('h9699)
	) name11203 (
		\a[2] ,
		_w10960_,
		_w10961_,
		_w10966_,
		_w11237_
	);
	LUT4 #(
		.INIT('h2b00)
	) name11204 (
		_w10969_,
		_w10975_,
		_w11233_,
		_w11237_,
		_w11238_
	);
	LUT2 #(
		.INIT('h4)
	) name11205 (
		_w10954_,
		_w10958_,
		_w11239_
	);
	LUT2 #(
		.INIT('h9)
	) name11206 (
		_w10954_,
		_w10958_,
		_w11240_
	);
	LUT4 #(
		.INIT('h5501)
	) name11207 (
		_w10959_,
		_w10968_,
		_w11238_,
		_w11239_,
		_w11241_
	);
	LUT4 #(
		.INIT('h2122)
	) name11208 (
		\a[2] ,
		_w10946_,
		_w10947_,
		_w10951_,
		_w11242_
	);
	LUT4 #(
		.INIT('h9699)
	) name11209 (
		\a[2] ,
		_w10946_,
		_w10947_,
		_w10951_,
		_w11243_
	);
	LUT3 #(
		.INIT('h54)
	) name11210 (
		_w10953_,
		_w11241_,
		_w11242_,
		_w11244_
	);
	LUT4 #(
		.INIT('h9699)
	) name11211 (
		\a[2] ,
		_w10937_,
		_w10938_,
		_w10943_,
		_w11245_
	);
	LUT4 #(
		.INIT('h2b00)
	) name11212 (
		_w10946_,
		_w10952_,
		_w11241_,
		_w11245_,
		_w11246_
	);
	LUT2 #(
		.INIT('h4)
	) name11213 (
		_w10930_,
		_w10935_,
		_w11247_
	);
	LUT2 #(
		.INIT('h9)
	) name11214 (
		_w10930_,
		_w10935_,
		_w11248_
	);
	LUT4 #(
		.INIT('h5501)
	) name11215 (
		_w10936_,
		_w10945_,
		_w11246_,
		_w11247_,
		_w11249_
	);
	LUT4 #(
		.INIT('h2122)
	) name11216 (
		\a[2] ,
		_w10923_,
		_w10924_,
		_w10927_,
		_w11250_
	);
	LUT4 #(
		.INIT('h9699)
	) name11217 (
		\a[2] ,
		_w10923_,
		_w10924_,
		_w10927_,
		_w11251_
	);
	LUT4 #(
		.INIT('h088a)
	) name11218 (
		_w10922_,
		_w10923_,
		_w10928_,
		_w11249_,
		_w11252_
	);
	LUT2 #(
		.INIT('h1)
	) name11219 (
		_w10921_,
		_w11252_,
		_w11253_
	);
	LUT3 #(
		.INIT('h54)
	) name11220 (
		_w10597_,
		_w10598_,
		_w11253_,
		_w11254_
	);
	LUT3 #(
		.INIT('h54)
	) name11221 (
		_w10578_,
		_w10579_,
		_w11254_,
		_w11255_
	);
	LUT3 #(
		.INIT('h54)
	) name11222 (
		_w10266_,
		_w10267_,
		_w11255_,
		_w11256_
	);
	LUT2 #(
		.INIT('h4)
	) name11223 (
		_w9703_,
		_w9975_,
		_w11257_
	);
	LUT2 #(
		.INIT('h9)
	) name11224 (
		_w9703_,
		_w9975_,
		_w11258_
	);
	LUT3 #(
		.INIT('h54)
	) name11225 (
		_w9976_,
		_w11256_,
		_w11257_,
		_w11259_
	);
	LUT3 #(
		.INIT('h96)
	) name11226 (
		_w9443_,
		_w9700_,
		_w9701_,
		_w11260_
	);
	LUT4 #(
		.INIT('h2b00)
	) name11227 (
		_w9703_,
		_w9975_,
		_w11256_,
		_w11260_,
		_w11261_
	);
	LUT4 #(
		.INIT('h1115)
	) name11228 (
		_w9445_,
		_w9446_,
		_w9702_,
		_w11261_,
		_w11262_
	);
	LUT3 #(
		.INIT('h90)
	) name11229 (
		_w8989_,
		_w8991_,
		_w9211_,
		_w11263_
	);
	LUT3 #(
		.INIT('h69)
	) name11230 (
		_w8989_,
		_w8991_,
		_w9211_,
		_w11264_
	);
	LUT3 #(
		.INIT('h54)
	) name11231 (
		_w9212_,
		_w11262_,
		_w11263_,
		_w11265_
	);
	LUT2 #(
		.INIT('h6)
	) name11232 (
		_w8992_,
		_w8993_,
		_w11266_
	);
	LUT4 #(
		.INIT('hba00)
	) name11233 (
		_w9212_,
		_w11262_,
		_w11264_,
		_w11266_,
		_w11267_
	);
	LUT4 #(
		.INIT('h4445)
	) name11234 (
		_w8792_,
		_w8793_,
		_w8994_,
		_w11267_,
		_w11268_
	);
	LUT2 #(
		.INIT('h4)
	) name11235 (
		_w8542_,
		_w8615_,
		_w11269_
	);
	LUT2 #(
		.INIT('h9)
	) name11236 (
		_w8542_,
		_w8615_,
		_w11270_
	);
	LUT3 #(
		.INIT('h54)
	) name11237 (
		_w8616_,
		_w11268_,
		_w11269_,
		_w11271_
	);
	LUT2 #(
		.INIT('h9)
	) name11238 (
		_w8539_,
		_w8540_,
		_w11272_
	);
	LUT4 #(
		.INIT('h2b00)
	) name11239 (
		_w8542_,
		_w8615_,
		_w11268_,
		_w11272_,
		_w11273_
	);
	LUT4 #(
		.INIT('h4445)
	) name11240 (
		_w8464_,
		_w8465_,
		_w8541_,
		_w11273_,
		_w11274_
	);
	LUT4 #(
		.INIT('h4054)
	) name11241 (
		_w8078_,
		_w8084_,
		_w8145_,
		_w8148_,
		_w11275_
	);
	LUT4 #(
		.INIT('h6566)
	) name11242 (
		_w8078_,
		_w8146_,
		_w8147_,
		_w8148_,
		_w11276_
	);
	LUT3 #(
		.INIT('h54)
	) name11243 (
		_w8150_,
		_w11274_,
		_w11275_,
		_w11277_
	);
	LUT4 #(
		.INIT('hae51)
	) name11244 (
		_w8072_,
		_w8073_,
		_w8074_,
		_w8076_,
		_w11278_
	);
	LUT4 #(
		.INIT('h2b00)
	) name11245 (
		_w8078_,
		_w8149_,
		_w11274_,
		_w11278_,
		_w11279_
	);
	LUT4 #(
		.INIT('h4445)
	) name11246 (
		_w7933_,
		_w7934_,
		_w8077_,
		_w11279_,
		_w11280_
	);
	LUT2 #(
		.INIT('h4)
	) name11247 (
		_w7751_,
		_w7815_,
		_w11281_
	);
	LUT2 #(
		.INIT('h9)
	) name11248 (
		_w7751_,
		_w7815_,
		_w11282_
	);
	LUT3 #(
		.INIT('h54)
	) name11249 (
		_w7816_,
		_w11280_,
		_w11281_,
		_w11283_
	);
	LUT4 #(
		.INIT('hae51)
	) name11250 (
		_w7744_,
		_w7745_,
		_w7746_,
		_w7749_,
		_w11284_
	);
	LUT4 #(
		.INIT('h2b00)
	) name11251 (
		_w7751_,
		_w7815_,
		_w11280_,
		_w11284_,
		_w11285_
	);
	LUT4 #(
		.INIT('h4445)
	) name11252 (
		_w7693_,
		_w7694_,
		_w7750_,
		_w11285_,
		_w11286_
	);
	LUT3 #(
		.INIT('hd4)
	) name11253 (
		_w7376_,
		_w7383_,
		_w7186_,
		_w11287_
	);
	LUT4 #(
		.INIT('h04c8)
	) name11254 (
		_w2622_,
		_w2874_,
		_w6978_,
		_w6980_,
		_w11288_
	);
	LUT4 #(
		.INIT('h007b)
	) name11255 (
		_w2546_,
		_w2975_,
		_w6981_,
		_w11288_,
		_w11289_
	);
	LUT3 #(
		.INIT('h70)
	) name11256 (
		_w2986_,
		_w6996_,
		_w11289_,
		_w11290_
	);
	LUT4 #(
		.INIT('h95aa)
	) name11257 (
		\a[26] ,
		_w2875_,
		_w7500_,
		_w11290_,
		_w11291_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11258 (
		_w2549_,
		_w2983_,
		_w6972_,
		_w6974_,
		_w11292_
	);
	LUT4 #(
		.INIT('h007d)
	) name11259 (
		_w2617_,
		_w2872_,
		_w6975_,
		_w11292_,
		_w11293_
	);
	LUT3 #(
		.INIT('h70)
	) name11260 (
		_w2854_,
		_w7002_,
		_w11293_,
		_w11294_
	);
	LUT4 #(
		.INIT('h95aa)
	) name11261 (
		\a[29] ,
		_w2550_,
		_w7426_,
		_w11294_,
		_w11295_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11262 (
		_w376_,
		_w3257_,
		_w6964_,
		_w6966_,
		_w11296_
	);
	LUT4 #(
		.INIT('h007d)
	) name11263 (
		_w2407_,
		_w6967_,
		_w6969_,
		_w11296_,
		_w11297_
	);
	LUT3 #(
		.INIT('h70)
	) name11264 (
		_w2527_,
		_w7008_,
		_w11297_,
		_w11298_
	);
	LUT3 #(
		.INIT('h70)
	) name11265 (
		_w377_,
		_w7403_,
		_w11298_,
		_w11299_
	);
	LUT4 #(
		.INIT('h4544)
	) name11266 (
		_w7279_,
		_w7280_,
		_w7282_,
		_w7287_,
		_w11300_
	);
	LUT4 #(
		.INIT('h8001)
	) name11267 (
		\a[17] ,
		\a[18] ,
		\a[19] ,
		\a[20] ,
		_w11301_
	);
	LUT4 #(
		.INIT('h559a)
	) name11268 (
		\a[20] ,
		_w7136_,
		_w7166_,
		_w11301_,
		_w11302_
	);
	LUT3 #(
		.INIT('h80)
	) name11269 (
		_w1774_,
		_w3447_,
		_w7318_,
		_w11303_
	);
	LUT3 #(
		.INIT('h80)
	) name11270 (
		_w674_,
		_w2159_,
		_w11303_,
		_w11304_
	);
	LUT2 #(
		.INIT('h8)
	) name11271 (
		_w974_,
		_w1401_,
		_w11305_
	);
	LUT4 #(
		.INIT('h2000)
	) name11272 (
		_w401_,
		_w389_,
		_w964_,
		_w942_,
		_w11306_
	);
	LUT4 #(
		.INIT('h8000)
	) name11273 (
		_w1465_,
		_w1467_,
		_w11305_,
		_w11306_,
		_w11307_
	);
	LUT3 #(
		.INIT('h80)
	) name11274 (
		_w1156_,
		_w1221_,
		_w2644_,
		_w11308_
	);
	LUT4 #(
		.INIT('h0777)
	) name11275 (
		_w106_,
		_w85_,
		_w56_,
		_w43_,
		_w11309_
	);
	LUT4 #(
		.INIT('h8000)
	) name11276 (
		_w1003_,
		_w1099_,
		_w1079_,
		_w11309_,
		_w11310_
	);
	LUT4 #(
		.INIT('h153f)
	) name11277 (
		_w106_,
		_w59_,
		_w72_,
		_w65_,
		_w11311_
	);
	LUT4 #(
		.INIT('h1000)
	) name11278 (
		_w308_,
		_w398_,
		_w1012_,
		_w11311_,
		_w11312_
	);
	LUT3 #(
		.INIT('h80)
	) name11279 (
		_w11308_,
		_w11310_,
		_w11312_,
		_w11313_
	);
	LUT4 #(
		.INIT('h8000)
	) name11280 (
		_w1236_,
		_w1240_,
		_w2247_,
		_w2249_,
		_w11314_
	);
	LUT4 #(
		.INIT('h8000)
	) name11281 (
		_w11304_,
		_w11307_,
		_w11313_,
		_w11314_,
		_w11315_
	);
	LUT2 #(
		.INIT('h8)
	) name11282 (
		_w1686_,
		_w11315_,
		_w11316_
	);
	LUT2 #(
		.INIT('h1)
	) name11283 (
		_w7217_,
		_w11316_,
		_w11317_
	);
	LUT2 #(
		.INIT('h8)
	) name11284 (
		_w7217_,
		_w11316_,
		_w11318_
	);
	LUT2 #(
		.INIT('h6)
	) name11285 (
		_w7217_,
		_w11316_,
		_w11319_
	);
	LUT4 #(
		.INIT('h6996)
	) name11286 (
		_w11302_,
		_w11319_,
		_w11300_,
		_w11299_,
		_w11320_
	);
	LUT4 #(
		.INIT('he11e)
	) name11287 (
		_w7289_,
		_w7375_,
		_w11320_,
		_w11295_,
		_w11321_
	);
	LUT3 #(
		.INIT('h69)
	) name11288 (
		_w11291_,
		_w11321_,
		_w11287_,
		_w11322_
	);
	LUT3 #(
		.INIT('h28)
	) name11289 (
		_w3249_,
		_w7136_,
		_w7168_,
		_w11323_
	);
	LUT4 #(
		.INIT('h028a)
	) name11290 (
		_w3262_,
		_w7136_,
		_w7166_,
		_w7167_,
		_w11324_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11291 (
		_w3214_,
		_w2411_,
		_w6983_,
		_w6993_,
		_w11325_
	);
	LUT3 #(
		.INIT('h01)
	) name11292 (
		_w11324_,
		_w11325_,
		_w11323_,
		_w11326_
	);
	LUT4 #(
		.INIT('h95aa)
	) name11293 (
		\a[23] ,
		_w37_,
		_w7696_,
		_w11326_,
		_w11327_
	);
	LUT4 #(
		.INIT('h0445)
	) name11294 (
		_w11327_,
		_w7384_,
		_w7415_,
		_w7179_,
		_w11328_
	);
	LUT4 #(
		.INIT('ha220)
	) name11295 (
		_w11327_,
		_w7384_,
		_w7415_,
		_w7179_,
		_w11329_
	);
	LUT4 #(
		.INIT('h599a)
	) name11296 (
		_w11327_,
		_w7384_,
		_w7415_,
		_w7179_,
		_w11330_
	);
	LUT2 #(
		.INIT('h6)
	) name11297 (
		_w11322_,
		_w11330_,
		_w11331_
	);
	LUT3 #(
		.INIT('h54)
	) name11298 (
		_w7496_,
		_w7497_,
		_w7416_,
		_w11332_
	);
	LUT2 #(
		.INIT('h2)
	) name11299 (
		_w11331_,
		_w11332_,
		_w11333_
	);
	LUT2 #(
		.INIT('h4)
	) name11300 (
		_w11331_,
		_w11332_,
		_w11334_
	);
	LUT2 #(
		.INIT('h9)
	) name11301 (
		_w11331_,
		_w11332_,
		_w11335_
	);
	LUT3 #(
		.INIT('h54)
	) name11302 (
		_w11333_,
		_w11286_,
		_w11334_,
		_w11336_
	);
	LUT3 #(
		.INIT('h51)
	) name11303 (
		_w11328_,
		_w11322_,
		_w11329_,
		_w11337_
	);
	LUT4 #(
		.INIT('h0a02)
	) name11304 (
		_w37_,
		_w7169_,
		_w7419_,
		_w7686_,
		_w11338_
	);
	LUT3 #(
		.INIT('h28)
	) name11305 (
		_w3214_,
		_w7136_,
		_w7168_,
		_w11339_
	);
	LUT4 #(
		.INIT('h781e)
	) name11306 (
		\a[20] ,
		\a[21] ,
		\a[22] ,
		\a[23] ,
		_w11340_
	);
	LUT3 #(
		.INIT('hb0)
	) name11307 (
		_w7136_,
		_w7166_,
		_w11340_,
		_w11341_
	);
	LUT3 #(
		.INIT('h40)
	) name11308 (
		_w3262_,
		_w7136_,
		_w7167_,
		_w11342_
	);
	LUT3 #(
		.INIT('h31)
	) name11309 (
		_w11341_,
		_w11339_,
		_w11342_,
		_w11343_
	);
	LUT3 #(
		.INIT('h9a)
	) name11310 (
		\a[23] ,
		_w11338_,
		_w11343_,
		_w11344_
	);
	LUT3 #(
		.INIT('he8)
	) name11311 (
		_w11291_,
		_w11321_,
		_w11287_,
		_w11345_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11312 (
		_w2875_,
		_w6998_,
		_w7133_,
		_w7134_,
		_w11346_
	);
	LUT4 #(
		.INIT('h04c8)
	) name11313 (
		_w2411_,
		_w2986_,
		_w6983_,
		_w6993_,
		_w11347_
	);
	LUT3 #(
		.INIT('h84)
	) name11314 (
		_w2546_,
		_w2874_,
		_w6981_,
		_w11348_
	);
	LUT3 #(
		.INIT('h07)
	) name11315 (
		_w2975_,
		_w6996_,
		_w11348_,
		_w11349_
	);
	LUT2 #(
		.INIT('h4)
	) name11316 (
		_w11347_,
		_w11349_,
		_w11350_
	);
	LUT3 #(
		.INIT('h9a)
	) name11317 (
		\a[26] ,
		_w11346_,
		_w11350_,
		_w11351_
	);
	LUT3 #(
		.INIT('h51)
	) name11318 (
		_w11317_,
		_w11302_,
		_w11318_,
		_w11352_
	);
	LUT4 #(
		.INIT('h2a02)
	) name11319 (
		_w7148_,
		_w7217_,
		_w11316_,
		_w11302_,
		_w11353_
	);
	LUT4 #(
		.INIT('h4054)
	) name11320 (
		_w7148_,
		_w7217_,
		_w11316_,
		_w11302_,
		_w11354_
	);
	LUT4 #(
		.INIT('h6656)
	) name11321 (
		_w7148_,
		_w11317_,
		_w11302_,
		_w11318_,
		_w11355_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11322 (
		_w377_,
		_w7010_,
		_w7121_,
		_w7122_,
		_w11356_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11323 (
		_w2527_,
		_w2983_,
		_w6972_,
		_w6974_,
		_w11357_
	);
	LUT3 #(
		.INIT('h82)
	) name11324 (
		_w376_,
		_w6967_,
		_w6969_,
		_w11358_
	);
	LUT3 #(
		.INIT('h07)
	) name11325 (
		_w2407_,
		_w7008_,
		_w11358_,
		_w11359_
	);
	LUT2 #(
		.INIT('h4)
	) name11326 (
		_w11357_,
		_w11359_,
		_w11360_
	);
	LUT2 #(
		.INIT('h4)
	) name11327 (
		_w11356_,
		_w11360_,
		_w11361_
	);
	LUT4 #(
		.INIT('h066f)
	) name11328 (
		_w11302_,
		_w11319_,
		_w11300_,
		_w11299_,
		_w11362_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11329 (
		_w2550_,
		_w7004_,
		_w7127_,
		_w7128_,
		_w11363_
	);
	LUT4 #(
		.INIT('h04c8)
	) name11330 (
		_w2622_,
		_w2854_,
		_w6978_,
		_w6980_,
		_w11364_
	);
	LUT3 #(
		.INIT('h82)
	) name11331 (
		_w2549_,
		_w2872_,
		_w6975_,
		_w11365_
	);
	LUT3 #(
		.INIT('h07)
	) name11332 (
		_w2617_,
		_w7002_,
		_w11365_,
		_w11366_
	);
	LUT2 #(
		.INIT('h4)
	) name11333 (
		_w11364_,
		_w11366_,
		_w11367_
	);
	LUT3 #(
		.INIT('h9a)
	) name11334 (
		\a[29] ,
		_w11363_,
		_w11367_,
		_w11368_
	);
	LUT4 #(
		.INIT('h6996)
	) name11335 (
		_w11355_,
		_w11361_,
		_w11362_,
		_w11368_,
		_w11369_
	);
	LUT4 #(
		.INIT('h1f01)
	) name11336 (
		_w7289_,
		_w7375_,
		_w11320_,
		_w11295_,
		_w11370_
	);
	LUT3 #(
		.INIT('h69)
	) name11337 (
		_w11369_,
		_w11370_,
		_w11351_,
		_w11371_
	);
	LUT3 #(
		.INIT('h69)
	) name11338 (
		_w11345_,
		_w11371_,
		_w11344_,
		_w11372_
	);
	LUT2 #(
		.INIT('h4)
	) name11339 (
		_w11337_,
		_w11372_,
		_w11373_
	);
	LUT2 #(
		.INIT('h9)
	) name11340 (
		_w11337_,
		_w11372_,
		_w11374_
	);
	LUT4 #(
		.INIT('h2b00)
	) name11341 (
		_w11331_,
		_w11332_,
		_w11286_,
		_w11374_,
		_w11375_
	);
	LUT4 #(
		.INIT('h00d4)
	) name11342 (
		_w11331_,
		_w11332_,
		_w11286_,
		_w11374_,
		_w11376_
	);
	LUT4 #(
		.INIT('h54ab)
	) name11343 (
		_w11333_,
		_w11286_,
		_w11334_,
		_w11374_,
		_w11377_
	);
	LUT4 #(
		.INIT('h1422)
	) name11344 (
		_w11333_,
		_w11286_,
		_w11334_,
		_w11374_,
		_w11378_
	);
	LUT3 #(
		.INIT('h56)
	) name11345 (
		_w7695_,
		_w7750_,
		_w11285_,
		_w11379_
	);
	LUT3 #(
		.INIT('h90)
	) name11346 (
		_w11286_,
		_w11335_,
		_w11379_,
		_w11380_
	);
	LUT4 #(
		.INIT('h00d4)
	) name11347 (
		_w7751_,
		_w7815_,
		_w11280_,
		_w11284_,
		_w11381_
	);
	LUT4 #(
		.INIT('h54ab)
	) name11348 (
		_w7816_,
		_w11280_,
		_w11281_,
		_w11284_,
		_w11382_
	);
	LUT4 #(
		.INIT('h2881)
	) name11349 (
		_w7695_,
		_w7748_,
		_w7749_,
		_w11283_,
		_w11383_
	);
	LUT4 #(
		.INIT('h9402)
	) name11350 (
		_w7751_,
		_w7815_,
		_w11280_,
		_w11284_,
		_w11384_
	);
	LUT3 #(
		.INIT('h56)
	) name11351 (
		_w7935_,
		_w8077_,
		_w11279_,
		_w11385_
	);
	LUT3 #(
		.INIT('h90)
	) name11352 (
		_w11280_,
		_w11282_,
		_w11385_,
		_w11386_
	);
	LUT4 #(
		.INIT('h00d4)
	) name11353 (
		_w8078_,
		_w8149_,
		_w11274_,
		_w11278_,
		_w11387_
	);
	LUT4 #(
		.INIT('h54ab)
	) name11354 (
		_w8150_,
		_w11274_,
		_w11275_,
		_w11278_,
		_w11388_
	);
	LUT4 #(
		.INIT('h6006)
	) name11355 (
		_w7935_,
		_w8077_,
		_w11277_,
		_w11278_,
		_w11389_
	);
	LUT4 #(
		.INIT('h9402)
	) name11356 (
		_w8078_,
		_w8149_,
		_w11274_,
		_w11278_,
		_w11390_
	);
	LUT3 #(
		.INIT('h56)
	) name11357 (
		_w8466_,
		_w8541_,
		_w11273_,
		_w11391_
	);
	LUT3 #(
		.INIT('h90)
	) name11358 (
		_w11274_,
		_w11276_,
		_w11391_,
		_w11392_
	);
	LUT4 #(
		.INIT('h00d4)
	) name11359 (
		_w8542_,
		_w8615_,
		_w11268_,
		_w11272_,
		_w11393_
	);
	LUT4 #(
		.INIT('h54ab)
	) name11360 (
		_w8616_,
		_w11268_,
		_w11269_,
		_w11272_,
		_w11394_
	);
	LUT4 #(
		.INIT('h8218)
	) name11361 (
		_w8466_,
		_w8539_,
		_w8540_,
		_w11271_,
		_w11395_
	);
	LUT4 #(
		.INIT('h9402)
	) name11362 (
		_w8542_,
		_w8615_,
		_w11268_,
		_w11272_,
		_w11396_
	);
	LUT3 #(
		.INIT('h56)
	) name11363 (
		_w8794_,
		_w8994_,
		_w11267_,
		_w11397_
	);
	LUT3 #(
		.INIT('h90)
	) name11364 (
		_w11268_,
		_w11270_,
		_w11397_,
		_w11398_
	);
	LUT4 #(
		.INIT('h0045)
	) name11365 (
		_w9212_,
		_w11262_,
		_w11264_,
		_w11266_,
		_w11399_
	);
	LUT4 #(
		.INIT('h54ab)
	) name11366 (
		_w9212_,
		_w11262_,
		_w11263_,
		_w11266_,
		_w11400_
	);
	LUT4 #(
		.INIT('h2881)
	) name11367 (
		_w8794_,
		_w8992_,
		_w8993_,
		_w11265_,
		_w11401_
	);
	LUT2 #(
		.INIT('h9)
	) name11368 (
		_w11262_,
		_w11264_,
		_w11402_
	);
	LUT3 #(
		.INIT('h56)
	) name11369 (
		_w9446_,
		_w9702_,
		_w11261_,
		_w11403_
	);
	LUT3 #(
		.INIT('h90)
	) name11370 (
		_w11262_,
		_w11264_,
		_w11403_,
		_w11404_
	);
	LUT4 #(
		.INIT('h00d4)
	) name11371 (
		_w9703_,
		_w9975_,
		_w11256_,
		_w11260_,
		_w11405_
	);
	LUT4 #(
		.INIT('h54ab)
	) name11372 (
		_w9976_,
		_w11256_,
		_w11257_,
		_w11260_,
		_w11406_
	);
	LUT4 #(
		.INIT('h6006)
	) name11373 (
		_w9446_,
		_w9702_,
		_w11259_,
		_w11260_,
		_w11407_
	);
	LUT4 #(
		.INIT('h9402)
	) name11374 (
		_w9703_,
		_w9975_,
		_w11256_,
		_w11260_,
		_w11408_
	);
	LUT2 #(
		.INIT('h9)
	) name11375 (
		_w10268_,
		_w11255_,
		_w11409_
	);
	LUT3 #(
		.INIT('h90)
	) name11376 (
		_w11256_,
		_w11258_,
		_w11409_,
		_w11410_
	);
	LUT2 #(
		.INIT('h9)
	) name11377 (
		_w10580_,
		_w11254_,
		_w11411_
	);
	LUT3 #(
		.INIT('h90)
	) name11378 (
		_w10268_,
		_w11255_,
		_w11411_,
		_w11412_
	);
	LUT2 #(
		.INIT('h9)
	) name11379 (
		_w10599_,
		_w11253_,
		_w11413_
	);
	LUT3 #(
		.INIT('h90)
	) name11380 (
		_w10580_,
		_w11254_,
		_w11413_,
		_w11414_
	);
	LUT4 #(
		.INIT('h6665)
	) name11381 (
		_w10922_,
		_w10929_,
		_w11249_,
		_w11250_,
		_w11415_
	);
	LUT3 #(
		.INIT('h90)
	) name11382 (
		_w10599_,
		_w11253_,
		_w11415_,
		_w11416_
	);
	LUT4 #(
		.INIT('h8224)
	) name11383 (
		_w10922_,
		_w10923_,
		_w10928_,
		_w11249_,
		_w11417_
	);
	LUT3 #(
		.INIT('h1e)
	) name11384 (
		_w10945_,
		_w11246_,
		_w11248_,
		_w11418_
	);
	LUT3 #(
		.INIT('h90)
	) name11385 (
		_w11249_,
		_w11251_,
		_w11418_,
		_w11419_
	);
	LUT4 #(
		.INIT('h00d4)
	) name11386 (
		_w10946_,
		_w10952_,
		_w11241_,
		_w11245_,
		_w11420_
	);
	LUT4 #(
		.INIT('h54ab)
	) name11387 (
		_w10953_,
		_w11241_,
		_w11242_,
		_w11245_,
		_w11421_
	);
	LUT4 #(
		.INIT('h9402)
	) name11388 (
		_w10937_,
		_w10944_,
		_w11244_,
		_w11248_,
		_w11422_
	);
	LUT4 #(
		.INIT('h9402)
	) name11389 (
		_w10946_,
		_w10952_,
		_w11241_,
		_w11245_,
		_w11423_
	);
	LUT3 #(
		.INIT('h1e)
	) name11390 (
		_w10968_,
		_w11238_,
		_w11240_,
		_w11424_
	);
	LUT3 #(
		.INIT('h90)
	) name11391 (
		_w11241_,
		_w11243_,
		_w11424_,
		_w11425_
	);
	LUT4 #(
		.INIT('h00d4)
	) name11392 (
		_w10969_,
		_w10975_,
		_w11233_,
		_w11237_,
		_w11426_
	);
	LUT4 #(
		.INIT('h54ab)
	) name11393 (
		_w10976_,
		_w11233_,
		_w11234_,
		_w11237_,
		_w11427_
	);
	LUT4 #(
		.INIT('h9402)
	) name11394 (
		_w10960_,
		_w10967_,
		_w11236_,
		_w11240_,
		_w11428_
	);
	LUT4 #(
		.INIT('h9402)
	) name11395 (
		_w10969_,
		_w10975_,
		_w11233_,
		_w11237_,
		_w11429_
	);
	LUT4 #(
		.INIT('h2940)
	) name11396 (
		_w10969_,
		_w10975_,
		_w11233_,
		_w11237_,
		_w11430_
	);
	LUT4 #(
		.INIT('h629d)
	) name11397 (
		_w10976_,
		_w11233_,
		_w11234_,
		_w11237_,
		_w11431_
	);
	LUT3 #(
		.INIT('h1e)
	) name11398 (
		_w10991_,
		_w11230_,
		_w11232_,
		_w11432_
	);
	LUT4 #(
		.INIT('h1051)
	) name11399 (
		_w10992_,
		_w10993_,
		_w11220_,
		_w11228_,
		_w11433_
	);
	LUT4 #(
		.INIT('h6566)
	) name11400 (
		_w10992_,
		_w11221_,
		_w11222_,
		_w11228_,
		_w11434_
	);
	LUT4 #(
		.INIT('hf090)
	) name11401 (
		_w11233_,
		_w11235_,
		_w11432_,
		_w11434_,
		_w11435_
	);
	LUT3 #(
		.INIT('h45)
	) name11402 (
		_w11429_,
		_w11430_,
		_w11435_,
		_w11436_
	);
	LUT4 #(
		.INIT('h2940)
	) name11403 (
		_w10960_,
		_w10967_,
		_w11236_,
		_w11240_,
		_w11437_
	);
	LUT4 #(
		.INIT('h1e2d)
	) name11404 (
		_w10968_,
		_w11238_,
		_w11240_,
		_w11426_,
		_w11438_
	);
	LUT3 #(
		.INIT('h54)
	) name11405 (
		_w11428_,
		_w11436_,
		_w11437_,
		_w11439_
	);
	LUT3 #(
		.INIT('h06)
	) name11406 (
		_w11241_,
		_w11243_,
		_w11424_,
		_w11440_
	);
	LUT3 #(
		.INIT('h69)
	) name11407 (
		_w11241_,
		_w11243_,
		_w11424_,
		_w11441_
	);
	LUT4 #(
		.INIT('h629d)
	) name11408 (
		_w10953_,
		_w11241_,
		_w11242_,
		_w11245_,
		_w11442_
	);
	LUT4 #(
		.INIT('hba00)
	) name11409 (
		_w11425_,
		_w11439_,
		_w11441_,
		_w11442_,
		_w11443_
	);
	LUT4 #(
		.INIT('h1e2d)
	) name11410 (
		_w10945_,
		_w11246_,
		_w11248_,
		_w11420_,
		_w11444_
	);
	LUT4 #(
		.INIT('h0155)
	) name11411 (
		_w11422_,
		_w11423_,
		_w11443_,
		_w11444_,
		_w11445_
	);
	LUT3 #(
		.INIT('h06)
	) name11412 (
		_w11249_,
		_w11251_,
		_w11418_,
		_w11446_
	);
	LUT3 #(
		.INIT('h69)
	) name11413 (
		_w11249_,
		_w11251_,
		_w11418_,
		_w11447_
	);
	LUT4 #(
		.INIT('h6959)
	) name11414 (
		_w10922_,
		_w10929_,
		_w11249_,
		_w11250_,
		_w11448_
	);
	LUT4 #(
		.INIT('hba00)
	) name11415 (
		_w11419_,
		_w11445_,
		_w11447_,
		_w11448_,
		_w11449_
	);
	LUT2 #(
		.INIT('h1)
	) name11416 (
		_w11417_,
		_w11449_,
		_w11450_
	);
	LUT3 #(
		.INIT('h06)
	) name11417 (
		_w10599_,
		_w11253_,
		_w11415_,
		_w11451_
	);
	LUT3 #(
		.INIT('h69)
	) name11418 (
		_w10599_,
		_w11253_,
		_w11415_,
		_w11452_
	);
	LUT3 #(
		.INIT('h54)
	) name11419 (
		_w11416_,
		_w11450_,
		_w11451_,
		_w11453_
	);
	LUT3 #(
		.INIT('h06)
	) name11420 (
		_w10580_,
		_w11254_,
		_w11413_,
		_w11454_
	);
	LUT3 #(
		.INIT('h69)
	) name11421 (
		_w10580_,
		_w11254_,
		_w11413_,
		_w11455_
	);
	LUT3 #(
		.INIT('h54)
	) name11422 (
		_w11414_,
		_w11453_,
		_w11454_,
		_w11456_
	);
	LUT3 #(
		.INIT('h06)
	) name11423 (
		_w10268_,
		_w11255_,
		_w11411_,
		_w11457_
	);
	LUT3 #(
		.INIT('h69)
	) name11424 (
		_w10268_,
		_w11255_,
		_w11411_,
		_w11458_
	);
	LUT3 #(
		.INIT('h54)
	) name11425 (
		_w11412_,
		_w11456_,
		_w11457_,
		_w11459_
	);
	LUT3 #(
		.INIT('h06)
	) name11426 (
		_w11256_,
		_w11258_,
		_w11409_,
		_w11460_
	);
	LUT3 #(
		.INIT('h69)
	) name11427 (
		_w11256_,
		_w11258_,
		_w11409_,
		_w11461_
	);
	LUT4 #(
		.INIT('h629d)
	) name11428 (
		_w9976_,
		_w11256_,
		_w11257_,
		_w11260_,
		_w11462_
	);
	LUT4 #(
		.INIT('hba00)
	) name11429 (
		_w11410_,
		_w11459_,
		_w11461_,
		_w11462_,
		_w11463_
	);
	LUT4 #(
		.INIT('h5659)
	) name11430 (
		_w9446_,
		_w9702_,
		_w11261_,
		_w11405_,
		_w11464_
	);
	LUT4 #(
		.INIT('h0155)
	) name11431 (
		_w11407_,
		_w11408_,
		_w11463_,
		_w11464_,
		_w11465_
	);
	LUT3 #(
		.INIT('h06)
	) name11432 (
		_w11262_,
		_w11264_,
		_w11403_,
		_w11466_
	);
	LUT3 #(
		.INIT('h69)
	) name11433 (
		_w11262_,
		_w11264_,
		_w11403_,
		_w11467_
	);
	LUT4 #(
		.INIT('h629d)
	) name11434 (
		_w9212_,
		_w11262_,
		_w11263_,
		_w11266_,
		_w11468_
	);
	LUT4 #(
		.INIT('h3713)
	) name11435 (
		_w11400_,
		_w11402_,
		_w11403_,
		_w11465_,
		_w11469_
	);
	LUT4 #(
		.INIT('h4228)
	) name11436 (
		_w8794_,
		_w8992_,
		_w8993_,
		_w11265_,
		_w11470_
	);
	LUT4 #(
		.INIT('h5659)
	) name11437 (
		_w8794_,
		_w8994_,
		_w11267_,
		_w11399_,
		_w11471_
	);
	LUT3 #(
		.INIT('h54)
	) name11438 (
		_w11401_,
		_w11469_,
		_w11470_,
		_w11472_
	);
	LUT3 #(
		.INIT('h06)
	) name11439 (
		_w11268_,
		_w11270_,
		_w11397_,
		_w11473_
	);
	LUT3 #(
		.INIT('h69)
	) name11440 (
		_w11268_,
		_w11270_,
		_w11397_,
		_w11474_
	);
	LUT4 #(
		.INIT('h629d)
	) name11441 (
		_w8616_,
		_w11268_,
		_w11269_,
		_w11272_,
		_w11475_
	);
	LUT4 #(
		.INIT('hba00)
	) name11442 (
		_w11398_,
		_w11472_,
		_w11474_,
		_w11475_,
		_w11476_
	);
	LUT4 #(
		.INIT('h5659)
	) name11443 (
		_w8466_,
		_w8541_,
		_w11273_,
		_w11393_,
		_w11477_
	);
	LUT4 #(
		.INIT('h0155)
	) name11444 (
		_w11395_,
		_w11396_,
		_w11476_,
		_w11477_,
		_w11478_
	);
	LUT3 #(
		.INIT('h06)
	) name11445 (
		_w11274_,
		_w11276_,
		_w11391_,
		_w11479_
	);
	LUT3 #(
		.INIT('h69)
	) name11446 (
		_w11274_,
		_w11276_,
		_w11391_,
		_w11480_
	);
	LUT4 #(
		.INIT('h629d)
	) name11447 (
		_w8150_,
		_w11274_,
		_w11275_,
		_w11278_,
		_w11481_
	);
	LUT4 #(
		.INIT('hba00)
	) name11448 (
		_w11392_,
		_w11478_,
		_w11480_,
		_w11481_,
		_w11482_
	);
	LUT4 #(
		.INIT('h5659)
	) name11449 (
		_w7935_,
		_w8077_,
		_w11279_,
		_w11387_,
		_w11483_
	);
	LUT4 #(
		.INIT('h0155)
	) name11450 (
		_w11389_,
		_w11390_,
		_w11482_,
		_w11483_,
		_w11484_
	);
	LUT3 #(
		.INIT('h06)
	) name11451 (
		_w11280_,
		_w11282_,
		_w11385_,
		_w11485_
	);
	LUT3 #(
		.INIT('h69)
	) name11452 (
		_w11280_,
		_w11282_,
		_w11385_,
		_w11486_
	);
	LUT4 #(
		.INIT('h629d)
	) name11453 (
		_w7816_,
		_w11280_,
		_w11281_,
		_w11284_,
		_w11487_
	);
	LUT4 #(
		.INIT('hba00)
	) name11454 (
		_w11386_,
		_w11484_,
		_w11486_,
		_w11487_,
		_w11488_
	);
	LUT4 #(
		.INIT('h5659)
	) name11455 (
		_w7695_,
		_w7750_,
		_w11285_,
		_w11381_,
		_w11489_
	);
	LUT4 #(
		.INIT('h0155)
	) name11456 (
		_w11383_,
		_w11384_,
		_w11488_,
		_w11489_,
		_w11490_
	);
	LUT3 #(
		.INIT('h06)
	) name11457 (
		_w11286_,
		_w11335_,
		_w11379_,
		_w11491_
	);
	LUT3 #(
		.INIT('h69)
	) name11458 (
		_w11286_,
		_w11335_,
		_w11379_,
		_w11492_
	);
	LUT4 #(
		.INIT('h8679)
	) name11459 (
		_w11333_,
		_w11286_,
		_w11335_,
		_w11374_,
		_w11493_
	);
	LUT4 #(
		.INIT('hba00)
	) name11460 (
		_w11380_,
		_w11490_,
		_w11492_,
		_w11493_,
		_w11494_
	);
	LUT4 #(
		.INIT('h028a)
	) name11461 (
		_w3214_,
		_w7136_,
		_w7166_,
		_w7167_,
		_w11495_
	);
	LUT2 #(
		.INIT('h1)
	) name11462 (
		_w11495_,
		_w11341_,
		_w11496_
	);
	LUT4 #(
		.INIT('h5700)
	) name11463 (
		_w37_,
		_w7418_,
		_w7419_,
		_w11496_,
		_w11497_
	);
	LUT2 #(
		.INIT('h6)
	) name11464 (
		\a[23] ,
		_w11497_,
		_w11498_
	);
	LUT3 #(
		.INIT('hd4)
	) name11465 (
		_w11369_,
		_w11370_,
		_w11351_,
		_w11499_
	);
	LUT4 #(
		.INIT('h0445)
	) name11466 (
		_w11498_,
		_w11369_,
		_w11370_,
		_w11351_,
		_w11500_
	);
	LUT4 #(
		.INIT('ha220)
	) name11467 (
		_w11498_,
		_w11369_,
		_w11370_,
		_w11351_,
		_w11501_
	);
	LUT4 #(
		.INIT('h599a)
	) name11468 (
		_w11498_,
		_w11369_,
		_w11370_,
		_w11351_,
		_w11502_
	);
	LUT4 #(
		.INIT('h6f06)
	) name11469 (
		_w11355_,
		_w11361_,
		_w11362_,
		_w11368_,
		_w11503_
	);
	LUT3 #(
		.INIT('h82)
	) name11470 (
		_w2550_,
		_w7129_,
		_w7131_,
		_w11504_
	);
	LUT3 #(
		.INIT('h84)
	) name11471 (
		_w2546_,
		_w2854_,
		_w6981_,
		_w11505_
	);
	LUT2 #(
		.INIT('h8)
	) name11472 (
		_w2549_,
		_w7002_,
		_w11506_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11473 (
		_w2617_,
		_w2622_,
		_w6978_,
		_w6980_,
		_w11507_
	);
	LUT2 #(
		.INIT('h1)
	) name11474 (
		_w11506_,
		_w11507_,
		_w11508_
	);
	LUT2 #(
		.INIT('h4)
	) name11475 (
		_w11505_,
		_w11508_,
		_w11509_
	);
	LUT3 #(
		.INIT('h9a)
	) name11476 (
		\a[29] ,
		_w11504_,
		_w11509_,
		_w11510_
	);
	LUT3 #(
		.INIT('h80)
	) name11477 (
		_w2015_,
		_w2573_,
		_w2696_,
		_w11511_
	);
	LUT4 #(
		.INIT('h135f)
	) name11478 (
		_w47_,
		_w93_,
		_w236_,
		_w166_,
		_w11512_
	);
	LUT4 #(
		.INIT('h8000)
	) name11479 (
		_w738_,
		_w957_,
		_w1248_,
		_w11512_,
		_w11513_
	);
	LUT4 #(
		.INIT('h1000)
	) name11480 (
		_w360_,
		_w443_,
		_w613_,
		_w2579_,
		_w11514_
	);
	LUT3 #(
		.INIT('h80)
	) name11481 (
		_w11511_,
		_w11513_,
		_w11514_,
		_w11515_
	);
	LUT3 #(
		.INIT('h80)
	) name11482 (
		_w739_,
		_w768_,
		_w1190_,
		_w11516_
	);
	LUT4 #(
		.INIT('h135f)
	) name11483 (
		_w56_,
		_w47_,
		_w166_,
		_w259_,
		_w11517_
	);
	LUT4 #(
		.INIT('h0777)
	) name11484 (
		_w122_,
		_w67_,
		_w41_,
		_w259_,
		_w11518_
	);
	LUT4 #(
		.INIT('h4000)
	) name11485 (
		_w476_,
		_w522_,
		_w11518_,
		_w11517_,
		_w11519_
	);
	LUT2 #(
		.INIT('h8)
	) name11486 (
		_w11516_,
		_w11519_,
		_w11520_
	);
	LUT3 #(
		.INIT('h80)
	) name11487 (
		_w646_,
		_w2690_,
		_w3802_,
		_w11521_
	);
	LUT3 #(
		.INIT('h80)
	) name11488 (
		_w11515_,
		_w11520_,
		_w11521_,
		_w11522_
	);
	LUT3 #(
		.INIT('h80)
	) name11489 (
		_w3106_,
		_w7195_,
		_w11522_,
		_w11523_
	);
	LUT2 #(
		.INIT('h9)
	) name11490 (
		_w7148_,
		_w11523_,
		_w11524_
	);
	LUT4 #(
		.INIT('h54ab)
	) name11491 (
		_w11353_,
		_w11354_,
		_w11361_,
		_w11524_,
		_w11525_
	);
	LUT3 #(
		.INIT('h82)
	) name11492 (
		_w377_,
		_w7123_,
		_w7125_,
		_w11526_
	);
	LUT3 #(
		.INIT('h82)
	) name11493 (
		_w2527_,
		_w2872_,
		_w6975_,
		_w11527_
	);
	LUT2 #(
		.INIT('h8)
	) name11494 (
		_w376_,
		_w7008_,
		_w11528_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11495 (
		_w2407_,
		_w2983_,
		_w6972_,
		_w6974_,
		_w11529_
	);
	LUT2 #(
		.INIT('h1)
	) name11496 (
		_w11528_,
		_w11529_,
		_w11530_
	);
	LUT2 #(
		.INIT('h4)
	) name11497 (
		_w11527_,
		_w11530_,
		_w11531_
	);
	LUT2 #(
		.INIT('h4)
	) name11498 (
		_w11526_,
		_w11531_,
		_w11532_
	);
	LUT3 #(
		.INIT('h96)
	) name11499 (
		_w11510_,
		_w11525_,
		_w11532_,
		_w11533_
	);
	LUT4 #(
		.INIT('h4114)
	) name11500 (
		_w11503_,
		_w11510_,
		_w11525_,
		_w11532_,
		_w11534_
	);
	LUT4 #(
		.INIT('h2882)
	) name11501 (
		_w11503_,
		_w11510_,
		_w11525_,
		_w11532_,
		_w11535_
	);
	LUT4 #(
		.INIT('h9669)
	) name11502 (
		_w11503_,
		_w11510_,
		_w11525_,
		_w11532_,
		_w11536_
	);
	LUT3 #(
		.INIT('h82)
	) name11503 (
		_w2875_,
		_w7135_,
		_w7172_,
		_w11537_
	);
	LUT3 #(
		.INIT('h28)
	) name11504 (
		_w2986_,
		_w7136_,
		_w7168_,
		_w11538_
	);
	LUT2 #(
		.INIT('h8)
	) name11505 (
		_w2874_,
		_w6996_,
		_w11539_
	);
	LUT4 #(
		.INIT('h04c8)
	) name11506 (
		_w2411_,
		_w2975_,
		_w6983_,
		_w6993_,
		_w11540_
	);
	LUT2 #(
		.INIT('h1)
	) name11507 (
		_w11539_,
		_w11540_,
		_w11541_
	);
	LUT2 #(
		.INIT('h4)
	) name11508 (
		_w11538_,
		_w11541_,
		_w11542_
	);
	LUT3 #(
		.INIT('h9a)
	) name11509 (
		\a[26] ,
		_w11537_,
		_w11542_,
		_w11543_
	);
	LUT2 #(
		.INIT('h9)
	) name11510 (
		_w11536_,
		_w11543_,
		_w11544_
	);
	LUT2 #(
		.INIT('h6)
	) name11511 (
		_w11502_,
		_w11544_,
		_w11545_
	);
	LUT3 #(
		.INIT('h17)
	) name11512 (
		_w11345_,
		_w11371_,
		_w11344_,
		_w11546_
	);
	LUT2 #(
		.INIT('h8)
	) name11513 (
		_w11545_,
		_w11546_,
		_w11547_
	);
	LUT2 #(
		.INIT('h1)
	) name11514 (
		_w11545_,
		_w11546_,
		_w11548_
	);
	LUT2 #(
		.INIT('h6)
	) name11515 (
		_w11545_,
		_w11546_,
		_w11549_
	);
	LUT3 #(
		.INIT('h56)
	) name11516 (
		_w11549_,
		_w11373_,
		_w11375_,
		_w11550_
	);
	LUT4 #(
		.INIT('h8218)
	) name11517 (
		_w11549_,
		_w11337_,
		_w11372_,
		_w11336_,
		_w11551_
	);
	LUT4 #(
		.INIT('h5659)
	) name11518 (
		_w11549_,
		_w11373_,
		_w11375_,
		_w11376_,
		_w11552_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11519 (
		_w35_,
		_w11378_,
		_w11494_,
		_w11552_,
		_w11553_
	);
	LUT4 #(
		.INIT('h2228)
	) name11520 (
		_w6324_,
		_w11549_,
		_w11373_,
		_w11375_,
		_w11554_
	);
	LUT3 #(
		.INIT('h82)
	) name11521 (
		_w5524_,
		_w11286_,
		_w11335_,
		_w11555_
	);
	LUT3 #(
		.INIT('h13)
	) name11522 (
		_w6031_,
		_w11555_,
		_w11377_,
		_w11556_
	);
	LUT2 #(
		.INIT('h4)
	) name11523 (
		_w11554_,
		_w11556_,
		_w11557_
	);
	LUT3 #(
		.INIT('h82)
	) name11524 (
		_w4459_,
		_w11478_,
		_w11480_,
		_w11558_
	);
	LUT3 #(
		.INIT('h82)
	) name11525 (
		_w4700_,
		_w11274_,
		_w11276_,
		_w11559_
	);
	LUT2 #(
		.INIT('h8)
	) name11526 (
		_w4458_,
		_w11394_,
		_w11560_
	);
	LUT4 #(
		.INIT('h2228)
	) name11527 (
		_w4684_,
		_w8466_,
		_w8541_,
		_w11273_,
		_w11561_
	);
	LUT2 #(
		.INIT('h1)
	) name11528 (
		_w11560_,
		_w11561_,
		_w11562_
	);
	LUT2 #(
		.INIT('h4)
	) name11529 (
		_w11559_,
		_w11562_,
		_w11563_
	);
	LUT3 #(
		.INIT('h82)
	) name11530 (
		_w4034_,
		_w11469_,
		_w11471_,
		_w11564_
	);
	LUT4 #(
		.INIT('h2228)
	) name11531 (
		_w4382_,
		_w8794_,
		_w8994_,
		_w11267_,
		_w11565_
	);
	LUT3 #(
		.INIT('h82)
	) name11532 (
		_w4033_,
		_w11262_,
		_w11264_,
		_w11566_
	);
	LUT3 #(
		.INIT('h07)
	) name11533 (
		_w4367_,
		_w11400_,
		_w11566_,
		_w11567_
	);
	LUT2 #(
		.INIT('h4)
	) name11534 (
		_w11565_,
		_w11567_,
		_w11568_
	);
	LUT4 #(
		.INIT('h54ab)
	) name11535 (
		_w11425_,
		_w11439_,
		_w11440_,
		_w11442_,
		_w11569_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11536 (
		_w3214_,
		_w10968_,
		_w11238_,
		_w11240_,
		_w11570_
	);
	LUT4 #(
		.INIT('h007d)
	) name11537 (
		_w3249_,
		_w11241_,
		_w11243_,
		_w11570_,
		_w11571_
	);
	LUT3 #(
		.INIT('h70)
	) name11538 (
		_w3262_,
		_w11421_,
		_w11571_,
		_w11572_
	);
	LUT4 #(
		.INIT('h95aa)
	) name11539 (
		\a[23] ,
		_w37_,
		_w11569_,
		_w11572_,
		_w11573_
	);
	LUT3 #(
		.INIT('h28)
	) name11540 (
		_w2875_,
		_w11431_,
		_w11435_,
		_w11574_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11541 (
		_w2874_,
		_w10991_,
		_w11230_,
		_w11232_,
		_w11575_
	);
	LUT4 #(
		.INIT('h007d)
	) name11542 (
		_w2975_,
		_w11233_,
		_w11235_,
		_w11575_,
		_w11576_
	);
	LUT3 #(
		.INIT('h70)
	) name11543 (
		_w2986_,
		_w11427_,
		_w11576_,
		_w11577_
	);
	LUT3 #(
		.INIT('h9a)
	) name11544 (
		\a[26] ,
		_w11574_,
		_w11577_,
		_w11578_
	);
	LUT2 #(
		.INIT('h4)
	) name11545 (
		_w2548_,
		_w11434_,
		_w11579_
	);
	LUT4 #(
		.INIT('h4029)
	) name11546 (
		_w10983_,
		_w10990_,
		_w11229_,
		_w11232_,
		_w11580_
	);
	LUT4 #(
		.INIT('he1d2)
	) name11547 (
		_w10991_,
		_w11230_,
		_w11232_,
		_w11433_,
		_w11581_
	);
	LUT2 #(
		.INIT('h8)
	) name11548 (
		_w2975_,
		_w11434_,
		_w11582_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11549 (
		_w2986_,
		_w10991_,
		_w11230_,
		_w11232_,
		_w11583_
	);
	LUT4 #(
		.INIT('h000d)
	) name11550 (
		_w2875_,
		_w11581_,
		_w11582_,
		_w11583_,
		_w11584_
	);
	LUT2 #(
		.INIT('h4)
	) name11551 (
		_w2873_,
		_w11434_,
		_w11585_
	);
	LUT3 #(
		.INIT('h8a)
	) name11552 (
		\a[26] ,
		_w2873_,
		_w11434_,
		_w11586_
	);
	LUT2 #(
		.INIT('h8)
	) name11553 (
		_w11584_,
		_w11586_,
		_w11587_
	);
	LUT4 #(
		.INIT('h2882)
	) name11554 (
		_w2875_,
		_w11233_,
		_w11235_,
		_w11580_,
		_w11588_
	);
	LUT3 #(
		.INIT('h82)
	) name11555 (
		_w2986_,
		_w11233_,
		_w11235_,
		_w11589_
	);
	LUT2 #(
		.INIT('h8)
	) name11556 (
		_w2874_,
		_w11434_,
		_w11590_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11557 (
		_w2975_,
		_w10991_,
		_w11230_,
		_w11232_,
		_w11591_
	);
	LUT2 #(
		.INIT('h1)
	) name11558 (
		_w11590_,
		_w11591_,
		_w11592_
	);
	LUT3 #(
		.INIT('h10)
	) name11559 (
		_w11589_,
		_w11588_,
		_w11592_,
		_w11593_
	);
	LUT3 #(
		.INIT('h80)
	) name11560 (
		_w11579_,
		_w11587_,
		_w11593_,
		_w11594_
	);
	LUT3 #(
		.INIT('h15)
	) name11561 (
		_w11579_,
		_w11587_,
		_w11593_,
		_w11595_
	);
	LUT3 #(
		.INIT('h6a)
	) name11562 (
		_w11579_,
		_w11587_,
		_w11593_,
		_w11596_
	);
	LUT2 #(
		.INIT('h9)
	) name11563 (
		_w11578_,
		_w11596_,
		_w11597_
	);
	LUT2 #(
		.INIT('h4)
	) name11564 (
		_w11573_,
		_w11597_,
		_w11598_
	);
	LUT3 #(
		.INIT('h82)
	) name11565 (
		_w37_,
		_w11439_,
		_w11441_,
		_w11599_
	);
	LUT3 #(
		.INIT('h82)
	) name11566 (
		_w3262_,
		_w11241_,
		_w11243_,
		_w11600_
	);
	LUT2 #(
		.INIT('h8)
	) name11567 (
		_w3214_,
		_w11427_,
		_w11601_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11568 (
		_w3249_,
		_w10968_,
		_w11238_,
		_w11240_,
		_w11602_
	);
	LUT2 #(
		.INIT('h1)
	) name11569 (
		_w11601_,
		_w11602_,
		_w11603_
	);
	LUT2 #(
		.INIT('h4)
	) name11570 (
		_w11600_,
		_w11603_,
		_w11604_
	);
	LUT3 #(
		.INIT('h8a)
	) name11571 (
		\a[26] ,
		_w11585_,
		_w11584_,
		_w11605_
	);
	LUT2 #(
		.INIT('h9)
	) name11572 (
		_w11593_,
		_w11605_,
		_w11606_
	);
	LUT4 #(
		.INIT('h6500)
	) name11573 (
		\a[23] ,
		_w11599_,
		_w11604_,
		_w11606_,
		_w11607_
	);
	LUT3 #(
		.INIT('h82)
	) name11574 (
		_w37_,
		_w11436_,
		_w11438_,
		_w11608_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11575 (
		_w3262_,
		_w10968_,
		_w11238_,
		_w11240_,
		_w11609_
	);
	LUT3 #(
		.INIT('h82)
	) name11576 (
		_w3214_,
		_w11233_,
		_w11235_,
		_w11610_
	);
	LUT3 #(
		.INIT('h07)
	) name11577 (
		_w3249_,
		_w11427_,
		_w11610_,
		_w11611_
	);
	LUT2 #(
		.INIT('h4)
	) name11578 (
		_w11609_,
		_w11611_,
		_w11612_
	);
	LUT3 #(
		.INIT('h20)
	) name11579 (
		\a[26] ,
		_w2873_,
		_w11434_,
		_w11613_
	);
	LUT2 #(
		.INIT('h9)
	) name11580 (
		_w11584_,
		_w11613_,
		_w11614_
	);
	LUT4 #(
		.INIT('h6500)
	) name11581 (
		\a[23] ,
		_w11608_,
		_w11612_,
		_w11614_,
		_w11615_
	);
	LUT2 #(
		.INIT('h8)
	) name11582 (
		_w3249_,
		_w11434_,
		_w11616_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11583 (
		_w3262_,
		_w10991_,
		_w11230_,
		_w11232_,
		_w11617_
	);
	LUT4 #(
		.INIT('h000d)
	) name11584 (
		_w37_,
		_w11581_,
		_w11616_,
		_w11617_,
		_w11618_
	);
	LUT2 #(
		.INIT('h4)
	) name11585 (
		_w36_,
		_w11434_,
		_w11619_
	);
	LUT3 #(
		.INIT('h8a)
	) name11586 (
		\a[23] ,
		_w36_,
		_w11434_,
		_w11620_
	);
	LUT2 #(
		.INIT('h8)
	) name11587 (
		_w11618_,
		_w11620_,
		_w11621_
	);
	LUT4 #(
		.INIT('h2882)
	) name11588 (
		_w37_,
		_w11233_,
		_w11235_,
		_w11580_,
		_w11622_
	);
	LUT3 #(
		.INIT('h82)
	) name11589 (
		_w3262_,
		_w11233_,
		_w11235_,
		_w11623_
	);
	LUT2 #(
		.INIT('h8)
	) name11590 (
		_w3214_,
		_w11434_,
		_w11624_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11591 (
		_w3249_,
		_w10991_,
		_w11230_,
		_w11232_,
		_w11625_
	);
	LUT2 #(
		.INIT('h1)
	) name11592 (
		_w11624_,
		_w11625_,
		_w11626_
	);
	LUT3 #(
		.INIT('h10)
	) name11593 (
		_w11623_,
		_w11622_,
		_w11626_,
		_w11627_
	);
	LUT3 #(
		.INIT('h80)
	) name11594 (
		_w11585_,
		_w11621_,
		_w11627_,
		_w11628_
	);
	LUT3 #(
		.INIT('h28)
	) name11595 (
		_w37_,
		_w11431_,
		_w11435_,
		_w11629_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11596 (
		_w3214_,
		_w10991_,
		_w11230_,
		_w11232_,
		_w11630_
	);
	LUT4 #(
		.INIT('h007d)
	) name11597 (
		_w3249_,
		_w11233_,
		_w11235_,
		_w11630_,
		_w11631_
	);
	LUT3 #(
		.INIT('h70)
	) name11598 (
		_w3262_,
		_w11427_,
		_w11631_,
		_w11632_
	);
	LUT3 #(
		.INIT('h9a)
	) name11599 (
		\a[23] ,
		_w11629_,
		_w11632_,
		_w11633_
	);
	LUT3 #(
		.INIT('h15)
	) name11600 (
		_w11585_,
		_w11621_,
		_w11627_,
		_w11634_
	);
	LUT3 #(
		.INIT('h6a)
	) name11601 (
		_w11585_,
		_w11621_,
		_w11627_,
		_w11635_
	);
	LUT3 #(
		.INIT('h54)
	) name11602 (
		_w11628_,
		_w11633_,
		_w11634_,
		_w11636_
	);
	LUT4 #(
		.INIT('h009a)
	) name11603 (
		\a[23] ,
		_w11608_,
		_w11612_,
		_w11614_,
		_w11637_
	);
	LUT4 #(
		.INIT('h9a65)
	) name11604 (
		\a[23] ,
		_w11608_,
		_w11612_,
		_w11614_,
		_w11638_
	);
	LUT3 #(
		.INIT('h54)
	) name11605 (
		_w11615_,
		_w11636_,
		_w11637_,
		_w11639_
	);
	LUT4 #(
		.INIT('h009a)
	) name11606 (
		\a[23] ,
		_w11599_,
		_w11604_,
		_w11606_,
		_w11640_
	);
	LUT4 #(
		.INIT('h9a65)
	) name11607 (
		\a[23] ,
		_w11599_,
		_w11604_,
		_w11606_,
		_w11641_
	);
	LUT3 #(
		.INIT('h54)
	) name11608 (
		_w11607_,
		_w11639_,
		_w11640_,
		_w11642_
	);
	LUT2 #(
		.INIT('h2)
	) name11609 (
		_w11573_,
		_w11597_,
		_w11643_
	);
	LUT2 #(
		.INIT('h9)
	) name11610 (
		_w11573_,
		_w11597_,
		_w11644_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11611 (
		_w37_,
		_w11423_,
		_w11443_,
		_w11444_,
		_w11645_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11612 (
		_w3262_,
		_w10945_,
		_w11246_,
		_w11248_,
		_w11646_
	);
	LUT3 #(
		.INIT('h82)
	) name11613 (
		_w3214_,
		_w11241_,
		_w11243_,
		_w11647_
	);
	LUT3 #(
		.INIT('h07)
	) name11614 (
		_w3249_,
		_w11421_,
		_w11647_,
		_w11648_
	);
	LUT2 #(
		.INIT('h4)
	) name11615 (
		_w11646_,
		_w11648_,
		_w11649_
	);
	LUT3 #(
		.INIT('h32)
	) name11616 (
		_w11578_,
		_w11594_,
		_w11595_,
		_w11650_
	);
	LUT3 #(
		.INIT('h82)
	) name11617 (
		_w2875_,
		_w11436_,
		_w11438_,
		_w11651_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11618 (
		_w2986_,
		_w10968_,
		_w11238_,
		_w11240_,
		_w11652_
	);
	LUT3 #(
		.INIT('h82)
	) name11619 (
		_w2874_,
		_w11233_,
		_w11235_,
		_w11653_
	);
	LUT3 #(
		.INIT('h07)
	) name11620 (
		_w2975_,
		_w11427_,
		_w11653_,
		_w11654_
	);
	LUT2 #(
		.INIT('h4)
	) name11621 (
		_w11652_,
		_w11654_,
		_w11655_
	);
	LUT3 #(
		.INIT('h20)
	) name11622 (
		\a[29] ,
		_w2548_,
		_w11434_,
		_w11656_
	);
	LUT2 #(
		.INIT('h8)
	) name11623 (
		_w2617_,
		_w11434_,
		_w11657_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11624 (
		_w2854_,
		_w10991_,
		_w11230_,
		_w11232_,
		_w11658_
	);
	LUT4 #(
		.INIT('h000d)
	) name11625 (
		_w2550_,
		_w11581_,
		_w11657_,
		_w11658_,
		_w11659_
	);
	LUT2 #(
		.INIT('h9)
	) name11626 (
		_w11656_,
		_w11659_,
		_w11660_
	);
	LUT4 #(
		.INIT('h6500)
	) name11627 (
		\a[26] ,
		_w11651_,
		_w11655_,
		_w11660_,
		_w11661_
	);
	LUT4 #(
		.INIT('h009a)
	) name11628 (
		\a[26] ,
		_w11651_,
		_w11655_,
		_w11660_,
		_w11662_
	);
	LUT4 #(
		.INIT('h9a65)
	) name11629 (
		\a[26] ,
		_w11651_,
		_w11655_,
		_w11660_,
		_w11663_
	);
	LUT2 #(
		.INIT('h9)
	) name11630 (
		_w11650_,
		_w11663_,
		_w11664_
	);
	LUT4 #(
		.INIT('h6500)
	) name11631 (
		\a[23] ,
		_w11645_,
		_w11649_,
		_w11664_,
		_w11665_
	);
	LUT4 #(
		.INIT('h9a65)
	) name11632 (
		\a[23] ,
		_w11645_,
		_w11649_,
		_w11664_,
		_w11666_
	);
	LUT4 #(
		.INIT('h4d00)
	) name11633 (
		_w11573_,
		_w11597_,
		_w11642_,
		_w11666_,
		_w11667_
	);
	LUT4 #(
		.INIT('h54ab)
	) name11634 (
		_w11598_,
		_w11642_,
		_w11643_,
		_w11666_,
		_w11668_
	);
	LUT3 #(
		.INIT('h82)
	) name11635 (
		_w3311_,
		_w11249_,
		_w11251_,
		_w11669_
	);
	LUT3 #(
		.INIT('h07)
	) name11636 (
		_w3645_,
		_w11415_,
		_w11669_,
		_w11670_
	);
	LUT4 #(
		.INIT('h7d00)
	) name11637 (
		_w3654_,
		_w10599_,
		_w11253_,
		_w11670_,
		_w11671_
	);
	LUT4 #(
		.INIT('h7d00)
	) name11638 (
		_w3312_,
		_w11450_,
		_w11452_,
		_w11671_,
		_w11672_
	);
	LUT3 #(
		.INIT('h84)
	) name11639 (
		\a[20] ,
		_w11668_,
		_w11672_,
		_w11673_
	);
	LUT2 #(
		.INIT('h9)
	) name11640 (
		_w11642_,
		_w11644_,
		_w11674_
	);
	LUT4 #(
		.INIT('h54ab)
	) name11641 (
		_w11419_,
		_w11445_,
		_w11446_,
		_w11448_,
		_w11675_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11642 (
		_w3311_,
		_w10945_,
		_w11246_,
		_w11248_,
		_w11676_
	);
	LUT4 #(
		.INIT('h007d)
	) name11643 (
		_w3645_,
		_w11249_,
		_w11251_,
		_w11676_,
		_w11677_
	);
	LUT3 #(
		.INIT('h70)
	) name11644 (
		_w3654_,
		_w11415_,
		_w11677_,
		_w11678_
	);
	LUT4 #(
		.INIT('h95aa)
	) name11645 (
		\a[20] ,
		_w3312_,
		_w11675_,
		_w11678_,
		_w11679_
	);
	LUT2 #(
		.INIT('h2)
	) name11646 (
		_w11674_,
		_w11679_,
		_w11680_
	);
	LUT2 #(
		.INIT('h9)
	) name11647 (
		_w11639_,
		_w11641_,
		_w11681_
	);
	LUT3 #(
		.INIT('h82)
	) name11648 (
		_w3312_,
		_w11445_,
		_w11447_,
		_w11682_
	);
	LUT3 #(
		.INIT('h82)
	) name11649 (
		_w3654_,
		_w11249_,
		_w11251_,
		_w11683_
	);
	LUT2 #(
		.INIT('h8)
	) name11650 (
		_w3311_,
		_w11421_,
		_w11684_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11651 (
		_w3645_,
		_w10945_,
		_w11246_,
		_w11248_,
		_w11685_
	);
	LUT2 #(
		.INIT('h1)
	) name11652 (
		_w11684_,
		_w11685_,
		_w11686_
	);
	LUT2 #(
		.INIT('h4)
	) name11653 (
		_w11683_,
		_w11686_,
		_w11687_
	);
	LUT4 #(
		.INIT('h4844)
	) name11654 (
		\a[20] ,
		_w11681_,
		_w11682_,
		_w11687_,
		_w11688_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11655 (
		_w3312_,
		_w11423_,
		_w11443_,
		_w11444_,
		_w11689_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11656 (
		_w3654_,
		_w10945_,
		_w11246_,
		_w11248_,
		_w11690_
	);
	LUT3 #(
		.INIT('h82)
	) name11657 (
		_w3311_,
		_w11241_,
		_w11243_,
		_w11691_
	);
	LUT3 #(
		.INIT('h07)
	) name11658 (
		_w3645_,
		_w11421_,
		_w11691_,
		_w11692_
	);
	LUT2 #(
		.INIT('h4)
	) name11659 (
		_w11690_,
		_w11692_,
		_w11693_
	);
	LUT2 #(
		.INIT('h9)
	) name11660 (
		_w11636_,
		_w11638_,
		_w11694_
	);
	LUT4 #(
		.INIT('h6500)
	) name11661 (
		\a[20] ,
		_w11689_,
		_w11693_,
		_w11694_,
		_w11695_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11662 (
		_w3311_,
		_w10968_,
		_w11238_,
		_w11240_,
		_w11696_
	);
	LUT4 #(
		.INIT('h007d)
	) name11663 (
		_w3645_,
		_w11241_,
		_w11243_,
		_w11696_,
		_w11697_
	);
	LUT3 #(
		.INIT('h70)
	) name11664 (
		_w3654_,
		_w11421_,
		_w11697_,
		_w11698_
	);
	LUT4 #(
		.INIT('h95aa)
	) name11665 (
		\a[20] ,
		_w3312_,
		_w11569_,
		_w11698_,
		_w11699_
	);
	LUT2 #(
		.INIT('h9)
	) name11666 (
		_w11633_,
		_w11635_,
		_w11700_
	);
	LUT2 #(
		.INIT('h4)
	) name11667 (
		_w11699_,
		_w11700_,
		_w11701_
	);
	LUT3 #(
		.INIT('h82)
	) name11668 (
		_w3312_,
		_w11439_,
		_w11441_,
		_w11702_
	);
	LUT3 #(
		.INIT('h82)
	) name11669 (
		_w3654_,
		_w11241_,
		_w11243_,
		_w11703_
	);
	LUT2 #(
		.INIT('h8)
	) name11670 (
		_w3311_,
		_w11427_,
		_w11704_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11671 (
		_w3645_,
		_w10968_,
		_w11238_,
		_w11240_,
		_w11705_
	);
	LUT2 #(
		.INIT('h1)
	) name11672 (
		_w11704_,
		_w11705_,
		_w11706_
	);
	LUT2 #(
		.INIT('h4)
	) name11673 (
		_w11703_,
		_w11706_,
		_w11707_
	);
	LUT3 #(
		.INIT('h8a)
	) name11674 (
		\a[23] ,
		_w11619_,
		_w11618_,
		_w11708_
	);
	LUT2 #(
		.INIT('h9)
	) name11675 (
		_w11627_,
		_w11708_,
		_w11709_
	);
	LUT4 #(
		.INIT('h6500)
	) name11676 (
		\a[20] ,
		_w11702_,
		_w11707_,
		_w11709_,
		_w11710_
	);
	LUT3 #(
		.INIT('h82)
	) name11677 (
		_w3312_,
		_w11436_,
		_w11438_,
		_w11711_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11678 (
		_w3654_,
		_w10968_,
		_w11238_,
		_w11240_,
		_w11712_
	);
	LUT3 #(
		.INIT('h82)
	) name11679 (
		_w3311_,
		_w11233_,
		_w11235_,
		_w11713_
	);
	LUT3 #(
		.INIT('h07)
	) name11680 (
		_w3645_,
		_w11427_,
		_w11713_,
		_w11714_
	);
	LUT2 #(
		.INIT('h4)
	) name11681 (
		_w11712_,
		_w11714_,
		_w11715_
	);
	LUT3 #(
		.INIT('h20)
	) name11682 (
		\a[23] ,
		_w36_,
		_w11434_,
		_w11716_
	);
	LUT2 #(
		.INIT('h9)
	) name11683 (
		_w11618_,
		_w11716_,
		_w11717_
	);
	LUT4 #(
		.INIT('h6500)
	) name11684 (
		\a[20] ,
		_w11711_,
		_w11715_,
		_w11717_,
		_w11718_
	);
	LUT2 #(
		.INIT('h8)
	) name11685 (
		_w3645_,
		_w11434_,
		_w11719_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11686 (
		_w3654_,
		_w10991_,
		_w11230_,
		_w11232_,
		_w11720_
	);
	LUT4 #(
		.INIT('h000d)
	) name11687 (
		_w3312_,
		_w11581_,
		_w11719_,
		_w11720_,
		_w11721_
	);
	LUT2 #(
		.INIT('h4)
	) name11688 (
		_w3310_,
		_w11434_,
		_w11722_
	);
	LUT3 #(
		.INIT('h8a)
	) name11689 (
		\a[20] ,
		_w3310_,
		_w11434_,
		_w11723_
	);
	LUT2 #(
		.INIT('h8)
	) name11690 (
		_w11721_,
		_w11723_,
		_w11724_
	);
	LUT4 #(
		.INIT('h2882)
	) name11691 (
		_w3312_,
		_w11233_,
		_w11235_,
		_w11580_,
		_w11725_
	);
	LUT3 #(
		.INIT('h82)
	) name11692 (
		_w3654_,
		_w11233_,
		_w11235_,
		_w11726_
	);
	LUT2 #(
		.INIT('h8)
	) name11693 (
		_w3311_,
		_w11434_,
		_w11727_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11694 (
		_w3645_,
		_w10991_,
		_w11230_,
		_w11232_,
		_w11728_
	);
	LUT2 #(
		.INIT('h1)
	) name11695 (
		_w11727_,
		_w11728_,
		_w11729_
	);
	LUT3 #(
		.INIT('h10)
	) name11696 (
		_w11726_,
		_w11725_,
		_w11729_,
		_w11730_
	);
	LUT3 #(
		.INIT('h80)
	) name11697 (
		_w11619_,
		_w11724_,
		_w11730_,
		_w11731_
	);
	LUT3 #(
		.INIT('h28)
	) name11698 (
		_w3312_,
		_w11431_,
		_w11435_,
		_w11732_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11699 (
		_w3311_,
		_w10991_,
		_w11230_,
		_w11232_,
		_w11733_
	);
	LUT4 #(
		.INIT('h007d)
	) name11700 (
		_w3645_,
		_w11233_,
		_w11235_,
		_w11733_,
		_w11734_
	);
	LUT3 #(
		.INIT('h70)
	) name11701 (
		_w3654_,
		_w11427_,
		_w11734_,
		_w11735_
	);
	LUT3 #(
		.INIT('h9a)
	) name11702 (
		\a[20] ,
		_w11732_,
		_w11735_,
		_w11736_
	);
	LUT3 #(
		.INIT('h15)
	) name11703 (
		_w11619_,
		_w11724_,
		_w11730_,
		_w11737_
	);
	LUT3 #(
		.INIT('h6a)
	) name11704 (
		_w11619_,
		_w11724_,
		_w11730_,
		_w11738_
	);
	LUT3 #(
		.INIT('h54)
	) name11705 (
		_w11731_,
		_w11736_,
		_w11737_,
		_w11739_
	);
	LUT4 #(
		.INIT('h009a)
	) name11706 (
		\a[20] ,
		_w11711_,
		_w11715_,
		_w11717_,
		_w11740_
	);
	LUT4 #(
		.INIT('h9a65)
	) name11707 (
		\a[20] ,
		_w11711_,
		_w11715_,
		_w11717_,
		_w11741_
	);
	LUT3 #(
		.INIT('h54)
	) name11708 (
		_w11718_,
		_w11739_,
		_w11740_,
		_w11742_
	);
	LUT4 #(
		.INIT('h009a)
	) name11709 (
		\a[20] ,
		_w11702_,
		_w11707_,
		_w11709_,
		_w11743_
	);
	LUT4 #(
		.INIT('h9a65)
	) name11710 (
		\a[20] ,
		_w11702_,
		_w11707_,
		_w11709_,
		_w11744_
	);
	LUT3 #(
		.INIT('h54)
	) name11711 (
		_w11710_,
		_w11742_,
		_w11743_,
		_w11745_
	);
	LUT2 #(
		.INIT('h2)
	) name11712 (
		_w11699_,
		_w11700_,
		_w11746_
	);
	LUT2 #(
		.INIT('h9)
	) name11713 (
		_w11699_,
		_w11700_,
		_w11747_
	);
	LUT4 #(
		.INIT('h9a65)
	) name11714 (
		\a[20] ,
		_w11689_,
		_w11693_,
		_w11694_,
		_w11748_
	);
	LUT4 #(
		.INIT('h4d00)
	) name11715 (
		_w11699_,
		_w11700_,
		_w11745_,
		_w11748_,
		_w11749_
	);
	LUT4 #(
		.INIT('h9699)
	) name11716 (
		\a[20] ,
		_w11681_,
		_w11682_,
		_w11687_,
		_w11750_
	);
	LUT4 #(
		.INIT('h0155)
	) name11717 (
		_w11688_,
		_w11695_,
		_w11749_,
		_w11750_,
		_w11751_
	);
	LUT2 #(
		.INIT('h4)
	) name11718 (
		_w11674_,
		_w11679_,
		_w11752_
	);
	LUT2 #(
		.INIT('h9)
	) name11719 (
		_w11674_,
		_w11679_,
		_w11753_
	);
	LUT3 #(
		.INIT('h54)
	) name11720 (
		_w11680_,
		_w11751_,
		_w11752_,
		_w11754_
	);
	LUT3 #(
		.INIT('h12)
	) name11721 (
		\a[20] ,
		_w11668_,
		_w11672_,
		_w11755_
	);
	LUT3 #(
		.INIT('h69)
	) name11722 (
		\a[20] ,
		_w11668_,
		_w11672_,
		_w11756_
	);
	LUT3 #(
		.INIT('h54)
	) name11723 (
		_w11673_,
		_w11754_,
		_w11755_,
		_w11757_
	);
	LUT2 #(
		.INIT('h8)
	) name11724 (
		_w3311_,
		_w11415_,
		_w11758_
	);
	LUT4 #(
		.INIT('h007d)
	) name11725 (
		_w3645_,
		_w10599_,
		_w11253_,
		_w11758_,
		_w11759_
	);
	LUT4 #(
		.INIT('h7d00)
	) name11726 (
		_w3654_,
		_w10580_,
		_w11254_,
		_w11759_,
		_w11760_
	);
	LUT4 #(
		.INIT('h7d00)
	) name11727 (
		_w3312_,
		_w11453_,
		_w11455_,
		_w11760_,
		_w11761_
	);
	LUT3 #(
		.INIT('h32)
	) name11728 (
		_w11650_,
		_w11661_,
		_w11662_,
		_w11762_
	);
	LUT3 #(
		.INIT('h82)
	) name11729 (
		_w2875_,
		_w11439_,
		_w11441_,
		_w11763_
	);
	LUT3 #(
		.INIT('h82)
	) name11730 (
		_w2986_,
		_w11241_,
		_w11243_,
		_w11764_
	);
	LUT2 #(
		.INIT('h8)
	) name11731 (
		_w2874_,
		_w11427_,
		_w11765_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11732 (
		_w2975_,
		_w10968_,
		_w11238_,
		_w11240_,
		_w11766_
	);
	LUT2 #(
		.INIT('h1)
	) name11733 (
		_w11765_,
		_w11766_,
		_w11767_
	);
	LUT2 #(
		.INIT('h4)
	) name11734 (
		_w11764_,
		_w11767_,
		_w11768_
	);
	LUT3 #(
		.INIT('h8a)
	) name11735 (
		\a[29] ,
		_w2548_,
		_w11434_,
		_w11769_
	);
	LUT2 #(
		.INIT('h8)
	) name11736 (
		_w11659_,
		_w11769_,
		_w11770_
	);
	LUT3 #(
		.INIT('h8a)
	) name11737 (
		\a[29] ,
		_w11579_,
		_w11659_,
		_w11771_
	);
	LUT4 #(
		.INIT('h2882)
	) name11738 (
		_w2550_,
		_w11233_,
		_w11235_,
		_w11580_,
		_w11772_
	);
	LUT3 #(
		.INIT('h82)
	) name11739 (
		_w2854_,
		_w11233_,
		_w11235_,
		_w11773_
	);
	LUT2 #(
		.INIT('h8)
	) name11740 (
		_w2549_,
		_w11434_,
		_w11774_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11741 (
		_w2617_,
		_w10991_,
		_w11230_,
		_w11232_,
		_w11775_
	);
	LUT2 #(
		.INIT('h1)
	) name11742 (
		_w11774_,
		_w11775_,
		_w11776_
	);
	LUT3 #(
		.INIT('h10)
	) name11743 (
		_w11773_,
		_w11772_,
		_w11776_,
		_w11777_
	);
	LUT2 #(
		.INIT('h9)
	) name11744 (
		_w11771_,
		_w11777_,
		_w11778_
	);
	LUT4 #(
		.INIT('h6500)
	) name11745 (
		\a[26] ,
		_w11763_,
		_w11768_,
		_w11778_,
		_w11779_
	);
	LUT4 #(
		.INIT('h009a)
	) name11746 (
		\a[26] ,
		_w11763_,
		_w11768_,
		_w11778_,
		_w11780_
	);
	LUT4 #(
		.INIT('h9a65)
	) name11747 (
		\a[26] ,
		_w11763_,
		_w11768_,
		_w11778_,
		_w11781_
	);
	LUT2 #(
		.INIT('h9)
	) name11748 (
		_w11762_,
		_w11781_,
		_w11782_
	);
	LUT3 #(
		.INIT('h82)
	) name11749 (
		_w37_,
		_w11445_,
		_w11447_,
		_w11783_
	);
	LUT3 #(
		.INIT('h82)
	) name11750 (
		_w3262_,
		_w11249_,
		_w11251_,
		_w11784_
	);
	LUT2 #(
		.INIT('h8)
	) name11751 (
		_w3214_,
		_w11421_,
		_w11785_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11752 (
		_w3249_,
		_w10945_,
		_w11246_,
		_w11248_,
		_w11786_
	);
	LUT2 #(
		.INIT('h1)
	) name11753 (
		_w11785_,
		_w11786_,
		_w11787_
	);
	LUT2 #(
		.INIT('h4)
	) name11754 (
		_w11784_,
		_w11787_,
		_w11788_
	);
	LUT4 #(
		.INIT('h4844)
	) name11755 (
		\a[23] ,
		_w11782_,
		_w11783_,
		_w11788_,
		_w11789_
	);
	LUT4 #(
		.INIT('h9699)
	) name11756 (
		\a[23] ,
		_w11782_,
		_w11783_,
		_w11788_,
		_w11790_
	);
	LUT3 #(
		.INIT('h1e)
	) name11757 (
		_w11665_,
		_w11667_,
		_w11790_,
		_w11791_
	);
	LUT3 #(
		.INIT('h90)
	) name11758 (
		\a[20] ,
		_w11761_,
		_w11791_,
		_w11792_
	);
	LUT3 #(
		.INIT('h06)
	) name11759 (
		\a[20] ,
		_w11761_,
		_w11791_,
		_w11793_
	);
	LUT3 #(
		.INIT('h69)
	) name11760 (
		\a[20] ,
		_w11761_,
		_w11791_,
		_w11794_
	);
	LUT2 #(
		.INIT('h9)
	) name11761 (
		_w11757_,
		_w11794_,
		_w11795_
	);
	LUT4 #(
		.INIT('h54ab)
	) name11762 (
		_w11410_,
		_w11459_,
		_w11460_,
		_w11462_,
		_w11796_
	);
	LUT3 #(
		.INIT('h82)
	) name11763 (
		_w3709_,
		_w10268_,
		_w11255_,
		_w11797_
	);
	LUT4 #(
		.INIT('h007d)
	) name11764 (
		_w3877_,
		_w11256_,
		_w11258_,
		_w11797_,
		_w11798_
	);
	LUT3 #(
		.INIT('h70)
	) name11765 (
		_w3886_,
		_w11406_,
		_w11798_,
		_w11799_
	);
	LUT4 #(
		.INIT('h95aa)
	) name11766 (
		\a[17] ,
		_w3710_,
		_w11796_,
		_w11799_,
		_w11800_
	);
	LUT2 #(
		.INIT('h2)
	) name11767 (
		_w11795_,
		_w11800_,
		_w11801_
	);
	LUT3 #(
		.INIT('h82)
	) name11768 (
		_w3709_,
		_w10580_,
		_w11254_,
		_w11802_
	);
	LUT4 #(
		.INIT('h007d)
	) name11769 (
		_w3877_,
		_w10268_,
		_w11255_,
		_w11802_,
		_w11803_
	);
	LUT4 #(
		.INIT('h7d00)
	) name11770 (
		_w3886_,
		_w11256_,
		_w11258_,
		_w11803_,
		_w11804_
	);
	LUT4 #(
		.INIT('h7d00)
	) name11771 (
		_w3710_,
		_w11459_,
		_w11461_,
		_w11804_,
		_w11805_
	);
	LUT2 #(
		.INIT('h9)
	) name11772 (
		_w11754_,
		_w11756_,
		_w11806_
	);
	LUT3 #(
		.INIT('h90)
	) name11773 (
		\a[17] ,
		_w11805_,
		_w11806_,
		_w11807_
	);
	LUT3 #(
		.INIT('h82)
	) name11774 (
		_w3709_,
		_w10599_,
		_w11253_,
		_w11808_
	);
	LUT4 #(
		.INIT('h007d)
	) name11775 (
		_w3877_,
		_w10580_,
		_w11254_,
		_w11808_,
		_w11809_
	);
	LUT4 #(
		.INIT('h7d00)
	) name11776 (
		_w3886_,
		_w10268_,
		_w11255_,
		_w11809_,
		_w11810_
	);
	LUT4 #(
		.INIT('h7d00)
	) name11777 (
		_w3710_,
		_w11456_,
		_w11458_,
		_w11810_,
		_w11811_
	);
	LUT2 #(
		.INIT('h9)
	) name11778 (
		_w11751_,
		_w11753_,
		_w11812_
	);
	LUT3 #(
		.INIT('h90)
	) name11779 (
		\a[17] ,
		_w11811_,
		_w11812_,
		_w11813_
	);
	LUT2 #(
		.INIT('h8)
	) name11780 (
		_w3709_,
		_w11415_,
		_w11814_
	);
	LUT4 #(
		.INIT('h007d)
	) name11781 (
		_w3877_,
		_w10599_,
		_w11253_,
		_w11814_,
		_w11815_
	);
	LUT4 #(
		.INIT('h7d00)
	) name11782 (
		_w3886_,
		_w10580_,
		_w11254_,
		_w11815_,
		_w11816_
	);
	LUT4 #(
		.INIT('h7d00)
	) name11783 (
		_w3710_,
		_w11453_,
		_w11455_,
		_w11816_,
		_w11817_
	);
	LUT3 #(
		.INIT('h1e)
	) name11784 (
		_w11695_,
		_w11749_,
		_w11750_,
		_w11818_
	);
	LUT3 #(
		.INIT('h90)
	) name11785 (
		\a[17] ,
		_w11817_,
		_w11818_,
		_w11819_
	);
	LUT4 #(
		.INIT('h54ab)
	) name11786 (
		_w11701_,
		_w11745_,
		_w11746_,
		_w11748_,
		_w11820_
	);
	LUT3 #(
		.INIT('h82)
	) name11787 (
		_w3709_,
		_w11249_,
		_w11251_,
		_w11821_
	);
	LUT3 #(
		.INIT('h07)
	) name11788 (
		_w3877_,
		_w11415_,
		_w11821_,
		_w11822_
	);
	LUT4 #(
		.INIT('h7d00)
	) name11789 (
		_w3886_,
		_w10599_,
		_w11253_,
		_w11822_,
		_w11823_
	);
	LUT4 #(
		.INIT('h7d00)
	) name11790 (
		_w3710_,
		_w11450_,
		_w11452_,
		_w11823_,
		_w11824_
	);
	LUT3 #(
		.INIT('h84)
	) name11791 (
		\a[17] ,
		_w11820_,
		_w11824_,
		_w11825_
	);
	LUT2 #(
		.INIT('h9)
	) name11792 (
		_w11745_,
		_w11747_,
		_w11826_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11793 (
		_w3709_,
		_w10945_,
		_w11246_,
		_w11248_,
		_w11827_
	);
	LUT4 #(
		.INIT('h007d)
	) name11794 (
		_w3877_,
		_w11249_,
		_w11251_,
		_w11827_,
		_w11828_
	);
	LUT3 #(
		.INIT('h70)
	) name11795 (
		_w3886_,
		_w11415_,
		_w11828_,
		_w11829_
	);
	LUT4 #(
		.INIT('h95aa)
	) name11796 (
		\a[17] ,
		_w3710_,
		_w11675_,
		_w11829_,
		_w11830_
	);
	LUT2 #(
		.INIT('h2)
	) name11797 (
		_w11826_,
		_w11830_,
		_w11831_
	);
	LUT2 #(
		.INIT('h9)
	) name11798 (
		_w11742_,
		_w11744_,
		_w11832_
	);
	LUT3 #(
		.INIT('h82)
	) name11799 (
		_w3710_,
		_w11445_,
		_w11447_,
		_w11833_
	);
	LUT3 #(
		.INIT('h82)
	) name11800 (
		_w3886_,
		_w11249_,
		_w11251_,
		_w11834_
	);
	LUT2 #(
		.INIT('h8)
	) name11801 (
		_w3709_,
		_w11421_,
		_w11835_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11802 (
		_w3877_,
		_w10945_,
		_w11246_,
		_w11248_,
		_w11836_
	);
	LUT2 #(
		.INIT('h1)
	) name11803 (
		_w11835_,
		_w11836_,
		_w11837_
	);
	LUT2 #(
		.INIT('h4)
	) name11804 (
		_w11834_,
		_w11837_,
		_w11838_
	);
	LUT4 #(
		.INIT('h4844)
	) name11805 (
		\a[17] ,
		_w11832_,
		_w11833_,
		_w11838_,
		_w11839_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11806 (
		_w3710_,
		_w11423_,
		_w11443_,
		_w11444_,
		_w11840_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11807 (
		_w3886_,
		_w10945_,
		_w11246_,
		_w11248_,
		_w11841_
	);
	LUT3 #(
		.INIT('h82)
	) name11808 (
		_w3709_,
		_w11241_,
		_w11243_,
		_w11842_
	);
	LUT3 #(
		.INIT('h07)
	) name11809 (
		_w3877_,
		_w11421_,
		_w11842_,
		_w11843_
	);
	LUT2 #(
		.INIT('h4)
	) name11810 (
		_w11841_,
		_w11843_,
		_w11844_
	);
	LUT2 #(
		.INIT('h9)
	) name11811 (
		_w11739_,
		_w11741_,
		_w11845_
	);
	LUT4 #(
		.INIT('h6500)
	) name11812 (
		\a[17] ,
		_w11840_,
		_w11844_,
		_w11845_,
		_w11846_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11813 (
		_w3709_,
		_w10968_,
		_w11238_,
		_w11240_,
		_w11847_
	);
	LUT4 #(
		.INIT('h007d)
	) name11814 (
		_w3877_,
		_w11241_,
		_w11243_,
		_w11847_,
		_w11848_
	);
	LUT3 #(
		.INIT('h70)
	) name11815 (
		_w3886_,
		_w11421_,
		_w11848_,
		_w11849_
	);
	LUT4 #(
		.INIT('h95aa)
	) name11816 (
		\a[17] ,
		_w3710_,
		_w11569_,
		_w11849_,
		_w11850_
	);
	LUT2 #(
		.INIT('h9)
	) name11817 (
		_w11736_,
		_w11738_,
		_w11851_
	);
	LUT2 #(
		.INIT('h4)
	) name11818 (
		_w11850_,
		_w11851_,
		_w11852_
	);
	LUT3 #(
		.INIT('h82)
	) name11819 (
		_w3710_,
		_w11439_,
		_w11441_,
		_w11853_
	);
	LUT3 #(
		.INIT('h82)
	) name11820 (
		_w3886_,
		_w11241_,
		_w11243_,
		_w11854_
	);
	LUT2 #(
		.INIT('h8)
	) name11821 (
		_w3709_,
		_w11427_,
		_w11855_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11822 (
		_w3877_,
		_w10968_,
		_w11238_,
		_w11240_,
		_w11856_
	);
	LUT2 #(
		.INIT('h1)
	) name11823 (
		_w11855_,
		_w11856_,
		_w11857_
	);
	LUT2 #(
		.INIT('h4)
	) name11824 (
		_w11854_,
		_w11857_,
		_w11858_
	);
	LUT3 #(
		.INIT('h8a)
	) name11825 (
		\a[20] ,
		_w11722_,
		_w11721_,
		_w11859_
	);
	LUT2 #(
		.INIT('h9)
	) name11826 (
		_w11730_,
		_w11859_,
		_w11860_
	);
	LUT4 #(
		.INIT('h6500)
	) name11827 (
		\a[17] ,
		_w11853_,
		_w11858_,
		_w11860_,
		_w11861_
	);
	LUT3 #(
		.INIT('h82)
	) name11828 (
		_w3710_,
		_w11436_,
		_w11438_,
		_w11862_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11829 (
		_w3886_,
		_w10968_,
		_w11238_,
		_w11240_,
		_w11863_
	);
	LUT3 #(
		.INIT('h82)
	) name11830 (
		_w3709_,
		_w11233_,
		_w11235_,
		_w11864_
	);
	LUT3 #(
		.INIT('h07)
	) name11831 (
		_w3877_,
		_w11427_,
		_w11864_,
		_w11865_
	);
	LUT2 #(
		.INIT('h4)
	) name11832 (
		_w11863_,
		_w11865_,
		_w11866_
	);
	LUT3 #(
		.INIT('h20)
	) name11833 (
		\a[20] ,
		_w3310_,
		_w11434_,
		_w11867_
	);
	LUT2 #(
		.INIT('h9)
	) name11834 (
		_w11721_,
		_w11867_,
		_w11868_
	);
	LUT4 #(
		.INIT('h6500)
	) name11835 (
		\a[17] ,
		_w11862_,
		_w11866_,
		_w11868_,
		_w11869_
	);
	LUT2 #(
		.INIT('h8)
	) name11836 (
		_w3877_,
		_w11434_,
		_w11870_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11837 (
		_w3886_,
		_w10991_,
		_w11230_,
		_w11232_,
		_w11871_
	);
	LUT4 #(
		.INIT('h000d)
	) name11838 (
		_w3710_,
		_w11581_,
		_w11870_,
		_w11871_,
		_w11872_
	);
	LUT2 #(
		.INIT('h4)
	) name11839 (
		_w3708_,
		_w11434_,
		_w11873_
	);
	LUT3 #(
		.INIT('h8a)
	) name11840 (
		\a[17] ,
		_w3708_,
		_w11434_,
		_w11874_
	);
	LUT2 #(
		.INIT('h8)
	) name11841 (
		_w11872_,
		_w11874_,
		_w11875_
	);
	LUT4 #(
		.INIT('h2882)
	) name11842 (
		_w3710_,
		_w11233_,
		_w11235_,
		_w11580_,
		_w11876_
	);
	LUT3 #(
		.INIT('h82)
	) name11843 (
		_w3886_,
		_w11233_,
		_w11235_,
		_w11877_
	);
	LUT2 #(
		.INIT('h8)
	) name11844 (
		_w3709_,
		_w11434_,
		_w11878_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11845 (
		_w3877_,
		_w10991_,
		_w11230_,
		_w11232_,
		_w11879_
	);
	LUT2 #(
		.INIT('h1)
	) name11846 (
		_w11878_,
		_w11879_,
		_w11880_
	);
	LUT3 #(
		.INIT('h10)
	) name11847 (
		_w11877_,
		_w11876_,
		_w11880_,
		_w11881_
	);
	LUT3 #(
		.INIT('h80)
	) name11848 (
		_w11722_,
		_w11875_,
		_w11881_,
		_w11882_
	);
	LUT3 #(
		.INIT('h28)
	) name11849 (
		_w3710_,
		_w11431_,
		_w11435_,
		_w11883_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11850 (
		_w3709_,
		_w10991_,
		_w11230_,
		_w11232_,
		_w11884_
	);
	LUT4 #(
		.INIT('h007d)
	) name11851 (
		_w3877_,
		_w11233_,
		_w11235_,
		_w11884_,
		_w11885_
	);
	LUT3 #(
		.INIT('h70)
	) name11852 (
		_w3886_,
		_w11427_,
		_w11885_,
		_w11886_
	);
	LUT3 #(
		.INIT('h9a)
	) name11853 (
		\a[17] ,
		_w11883_,
		_w11886_,
		_w11887_
	);
	LUT3 #(
		.INIT('h15)
	) name11854 (
		_w11722_,
		_w11875_,
		_w11881_,
		_w11888_
	);
	LUT3 #(
		.INIT('h6a)
	) name11855 (
		_w11722_,
		_w11875_,
		_w11881_,
		_w11889_
	);
	LUT3 #(
		.INIT('h54)
	) name11856 (
		_w11882_,
		_w11887_,
		_w11888_,
		_w11890_
	);
	LUT4 #(
		.INIT('h009a)
	) name11857 (
		\a[17] ,
		_w11862_,
		_w11866_,
		_w11868_,
		_w11891_
	);
	LUT4 #(
		.INIT('h9a65)
	) name11858 (
		\a[17] ,
		_w11862_,
		_w11866_,
		_w11868_,
		_w11892_
	);
	LUT3 #(
		.INIT('h54)
	) name11859 (
		_w11869_,
		_w11890_,
		_w11891_,
		_w11893_
	);
	LUT4 #(
		.INIT('h009a)
	) name11860 (
		\a[17] ,
		_w11853_,
		_w11858_,
		_w11860_,
		_w11894_
	);
	LUT4 #(
		.INIT('h9a65)
	) name11861 (
		\a[17] ,
		_w11853_,
		_w11858_,
		_w11860_,
		_w11895_
	);
	LUT3 #(
		.INIT('h54)
	) name11862 (
		_w11861_,
		_w11893_,
		_w11894_,
		_w11896_
	);
	LUT2 #(
		.INIT('h2)
	) name11863 (
		_w11850_,
		_w11851_,
		_w11897_
	);
	LUT2 #(
		.INIT('h9)
	) name11864 (
		_w11850_,
		_w11851_,
		_w11898_
	);
	LUT4 #(
		.INIT('h9a65)
	) name11865 (
		\a[17] ,
		_w11840_,
		_w11844_,
		_w11845_,
		_w11899_
	);
	LUT4 #(
		.INIT('h4d00)
	) name11866 (
		_w11850_,
		_w11851_,
		_w11896_,
		_w11899_,
		_w11900_
	);
	LUT4 #(
		.INIT('h9699)
	) name11867 (
		\a[17] ,
		_w11832_,
		_w11833_,
		_w11838_,
		_w11901_
	);
	LUT4 #(
		.INIT('h0155)
	) name11868 (
		_w11839_,
		_w11846_,
		_w11900_,
		_w11901_,
		_w11902_
	);
	LUT2 #(
		.INIT('h4)
	) name11869 (
		_w11826_,
		_w11830_,
		_w11903_
	);
	LUT2 #(
		.INIT('h9)
	) name11870 (
		_w11826_,
		_w11830_,
		_w11904_
	);
	LUT3 #(
		.INIT('h54)
	) name11871 (
		_w11831_,
		_w11902_,
		_w11903_,
		_w11905_
	);
	LUT3 #(
		.INIT('h12)
	) name11872 (
		\a[17] ,
		_w11820_,
		_w11824_,
		_w11906_
	);
	LUT3 #(
		.INIT('h69)
	) name11873 (
		\a[17] ,
		_w11820_,
		_w11824_,
		_w11907_
	);
	LUT3 #(
		.INIT('h54)
	) name11874 (
		_w11825_,
		_w11905_,
		_w11906_,
		_w11908_
	);
	LUT3 #(
		.INIT('h06)
	) name11875 (
		\a[17] ,
		_w11817_,
		_w11818_,
		_w11909_
	);
	LUT3 #(
		.INIT('h69)
	) name11876 (
		\a[17] ,
		_w11817_,
		_w11818_,
		_w11910_
	);
	LUT3 #(
		.INIT('h54)
	) name11877 (
		_w11819_,
		_w11908_,
		_w11909_,
		_w11911_
	);
	LUT3 #(
		.INIT('h06)
	) name11878 (
		\a[17] ,
		_w11811_,
		_w11812_,
		_w11912_
	);
	LUT3 #(
		.INIT('h69)
	) name11879 (
		\a[17] ,
		_w11811_,
		_w11812_,
		_w11913_
	);
	LUT3 #(
		.INIT('h54)
	) name11880 (
		_w11813_,
		_w11911_,
		_w11912_,
		_w11914_
	);
	LUT3 #(
		.INIT('h06)
	) name11881 (
		\a[17] ,
		_w11805_,
		_w11806_,
		_w11915_
	);
	LUT3 #(
		.INIT('h69)
	) name11882 (
		\a[17] ,
		_w11805_,
		_w11806_,
		_w11916_
	);
	LUT3 #(
		.INIT('h54)
	) name11883 (
		_w11807_,
		_w11914_,
		_w11915_,
		_w11917_
	);
	LUT2 #(
		.INIT('h4)
	) name11884 (
		_w11795_,
		_w11800_,
		_w11918_
	);
	LUT2 #(
		.INIT('h9)
	) name11885 (
		_w11795_,
		_w11800_,
		_w11919_
	);
	LUT3 #(
		.INIT('h32)
	) name11886 (
		_w11757_,
		_w11792_,
		_w11793_,
		_w11920_
	);
	LUT3 #(
		.INIT('h82)
	) name11887 (
		_w3311_,
		_w10599_,
		_w11253_,
		_w11921_
	);
	LUT4 #(
		.INIT('h007d)
	) name11888 (
		_w3645_,
		_w10580_,
		_w11254_,
		_w11921_,
		_w11922_
	);
	LUT4 #(
		.INIT('h7d00)
	) name11889 (
		_w3654_,
		_w10268_,
		_w11255_,
		_w11922_,
		_w11923_
	);
	LUT4 #(
		.INIT('h7d00)
	) name11890 (
		_w3312_,
		_w11456_,
		_w11458_,
		_w11923_,
		_w11924_
	);
	LUT4 #(
		.INIT('h010f)
	) name11891 (
		_w11665_,
		_w11667_,
		_w11789_,
		_w11790_,
		_w11925_
	);
	LUT3 #(
		.INIT('h32)
	) name11892 (
		_w11762_,
		_w11779_,
		_w11780_,
		_w11926_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11893 (
		_w2874_,
		_w10968_,
		_w11238_,
		_w11240_,
		_w11927_
	);
	LUT4 #(
		.INIT('h007d)
	) name11894 (
		_w2975_,
		_w11241_,
		_w11243_,
		_w11927_,
		_w11928_
	);
	LUT3 #(
		.INIT('h70)
	) name11895 (
		_w2986_,
		_w11421_,
		_w11928_,
		_w11929_
	);
	LUT4 #(
		.INIT('h95aa)
	) name11896 (
		\a[26] ,
		_w2875_,
		_w11569_,
		_w11929_,
		_w11930_
	);
	LUT3 #(
		.INIT('h28)
	) name11897 (
		_w2550_,
		_w11431_,
		_w11435_,
		_w11931_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11898 (
		_w2549_,
		_w10991_,
		_w11230_,
		_w11232_,
		_w11932_
	);
	LUT4 #(
		.INIT('h007d)
	) name11899 (
		_w2617_,
		_w11233_,
		_w11235_,
		_w11932_,
		_w11933_
	);
	LUT3 #(
		.INIT('h70)
	) name11900 (
		_w2854_,
		_w11427_,
		_w11933_,
		_w11934_
	);
	LUT3 #(
		.INIT('h9a)
	) name11901 (
		\a[29] ,
		_w11931_,
		_w11934_,
		_w11935_
	);
	LUT2 #(
		.INIT('h4)
	) name11902 (
		_w375_,
		_w11434_,
		_w11936_
	);
	LUT3 #(
		.INIT('h80)
	) name11903 (
		_w11770_,
		_w11777_,
		_w11936_,
		_w11937_
	);
	LUT3 #(
		.INIT('h07)
	) name11904 (
		_w11770_,
		_w11777_,
		_w11936_,
		_w11938_
	);
	LUT3 #(
		.INIT('h78)
	) name11905 (
		_w11770_,
		_w11777_,
		_w11936_,
		_w11939_
	);
	LUT2 #(
		.INIT('h9)
	) name11906 (
		_w11935_,
		_w11939_,
		_w11940_
	);
	LUT2 #(
		.INIT('h4)
	) name11907 (
		_w11930_,
		_w11940_,
		_w11941_
	);
	LUT2 #(
		.INIT('h2)
	) name11908 (
		_w11930_,
		_w11940_,
		_w11942_
	);
	LUT2 #(
		.INIT('h9)
	) name11909 (
		_w11930_,
		_w11940_,
		_w11943_
	);
	LUT2 #(
		.INIT('h9)
	) name11910 (
		_w11926_,
		_w11943_,
		_w11944_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11911 (
		_w3214_,
		_w10945_,
		_w11246_,
		_w11248_,
		_w11945_
	);
	LUT4 #(
		.INIT('h007d)
	) name11912 (
		_w3249_,
		_w11249_,
		_w11251_,
		_w11945_,
		_w11946_
	);
	LUT3 #(
		.INIT('h70)
	) name11913 (
		_w3262_,
		_w11415_,
		_w11946_,
		_w11947_
	);
	LUT4 #(
		.INIT('h95aa)
	) name11914 (
		\a[23] ,
		_w37_,
		_w11675_,
		_w11947_,
		_w11948_
	);
	LUT2 #(
		.INIT('h2)
	) name11915 (
		_w11944_,
		_w11948_,
		_w11949_
	);
	LUT2 #(
		.INIT('h4)
	) name11916 (
		_w11944_,
		_w11948_,
		_w11950_
	);
	LUT2 #(
		.INIT('h9)
	) name11917 (
		_w11944_,
		_w11948_,
		_w11951_
	);
	LUT2 #(
		.INIT('h9)
	) name11918 (
		_w11925_,
		_w11951_,
		_w11952_
	);
	LUT3 #(
		.INIT('h90)
	) name11919 (
		\a[20] ,
		_w11924_,
		_w11952_,
		_w11953_
	);
	LUT3 #(
		.INIT('h06)
	) name11920 (
		\a[20] ,
		_w11924_,
		_w11952_,
		_w11954_
	);
	LUT3 #(
		.INIT('h69)
	) name11921 (
		\a[20] ,
		_w11924_,
		_w11952_,
		_w11955_
	);
	LUT2 #(
		.INIT('h9)
	) name11922 (
		_w11920_,
		_w11955_,
		_w11956_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11923 (
		_w3710_,
		_w11408_,
		_w11463_,
		_w11464_,
		_w11957_
	);
	LUT4 #(
		.INIT('h2228)
	) name11924 (
		_w3886_,
		_w9446_,
		_w9702_,
		_w11261_,
		_w11958_
	);
	LUT3 #(
		.INIT('h82)
	) name11925 (
		_w3709_,
		_w11256_,
		_w11258_,
		_w11959_
	);
	LUT3 #(
		.INIT('h07)
	) name11926 (
		_w3877_,
		_w11406_,
		_w11959_,
		_w11960_
	);
	LUT2 #(
		.INIT('h4)
	) name11927 (
		_w11958_,
		_w11960_,
		_w11961_
	);
	LUT4 #(
		.INIT('h4844)
	) name11928 (
		\a[17] ,
		_w11956_,
		_w11957_,
		_w11961_,
		_w11962_
	);
	LUT4 #(
		.INIT('h9699)
	) name11929 (
		\a[17] ,
		_w11956_,
		_w11957_,
		_w11961_,
		_w11963_
	);
	LUT4 #(
		.INIT('h2b00)
	) name11930 (
		_w11795_,
		_w11800_,
		_w11917_,
		_w11963_,
		_w11964_
	);
	LUT4 #(
		.INIT('h54ab)
	) name11931 (
		_w11801_,
		_w11917_,
		_w11918_,
		_w11963_,
		_w11965_
	);
	LUT4 #(
		.INIT('h6500)
	) name11932 (
		\a[14] ,
		_w11564_,
		_w11568_,
		_w11965_,
		_w11966_
	);
	LUT4 #(
		.INIT('h54ab)
	) name11933 (
		_w11404_,
		_w11465_,
		_w11466_,
		_w11468_,
		_w11967_
	);
	LUT4 #(
		.INIT('h2228)
	) name11934 (
		_w4033_,
		_w9446_,
		_w9702_,
		_w11261_,
		_w11968_
	);
	LUT4 #(
		.INIT('h007d)
	) name11935 (
		_w4367_,
		_w11262_,
		_w11264_,
		_w11968_,
		_w11969_
	);
	LUT3 #(
		.INIT('h70)
	) name11936 (
		_w4382_,
		_w11400_,
		_w11969_,
		_w11970_
	);
	LUT4 #(
		.INIT('h95aa)
	) name11937 (
		\a[14] ,
		_w4034_,
		_w11967_,
		_w11970_,
		_w11971_
	);
	LUT2 #(
		.INIT('h9)
	) name11938 (
		_w11917_,
		_w11919_,
		_w11972_
	);
	LUT2 #(
		.INIT('h4)
	) name11939 (
		_w11971_,
		_w11972_,
		_w11973_
	);
	LUT2 #(
		.INIT('h9)
	) name11940 (
		_w11914_,
		_w11916_,
		_w11974_
	);
	LUT3 #(
		.INIT('h82)
	) name11941 (
		_w4034_,
		_w11465_,
		_w11467_,
		_w11975_
	);
	LUT3 #(
		.INIT('h82)
	) name11942 (
		_w4382_,
		_w11262_,
		_w11264_,
		_w11976_
	);
	LUT2 #(
		.INIT('h8)
	) name11943 (
		_w4033_,
		_w11406_,
		_w11977_
	);
	LUT4 #(
		.INIT('h2228)
	) name11944 (
		_w4367_,
		_w9446_,
		_w9702_,
		_w11261_,
		_w11978_
	);
	LUT2 #(
		.INIT('h1)
	) name11945 (
		_w11977_,
		_w11978_,
		_w11979_
	);
	LUT2 #(
		.INIT('h4)
	) name11946 (
		_w11976_,
		_w11979_,
		_w11980_
	);
	LUT4 #(
		.INIT('h4844)
	) name11947 (
		\a[14] ,
		_w11974_,
		_w11975_,
		_w11980_,
		_w11981_
	);
	LUT2 #(
		.INIT('h9)
	) name11948 (
		_w11911_,
		_w11913_,
		_w11982_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11949 (
		_w4034_,
		_w11408_,
		_w11463_,
		_w11464_,
		_w11983_
	);
	LUT4 #(
		.INIT('h2228)
	) name11950 (
		_w4382_,
		_w9446_,
		_w9702_,
		_w11261_,
		_w11984_
	);
	LUT3 #(
		.INIT('h82)
	) name11951 (
		_w4033_,
		_w11256_,
		_w11258_,
		_w11985_
	);
	LUT3 #(
		.INIT('h07)
	) name11952 (
		_w4367_,
		_w11406_,
		_w11985_,
		_w11986_
	);
	LUT2 #(
		.INIT('h4)
	) name11953 (
		_w11984_,
		_w11986_,
		_w11987_
	);
	LUT4 #(
		.INIT('h4844)
	) name11954 (
		\a[14] ,
		_w11982_,
		_w11983_,
		_w11987_,
		_w11988_
	);
	LUT2 #(
		.INIT('h9)
	) name11955 (
		_w11908_,
		_w11910_,
		_w11989_
	);
	LUT3 #(
		.INIT('h82)
	) name11956 (
		_w4033_,
		_w10268_,
		_w11255_,
		_w11990_
	);
	LUT4 #(
		.INIT('h007d)
	) name11957 (
		_w4367_,
		_w11256_,
		_w11258_,
		_w11990_,
		_w11991_
	);
	LUT3 #(
		.INIT('h70)
	) name11958 (
		_w4382_,
		_w11406_,
		_w11991_,
		_w11992_
	);
	LUT4 #(
		.INIT('h95aa)
	) name11959 (
		\a[14] ,
		_w4034_,
		_w11796_,
		_w11992_,
		_w11993_
	);
	LUT2 #(
		.INIT('h2)
	) name11960 (
		_w11989_,
		_w11993_,
		_w11994_
	);
	LUT3 #(
		.INIT('h82)
	) name11961 (
		_w4033_,
		_w10580_,
		_w11254_,
		_w11995_
	);
	LUT4 #(
		.INIT('h007d)
	) name11962 (
		_w4367_,
		_w10268_,
		_w11255_,
		_w11995_,
		_w11996_
	);
	LUT4 #(
		.INIT('h7d00)
	) name11963 (
		_w4382_,
		_w11256_,
		_w11258_,
		_w11996_,
		_w11997_
	);
	LUT4 #(
		.INIT('h7d00)
	) name11964 (
		_w4034_,
		_w11459_,
		_w11461_,
		_w11997_,
		_w11998_
	);
	LUT2 #(
		.INIT('h9)
	) name11965 (
		_w11905_,
		_w11907_,
		_w11999_
	);
	LUT3 #(
		.INIT('h90)
	) name11966 (
		\a[14] ,
		_w11998_,
		_w11999_,
		_w12000_
	);
	LUT3 #(
		.INIT('h82)
	) name11967 (
		_w4033_,
		_w10599_,
		_w11253_,
		_w12001_
	);
	LUT4 #(
		.INIT('h007d)
	) name11968 (
		_w4367_,
		_w10580_,
		_w11254_,
		_w12001_,
		_w12002_
	);
	LUT4 #(
		.INIT('h7d00)
	) name11969 (
		_w4382_,
		_w10268_,
		_w11255_,
		_w12002_,
		_w12003_
	);
	LUT4 #(
		.INIT('h7d00)
	) name11970 (
		_w4034_,
		_w11456_,
		_w11458_,
		_w12003_,
		_w12004_
	);
	LUT2 #(
		.INIT('h9)
	) name11971 (
		_w11902_,
		_w11904_,
		_w12005_
	);
	LUT3 #(
		.INIT('h90)
	) name11972 (
		\a[14] ,
		_w12004_,
		_w12005_,
		_w12006_
	);
	LUT2 #(
		.INIT('h8)
	) name11973 (
		_w4033_,
		_w11415_,
		_w12007_
	);
	LUT4 #(
		.INIT('h007d)
	) name11974 (
		_w4367_,
		_w10599_,
		_w11253_,
		_w12007_,
		_w12008_
	);
	LUT4 #(
		.INIT('h7d00)
	) name11975 (
		_w4382_,
		_w10580_,
		_w11254_,
		_w12008_,
		_w12009_
	);
	LUT4 #(
		.INIT('h7d00)
	) name11976 (
		_w4034_,
		_w11453_,
		_w11455_,
		_w12009_,
		_w12010_
	);
	LUT3 #(
		.INIT('h1e)
	) name11977 (
		_w11846_,
		_w11900_,
		_w11901_,
		_w12011_
	);
	LUT3 #(
		.INIT('h90)
	) name11978 (
		\a[14] ,
		_w12010_,
		_w12011_,
		_w12012_
	);
	LUT4 #(
		.INIT('h54ab)
	) name11979 (
		_w11852_,
		_w11896_,
		_w11897_,
		_w11899_,
		_w12013_
	);
	LUT3 #(
		.INIT('h82)
	) name11980 (
		_w4033_,
		_w11249_,
		_w11251_,
		_w12014_
	);
	LUT3 #(
		.INIT('h07)
	) name11981 (
		_w4367_,
		_w11415_,
		_w12014_,
		_w12015_
	);
	LUT4 #(
		.INIT('h7d00)
	) name11982 (
		_w4382_,
		_w10599_,
		_w11253_,
		_w12015_,
		_w12016_
	);
	LUT4 #(
		.INIT('h7d00)
	) name11983 (
		_w4034_,
		_w11450_,
		_w11452_,
		_w12016_,
		_w12017_
	);
	LUT3 #(
		.INIT('h84)
	) name11984 (
		\a[14] ,
		_w12013_,
		_w12017_,
		_w12018_
	);
	LUT2 #(
		.INIT('h9)
	) name11985 (
		_w11896_,
		_w11898_,
		_w12019_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11986 (
		_w4033_,
		_w10945_,
		_w11246_,
		_w11248_,
		_w12020_
	);
	LUT4 #(
		.INIT('h007d)
	) name11987 (
		_w4367_,
		_w11249_,
		_w11251_,
		_w12020_,
		_w12021_
	);
	LUT3 #(
		.INIT('h70)
	) name11988 (
		_w4382_,
		_w11415_,
		_w12021_,
		_w12022_
	);
	LUT4 #(
		.INIT('h95aa)
	) name11989 (
		\a[14] ,
		_w4034_,
		_w11675_,
		_w12022_,
		_w12023_
	);
	LUT2 #(
		.INIT('h2)
	) name11990 (
		_w12019_,
		_w12023_,
		_w12024_
	);
	LUT2 #(
		.INIT('h9)
	) name11991 (
		_w11893_,
		_w11895_,
		_w12025_
	);
	LUT3 #(
		.INIT('h82)
	) name11992 (
		_w4034_,
		_w11445_,
		_w11447_,
		_w12026_
	);
	LUT3 #(
		.INIT('h82)
	) name11993 (
		_w4382_,
		_w11249_,
		_w11251_,
		_w12027_
	);
	LUT2 #(
		.INIT('h8)
	) name11994 (
		_w4033_,
		_w11421_,
		_w12028_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11995 (
		_w4367_,
		_w10945_,
		_w11246_,
		_w11248_,
		_w12029_
	);
	LUT2 #(
		.INIT('h1)
	) name11996 (
		_w12028_,
		_w12029_,
		_w12030_
	);
	LUT2 #(
		.INIT('h4)
	) name11997 (
		_w12027_,
		_w12030_,
		_w12031_
	);
	LUT4 #(
		.INIT('h4844)
	) name11998 (
		\a[14] ,
		_w12025_,
		_w12026_,
		_w12031_,
		_w12032_
	);
	LUT4 #(
		.INIT('h02a8)
	) name11999 (
		_w4034_,
		_w11423_,
		_w11443_,
		_w11444_,
		_w12033_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12000 (
		_w4382_,
		_w10945_,
		_w11246_,
		_w11248_,
		_w12034_
	);
	LUT3 #(
		.INIT('h82)
	) name12001 (
		_w4033_,
		_w11241_,
		_w11243_,
		_w12035_
	);
	LUT3 #(
		.INIT('h07)
	) name12002 (
		_w4367_,
		_w11421_,
		_w12035_,
		_w12036_
	);
	LUT2 #(
		.INIT('h4)
	) name12003 (
		_w12034_,
		_w12036_,
		_w12037_
	);
	LUT2 #(
		.INIT('h9)
	) name12004 (
		_w11890_,
		_w11892_,
		_w12038_
	);
	LUT4 #(
		.INIT('h6500)
	) name12005 (
		\a[14] ,
		_w12033_,
		_w12037_,
		_w12038_,
		_w12039_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12006 (
		_w4033_,
		_w10968_,
		_w11238_,
		_w11240_,
		_w12040_
	);
	LUT4 #(
		.INIT('h007d)
	) name12007 (
		_w4367_,
		_w11241_,
		_w11243_,
		_w12040_,
		_w12041_
	);
	LUT3 #(
		.INIT('h70)
	) name12008 (
		_w4382_,
		_w11421_,
		_w12041_,
		_w12042_
	);
	LUT4 #(
		.INIT('h95aa)
	) name12009 (
		\a[14] ,
		_w4034_,
		_w11569_,
		_w12042_,
		_w12043_
	);
	LUT2 #(
		.INIT('h9)
	) name12010 (
		_w11887_,
		_w11889_,
		_w12044_
	);
	LUT2 #(
		.INIT('h4)
	) name12011 (
		_w12043_,
		_w12044_,
		_w12045_
	);
	LUT3 #(
		.INIT('h82)
	) name12012 (
		_w4034_,
		_w11439_,
		_w11441_,
		_w12046_
	);
	LUT3 #(
		.INIT('h82)
	) name12013 (
		_w4382_,
		_w11241_,
		_w11243_,
		_w12047_
	);
	LUT2 #(
		.INIT('h8)
	) name12014 (
		_w4033_,
		_w11427_,
		_w12048_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12015 (
		_w4367_,
		_w10968_,
		_w11238_,
		_w11240_,
		_w12049_
	);
	LUT2 #(
		.INIT('h1)
	) name12016 (
		_w12048_,
		_w12049_,
		_w12050_
	);
	LUT2 #(
		.INIT('h4)
	) name12017 (
		_w12047_,
		_w12050_,
		_w12051_
	);
	LUT3 #(
		.INIT('h8a)
	) name12018 (
		\a[17] ,
		_w11873_,
		_w11872_,
		_w12052_
	);
	LUT2 #(
		.INIT('h9)
	) name12019 (
		_w11881_,
		_w12052_,
		_w12053_
	);
	LUT4 #(
		.INIT('h6500)
	) name12020 (
		\a[14] ,
		_w12046_,
		_w12051_,
		_w12053_,
		_w12054_
	);
	LUT3 #(
		.INIT('h82)
	) name12021 (
		_w4034_,
		_w11436_,
		_w11438_,
		_w12055_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12022 (
		_w4382_,
		_w10968_,
		_w11238_,
		_w11240_,
		_w12056_
	);
	LUT3 #(
		.INIT('h82)
	) name12023 (
		_w4033_,
		_w11233_,
		_w11235_,
		_w12057_
	);
	LUT3 #(
		.INIT('h07)
	) name12024 (
		_w4367_,
		_w11427_,
		_w12057_,
		_w12058_
	);
	LUT2 #(
		.INIT('h4)
	) name12025 (
		_w12056_,
		_w12058_,
		_w12059_
	);
	LUT3 #(
		.INIT('h20)
	) name12026 (
		\a[17] ,
		_w3708_,
		_w11434_,
		_w12060_
	);
	LUT2 #(
		.INIT('h9)
	) name12027 (
		_w11872_,
		_w12060_,
		_w12061_
	);
	LUT4 #(
		.INIT('h6500)
	) name12028 (
		\a[14] ,
		_w12055_,
		_w12059_,
		_w12061_,
		_w12062_
	);
	LUT2 #(
		.INIT('h8)
	) name12029 (
		_w4367_,
		_w11434_,
		_w12063_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12030 (
		_w4382_,
		_w10991_,
		_w11230_,
		_w11232_,
		_w12064_
	);
	LUT4 #(
		.INIT('h000d)
	) name12031 (
		_w4034_,
		_w11581_,
		_w12063_,
		_w12064_,
		_w12065_
	);
	LUT2 #(
		.INIT('h4)
	) name12032 (
		_w4032_,
		_w11434_,
		_w12066_
	);
	LUT3 #(
		.INIT('h8a)
	) name12033 (
		\a[14] ,
		_w4032_,
		_w11434_,
		_w12067_
	);
	LUT2 #(
		.INIT('h8)
	) name12034 (
		_w12065_,
		_w12067_,
		_w12068_
	);
	LUT4 #(
		.INIT('h2882)
	) name12035 (
		_w4034_,
		_w11233_,
		_w11235_,
		_w11580_,
		_w12069_
	);
	LUT3 #(
		.INIT('h82)
	) name12036 (
		_w4382_,
		_w11233_,
		_w11235_,
		_w12070_
	);
	LUT2 #(
		.INIT('h8)
	) name12037 (
		_w4033_,
		_w11434_,
		_w12071_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12038 (
		_w4367_,
		_w10991_,
		_w11230_,
		_w11232_,
		_w12072_
	);
	LUT2 #(
		.INIT('h1)
	) name12039 (
		_w12071_,
		_w12072_,
		_w12073_
	);
	LUT3 #(
		.INIT('h10)
	) name12040 (
		_w12070_,
		_w12069_,
		_w12073_,
		_w12074_
	);
	LUT3 #(
		.INIT('h80)
	) name12041 (
		_w11873_,
		_w12068_,
		_w12074_,
		_w12075_
	);
	LUT3 #(
		.INIT('h28)
	) name12042 (
		_w4034_,
		_w11431_,
		_w11435_,
		_w12076_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12043 (
		_w4033_,
		_w10991_,
		_w11230_,
		_w11232_,
		_w12077_
	);
	LUT4 #(
		.INIT('h007d)
	) name12044 (
		_w4367_,
		_w11233_,
		_w11235_,
		_w12077_,
		_w12078_
	);
	LUT3 #(
		.INIT('h70)
	) name12045 (
		_w4382_,
		_w11427_,
		_w12078_,
		_w12079_
	);
	LUT3 #(
		.INIT('h9a)
	) name12046 (
		\a[14] ,
		_w12076_,
		_w12079_,
		_w12080_
	);
	LUT3 #(
		.INIT('h15)
	) name12047 (
		_w11873_,
		_w12068_,
		_w12074_,
		_w12081_
	);
	LUT3 #(
		.INIT('h6a)
	) name12048 (
		_w11873_,
		_w12068_,
		_w12074_,
		_w12082_
	);
	LUT3 #(
		.INIT('h54)
	) name12049 (
		_w12075_,
		_w12080_,
		_w12081_,
		_w12083_
	);
	LUT4 #(
		.INIT('h009a)
	) name12050 (
		\a[14] ,
		_w12055_,
		_w12059_,
		_w12061_,
		_w12084_
	);
	LUT4 #(
		.INIT('h9a65)
	) name12051 (
		\a[14] ,
		_w12055_,
		_w12059_,
		_w12061_,
		_w12085_
	);
	LUT3 #(
		.INIT('h54)
	) name12052 (
		_w12062_,
		_w12083_,
		_w12084_,
		_w12086_
	);
	LUT4 #(
		.INIT('h009a)
	) name12053 (
		\a[14] ,
		_w12046_,
		_w12051_,
		_w12053_,
		_w12087_
	);
	LUT4 #(
		.INIT('h9a65)
	) name12054 (
		\a[14] ,
		_w12046_,
		_w12051_,
		_w12053_,
		_w12088_
	);
	LUT3 #(
		.INIT('h54)
	) name12055 (
		_w12054_,
		_w12086_,
		_w12087_,
		_w12089_
	);
	LUT2 #(
		.INIT('h2)
	) name12056 (
		_w12043_,
		_w12044_,
		_w12090_
	);
	LUT2 #(
		.INIT('h9)
	) name12057 (
		_w12043_,
		_w12044_,
		_w12091_
	);
	LUT4 #(
		.INIT('h9a65)
	) name12058 (
		\a[14] ,
		_w12033_,
		_w12037_,
		_w12038_,
		_w12092_
	);
	LUT4 #(
		.INIT('h4d00)
	) name12059 (
		_w12043_,
		_w12044_,
		_w12089_,
		_w12092_,
		_w12093_
	);
	LUT4 #(
		.INIT('h9699)
	) name12060 (
		\a[14] ,
		_w12025_,
		_w12026_,
		_w12031_,
		_w12094_
	);
	LUT4 #(
		.INIT('h0155)
	) name12061 (
		_w12032_,
		_w12039_,
		_w12093_,
		_w12094_,
		_w12095_
	);
	LUT2 #(
		.INIT('h4)
	) name12062 (
		_w12019_,
		_w12023_,
		_w12096_
	);
	LUT2 #(
		.INIT('h9)
	) name12063 (
		_w12019_,
		_w12023_,
		_w12097_
	);
	LUT3 #(
		.INIT('h54)
	) name12064 (
		_w12024_,
		_w12095_,
		_w12096_,
		_w12098_
	);
	LUT3 #(
		.INIT('h12)
	) name12065 (
		\a[14] ,
		_w12013_,
		_w12017_,
		_w12099_
	);
	LUT3 #(
		.INIT('h69)
	) name12066 (
		\a[14] ,
		_w12013_,
		_w12017_,
		_w12100_
	);
	LUT3 #(
		.INIT('h54)
	) name12067 (
		_w12018_,
		_w12098_,
		_w12099_,
		_w12101_
	);
	LUT3 #(
		.INIT('h06)
	) name12068 (
		\a[14] ,
		_w12010_,
		_w12011_,
		_w12102_
	);
	LUT3 #(
		.INIT('h69)
	) name12069 (
		\a[14] ,
		_w12010_,
		_w12011_,
		_w12103_
	);
	LUT3 #(
		.INIT('h54)
	) name12070 (
		_w12012_,
		_w12101_,
		_w12102_,
		_w12104_
	);
	LUT3 #(
		.INIT('h06)
	) name12071 (
		\a[14] ,
		_w12004_,
		_w12005_,
		_w12105_
	);
	LUT3 #(
		.INIT('h69)
	) name12072 (
		\a[14] ,
		_w12004_,
		_w12005_,
		_w12106_
	);
	LUT3 #(
		.INIT('h54)
	) name12073 (
		_w12006_,
		_w12104_,
		_w12105_,
		_w12107_
	);
	LUT3 #(
		.INIT('h06)
	) name12074 (
		\a[14] ,
		_w11998_,
		_w11999_,
		_w12108_
	);
	LUT3 #(
		.INIT('h69)
	) name12075 (
		\a[14] ,
		_w11998_,
		_w11999_,
		_w12109_
	);
	LUT3 #(
		.INIT('h54)
	) name12076 (
		_w12000_,
		_w12107_,
		_w12108_,
		_w12110_
	);
	LUT2 #(
		.INIT('h4)
	) name12077 (
		_w11989_,
		_w11993_,
		_w12111_
	);
	LUT2 #(
		.INIT('h9)
	) name12078 (
		_w11989_,
		_w11993_,
		_w12112_
	);
	LUT4 #(
		.INIT('h9699)
	) name12079 (
		\a[14] ,
		_w11982_,
		_w11983_,
		_w11987_,
		_w12113_
	);
	LUT4 #(
		.INIT('h2b00)
	) name12080 (
		_w11989_,
		_w11993_,
		_w12110_,
		_w12113_,
		_w12114_
	);
	LUT4 #(
		.INIT('h9699)
	) name12081 (
		\a[14] ,
		_w11974_,
		_w11975_,
		_w11980_,
		_w12115_
	);
	LUT4 #(
		.INIT('h0155)
	) name12082 (
		_w11981_,
		_w11988_,
		_w12114_,
		_w12115_,
		_w12116_
	);
	LUT2 #(
		.INIT('h2)
	) name12083 (
		_w11971_,
		_w11972_,
		_w12117_
	);
	LUT2 #(
		.INIT('h9)
	) name12084 (
		_w11971_,
		_w11972_,
		_w12118_
	);
	LUT4 #(
		.INIT('h9a65)
	) name12085 (
		\a[14] ,
		_w11564_,
		_w11568_,
		_w11965_,
		_w12119_
	);
	LUT4 #(
		.INIT('h4d00)
	) name12086 (
		_w11971_,
		_w11972_,
		_w12116_,
		_w12119_,
		_w12120_
	);
	LUT3 #(
		.INIT('h82)
	) name12087 (
		_w3710_,
		_w11465_,
		_w11467_,
		_w12121_
	);
	LUT3 #(
		.INIT('h82)
	) name12088 (
		_w3886_,
		_w11262_,
		_w11264_,
		_w12122_
	);
	LUT2 #(
		.INIT('h8)
	) name12089 (
		_w3709_,
		_w11406_,
		_w12123_
	);
	LUT4 #(
		.INIT('h2228)
	) name12090 (
		_w3877_,
		_w9446_,
		_w9702_,
		_w11261_,
		_w12124_
	);
	LUT2 #(
		.INIT('h1)
	) name12091 (
		_w12123_,
		_w12124_,
		_w12125_
	);
	LUT2 #(
		.INIT('h4)
	) name12092 (
		_w12122_,
		_w12125_,
		_w12126_
	);
	LUT3 #(
		.INIT('h32)
	) name12093 (
		_w11920_,
		_w11953_,
		_w11954_,
		_w12127_
	);
	LUT3 #(
		.INIT('h32)
	) name12094 (
		_w11925_,
		_w11949_,
		_w11950_,
		_w12128_
	);
	LUT3 #(
		.INIT('h82)
	) name12095 (
		_w3214_,
		_w11249_,
		_w11251_,
		_w12129_
	);
	LUT3 #(
		.INIT('h07)
	) name12096 (
		_w3249_,
		_w11415_,
		_w12129_,
		_w12130_
	);
	LUT4 #(
		.INIT('h7d00)
	) name12097 (
		_w3262_,
		_w10599_,
		_w11253_,
		_w12130_,
		_w12131_
	);
	LUT4 #(
		.INIT('h7d00)
	) name12098 (
		_w37_,
		_w11450_,
		_w11452_,
		_w12131_,
		_w12132_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12099 (
		_w2875_,
		_w11423_,
		_w11443_,
		_w11444_,
		_w12133_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12100 (
		_w2986_,
		_w10945_,
		_w11246_,
		_w11248_,
		_w12134_
	);
	LUT3 #(
		.INIT('h82)
	) name12101 (
		_w2874_,
		_w11241_,
		_w11243_,
		_w12135_
	);
	LUT3 #(
		.INIT('h07)
	) name12102 (
		_w2975_,
		_w11421_,
		_w12135_,
		_w12136_
	);
	LUT2 #(
		.INIT('h4)
	) name12103 (
		_w12134_,
		_w12136_,
		_w12137_
	);
	LUT3 #(
		.INIT('h32)
	) name12104 (
		_w11935_,
		_w11937_,
		_w11938_,
		_w12138_
	);
	LUT3 #(
		.INIT('h82)
	) name12105 (
		_w2550_,
		_w11436_,
		_w11438_,
		_w12139_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12106 (
		_w2854_,
		_w10968_,
		_w11238_,
		_w11240_,
		_w12140_
	);
	LUT3 #(
		.INIT('h82)
	) name12107 (
		_w2549_,
		_w11233_,
		_w11235_,
		_w12141_
	);
	LUT3 #(
		.INIT('h07)
	) name12108 (
		_w2617_,
		_w11427_,
		_w12141_,
		_w12142_
	);
	LUT2 #(
		.INIT('h4)
	) name12109 (
		_w12140_,
		_w12142_,
		_w12143_
	);
	LUT3 #(
		.INIT('h80)
	) name12110 (
		_w950_,
		_w1198_,
		_w3350_,
		_w12144_
	);
	LUT4 #(
		.INIT('h0777)
	) name12111 (
		_w59_,
		_w43_,
		_w44_,
		_w201_,
		_w12145_
	);
	LUT2 #(
		.INIT('h4)
	) name12112 (
		_w165_,
		_w12145_,
		_w12146_
	);
	LUT4 #(
		.INIT('h8000)
	) name12113 (
		_w287_,
		_w807_,
		_w817_,
		_w860_,
		_w12147_
	);
	LUT3 #(
		.INIT('h80)
	) name12114 (
		_w12146_,
		_w12144_,
		_w12147_,
		_w12148_
	);
	LUT4 #(
		.INIT('h0777)
	) name12115 (
		_w85_,
		_w43_,
		_w46_,
		_w259_,
		_w12149_
	);
	LUT4 #(
		.INIT('h4000)
	) name12116 (
		_w268_,
		_w777_,
		_w894_,
		_w12149_,
		_w12150_
	);
	LUT4 #(
		.INIT('h8000)
	) name12117 (
		_w678_,
		_w1113_,
		_w1910_,
		_w1911_,
		_w12151_
	);
	LUT2 #(
		.INIT('h8)
	) name12118 (
		_w12150_,
		_w12151_,
		_w12152_
	);
	LUT4 #(
		.INIT('h8000)
	) name12119 (
		_w944_,
		_w1318_,
		_w1359_,
		_w2581_,
		_w12153_
	);
	LUT3 #(
		.INIT('h80)
	) name12120 (
		_w1279_,
		_w8306_,
		_w12153_,
		_w12154_
	);
	LUT3 #(
		.INIT('h80)
	) name12121 (
		_w12148_,
		_w12152_,
		_w12154_,
		_w12155_
	);
	LUT4 #(
		.INIT('h153f)
	) name12122 (
		_w85_,
		_w56_,
		_w158_,
		_w176_,
		_w12156_
	);
	LUT4 #(
		.INIT('h8000)
	) name12123 (
		_w125_,
		_w408_,
		_w411_,
		_w12156_,
		_w12157_
	);
	LUT2 #(
		.INIT('h8)
	) name12124 (
		_w3018_,
		_w12157_,
		_w12158_
	);
	LUT4 #(
		.INIT('h8000)
	) name12125 (
		_w1982_,
		_w2256_,
		_w2706_,
		_w4266_,
		_w12159_
	);
	LUT4 #(
		.INIT('h8000)
	) name12126 (
		_w387_,
		_w820_,
		_w908_,
		_w1158_,
		_w12160_
	);
	LUT3 #(
		.INIT('h80)
	) name12127 (
		_w7438_,
		_w12159_,
		_w12160_,
		_w12161_
	);
	LUT4 #(
		.INIT('h8000)
	) name12128 (
		_w4193_,
		_w8267_,
		_w12158_,
		_w12161_,
		_w12162_
	);
	LUT2 #(
		.INIT('h8)
	) name12129 (
		_w12155_,
		_w12162_,
		_w12163_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12130 (
		_w2527_,
		_w10991_,
		_w11230_,
		_w11232_,
		_w12164_
	);
	LUT2 #(
		.INIT('h8)
	) name12131 (
		_w2407_,
		_w11434_,
		_w12165_
	);
	LUT4 #(
		.INIT('h000d)
	) name12132 (
		_w377_,
		_w11581_,
		_w12164_,
		_w12165_,
		_w12166_
	);
	LUT2 #(
		.INIT('h6)
	) name12133 (
		_w12163_,
		_w12166_,
		_w12167_
	);
	LUT4 #(
		.INIT('h6500)
	) name12134 (
		\a[29] ,
		_w12139_,
		_w12143_,
		_w12167_,
		_w12168_
	);
	LUT4 #(
		.INIT('h009a)
	) name12135 (
		\a[29] ,
		_w12139_,
		_w12143_,
		_w12167_,
		_w12169_
	);
	LUT4 #(
		.INIT('h9a65)
	) name12136 (
		\a[29] ,
		_w12139_,
		_w12143_,
		_w12167_,
		_w12170_
	);
	LUT2 #(
		.INIT('h9)
	) name12137 (
		_w12138_,
		_w12170_,
		_w12171_
	);
	LUT4 #(
		.INIT('h6500)
	) name12138 (
		\a[26] ,
		_w12133_,
		_w12137_,
		_w12171_,
		_w12172_
	);
	LUT4 #(
		.INIT('h9a65)
	) name12139 (
		\a[26] ,
		_w12133_,
		_w12137_,
		_w12171_,
		_w12173_
	);
	LUT4 #(
		.INIT('h7100)
	) name12140 (
		_w11926_,
		_w11930_,
		_w11940_,
		_w12173_,
		_w12174_
	);
	LUT4 #(
		.INIT('h32cd)
	) name12141 (
		_w11926_,
		_w11941_,
		_w11942_,
		_w12173_,
		_w12175_
	);
	LUT3 #(
		.INIT('h90)
	) name12142 (
		\a[23] ,
		_w12132_,
		_w12175_,
		_w12176_
	);
	LUT3 #(
		.INIT('h06)
	) name12143 (
		\a[23] ,
		_w12132_,
		_w12175_,
		_w12177_
	);
	LUT3 #(
		.INIT('h69)
	) name12144 (
		\a[23] ,
		_w12132_,
		_w12175_,
		_w12178_
	);
	LUT2 #(
		.INIT('h9)
	) name12145 (
		_w12128_,
		_w12178_,
		_w12179_
	);
	LUT3 #(
		.INIT('h82)
	) name12146 (
		_w3311_,
		_w10580_,
		_w11254_,
		_w12180_
	);
	LUT4 #(
		.INIT('h007d)
	) name12147 (
		_w3645_,
		_w10268_,
		_w11255_,
		_w12180_,
		_w12181_
	);
	LUT4 #(
		.INIT('h7d00)
	) name12148 (
		_w3654_,
		_w11256_,
		_w11258_,
		_w12181_,
		_w12182_
	);
	LUT4 #(
		.INIT('h7d00)
	) name12149 (
		_w3312_,
		_w11459_,
		_w11461_,
		_w12182_,
		_w12183_
	);
	LUT3 #(
		.INIT('h84)
	) name12150 (
		\a[20] ,
		_w12179_,
		_w12183_,
		_w12184_
	);
	LUT3 #(
		.INIT('h12)
	) name12151 (
		\a[20] ,
		_w12179_,
		_w12183_,
		_w12185_
	);
	LUT3 #(
		.INIT('h69)
	) name12152 (
		\a[20] ,
		_w12179_,
		_w12183_,
		_w12186_
	);
	LUT2 #(
		.INIT('h9)
	) name12153 (
		_w12127_,
		_w12186_,
		_w12187_
	);
	LUT4 #(
		.INIT('h6500)
	) name12154 (
		\a[17] ,
		_w12121_,
		_w12126_,
		_w12187_,
		_w12188_
	);
	LUT4 #(
		.INIT('h9a65)
	) name12155 (
		\a[17] ,
		_w12121_,
		_w12126_,
		_w12187_,
		_w12189_
	);
	LUT3 #(
		.INIT('h1e)
	) name12156 (
		_w11962_,
		_w11964_,
		_w12189_,
		_w12190_
	);
	LUT3 #(
		.INIT('h82)
	) name12157 (
		_w4034_,
		_w11472_,
		_w11474_,
		_w12191_
	);
	LUT3 #(
		.INIT('h82)
	) name12158 (
		_w4382_,
		_w11268_,
		_w11270_,
		_w12192_
	);
	LUT2 #(
		.INIT('h8)
	) name12159 (
		_w4033_,
		_w11400_,
		_w12193_
	);
	LUT4 #(
		.INIT('h2228)
	) name12160 (
		_w4367_,
		_w8794_,
		_w8994_,
		_w11267_,
		_w12194_
	);
	LUT2 #(
		.INIT('h1)
	) name12161 (
		_w12193_,
		_w12194_,
		_w12195_
	);
	LUT2 #(
		.INIT('h4)
	) name12162 (
		_w12192_,
		_w12195_,
		_w12196_
	);
	LUT4 #(
		.INIT('h4844)
	) name12163 (
		\a[14] ,
		_w12190_,
		_w12191_,
		_w12196_,
		_w12197_
	);
	LUT4 #(
		.INIT('h9699)
	) name12164 (
		\a[14] ,
		_w12190_,
		_w12191_,
		_w12196_,
		_w12198_
	);
	LUT3 #(
		.INIT('h1e)
	) name12165 (
		_w11966_,
		_w12120_,
		_w12198_,
		_w12199_
	);
	LUT4 #(
		.INIT('h6500)
	) name12166 (
		\a[11] ,
		_w11558_,
		_w11563_,
		_w12199_,
		_w12200_
	);
	LUT4 #(
		.INIT('h54ab)
	) name12167 (
		_w11973_,
		_w12116_,
		_w12117_,
		_w12119_,
		_w12201_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12168 (
		_w4459_,
		_w11396_,
		_w11476_,
		_w11477_,
		_w12202_
	);
	LUT4 #(
		.INIT('h2228)
	) name12169 (
		_w4700_,
		_w8466_,
		_w8541_,
		_w11273_,
		_w12203_
	);
	LUT3 #(
		.INIT('h82)
	) name12170 (
		_w4458_,
		_w11268_,
		_w11270_,
		_w12204_
	);
	LUT3 #(
		.INIT('h07)
	) name12171 (
		_w4684_,
		_w11394_,
		_w12204_,
		_w12205_
	);
	LUT2 #(
		.INIT('h4)
	) name12172 (
		_w12203_,
		_w12205_,
		_w12206_
	);
	LUT4 #(
		.INIT('h4844)
	) name12173 (
		\a[11] ,
		_w12201_,
		_w12202_,
		_w12206_,
		_w12207_
	);
	LUT2 #(
		.INIT('h9)
	) name12174 (
		_w12116_,
		_w12118_,
		_w12208_
	);
	LUT4 #(
		.INIT('h54ab)
	) name12175 (
		_w11398_,
		_w11472_,
		_w11473_,
		_w11475_,
		_w12209_
	);
	LUT4 #(
		.INIT('h2228)
	) name12176 (
		_w4458_,
		_w8794_,
		_w8994_,
		_w11267_,
		_w12210_
	);
	LUT4 #(
		.INIT('h007d)
	) name12177 (
		_w4684_,
		_w11268_,
		_w11270_,
		_w12210_,
		_w12211_
	);
	LUT3 #(
		.INIT('h70)
	) name12178 (
		_w4700_,
		_w11394_,
		_w12211_,
		_w12212_
	);
	LUT4 #(
		.INIT('h95aa)
	) name12179 (
		\a[11] ,
		_w4459_,
		_w12209_,
		_w12212_,
		_w12213_
	);
	LUT2 #(
		.INIT('h2)
	) name12180 (
		_w12208_,
		_w12213_,
		_w12214_
	);
	LUT3 #(
		.INIT('h82)
	) name12181 (
		_w4459_,
		_w11472_,
		_w11474_,
		_w12215_
	);
	LUT3 #(
		.INIT('h82)
	) name12182 (
		_w4700_,
		_w11268_,
		_w11270_,
		_w12216_
	);
	LUT2 #(
		.INIT('h8)
	) name12183 (
		_w4458_,
		_w11400_,
		_w12217_
	);
	LUT4 #(
		.INIT('h2228)
	) name12184 (
		_w4684_,
		_w8794_,
		_w8994_,
		_w11267_,
		_w12218_
	);
	LUT2 #(
		.INIT('h1)
	) name12185 (
		_w12217_,
		_w12218_,
		_w12219_
	);
	LUT2 #(
		.INIT('h4)
	) name12186 (
		_w12216_,
		_w12219_,
		_w12220_
	);
	LUT3 #(
		.INIT('h1e)
	) name12187 (
		_w11988_,
		_w12114_,
		_w12115_,
		_w12221_
	);
	LUT4 #(
		.INIT('h6500)
	) name12188 (
		\a[11] ,
		_w12215_,
		_w12220_,
		_w12221_,
		_w12222_
	);
	LUT3 #(
		.INIT('h82)
	) name12189 (
		_w4459_,
		_w11469_,
		_w11471_,
		_w12223_
	);
	LUT4 #(
		.INIT('h2228)
	) name12190 (
		_w4700_,
		_w8794_,
		_w8994_,
		_w11267_,
		_w12224_
	);
	LUT3 #(
		.INIT('h82)
	) name12191 (
		_w4458_,
		_w11262_,
		_w11264_,
		_w12225_
	);
	LUT3 #(
		.INIT('h07)
	) name12192 (
		_w4684_,
		_w11400_,
		_w12225_,
		_w12226_
	);
	LUT2 #(
		.INIT('h4)
	) name12193 (
		_w12224_,
		_w12226_,
		_w12227_
	);
	LUT4 #(
		.INIT('h54ab)
	) name12194 (
		_w11994_,
		_w12110_,
		_w12111_,
		_w12113_,
		_w12228_
	);
	LUT4 #(
		.INIT('h6500)
	) name12195 (
		\a[11] ,
		_w12223_,
		_w12227_,
		_w12228_,
		_w12229_
	);
	LUT4 #(
		.INIT('h2228)
	) name12196 (
		_w4458_,
		_w9446_,
		_w9702_,
		_w11261_,
		_w12230_
	);
	LUT4 #(
		.INIT('h007d)
	) name12197 (
		_w4684_,
		_w11262_,
		_w11264_,
		_w12230_,
		_w12231_
	);
	LUT3 #(
		.INIT('h70)
	) name12198 (
		_w4700_,
		_w11400_,
		_w12231_,
		_w12232_
	);
	LUT4 #(
		.INIT('h95aa)
	) name12199 (
		\a[11] ,
		_w4459_,
		_w11967_,
		_w12232_,
		_w12233_
	);
	LUT2 #(
		.INIT('h9)
	) name12200 (
		_w12110_,
		_w12112_,
		_w12234_
	);
	LUT2 #(
		.INIT('h4)
	) name12201 (
		_w12233_,
		_w12234_,
		_w12235_
	);
	LUT2 #(
		.INIT('h9)
	) name12202 (
		_w12107_,
		_w12109_,
		_w12236_
	);
	LUT3 #(
		.INIT('h82)
	) name12203 (
		_w4459_,
		_w11465_,
		_w11467_,
		_w12237_
	);
	LUT3 #(
		.INIT('h82)
	) name12204 (
		_w4700_,
		_w11262_,
		_w11264_,
		_w12238_
	);
	LUT2 #(
		.INIT('h8)
	) name12205 (
		_w4458_,
		_w11406_,
		_w12239_
	);
	LUT4 #(
		.INIT('h2228)
	) name12206 (
		_w4684_,
		_w9446_,
		_w9702_,
		_w11261_,
		_w12240_
	);
	LUT2 #(
		.INIT('h1)
	) name12207 (
		_w12239_,
		_w12240_,
		_w12241_
	);
	LUT2 #(
		.INIT('h4)
	) name12208 (
		_w12238_,
		_w12241_,
		_w12242_
	);
	LUT4 #(
		.INIT('h4844)
	) name12209 (
		\a[11] ,
		_w12236_,
		_w12237_,
		_w12242_,
		_w12243_
	);
	LUT2 #(
		.INIT('h9)
	) name12210 (
		_w12104_,
		_w12106_,
		_w12244_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12211 (
		_w4459_,
		_w11408_,
		_w11463_,
		_w11464_,
		_w12245_
	);
	LUT4 #(
		.INIT('h2228)
	) name12212 (
		_w4700_,
		_w9446_,
		_w9702_,
		_w11261_,
		_w12246_
	);
	LUT3 #(
		.INIT('h82)
	) name12213 (
		_w4458_,
		_w11256_,
		_w11258_,
		_w12247_
	);
	LUT3 #(
		.INIT('h07)
	) name12214 (
		_w4684_,
		_w11406_,
		_w12247_,
		_w12248_
	);
	LUT2 #(
		.INIT('h4)
	) name12215 (
		_w12246_,
		_w12248_,
		_w12249_
	);
	LUT4 #(
		.INIT('h4844)
	) name12216 (
		\a[11] ,
		_w12244_,
		_w12245_,
		_w12249_,
		_w12250_
	);
	LUT2 #(
		.INIT('h9)
	) name12217 (
		_w12101_,
		_w12103_,
		_w12251_
	);
	LUT3 #(
		.INIT('h82)
	) name12218 (
		_w4458_,
		_w10268_,
		_w11255_,
		_w12252_
	);
	LUT4 #(
		.INIT('h007d)
	) name12219 (
		_w4684_,
		_w11256_,
		_w11258_,
		_w12252_,
		_w12253_
	);
	LUT3 #(
		.INIT('h70)
	) name12220 (
		_w4700_,
		_w11406_,
		_w12253_,
		_w12254_
	);
	LUT4 #(
		.INIT('h95aa)
	) name12221 (
		\a[11] ,
		_w4459_,
		_w11796_,
		_w12254_,
		_w12255_
	);
	LUT2 #(
		.INIT('h2)
	) name12222 (
		_w12251_,
		_w12255_,
		_w12256_
	);
	LUT3 #(
		.INIT('h82)
	) name12223 (
		_w4458_,
		_w10580_,
		_w11254_,
		_w12257_
	);
	LUT4 #(
		.INIT('h007d)
	) name12224 (
		_w4684_,
		_w10268_,
		_w11255_,
		_w12257_,
		_w12258_
	);
	LUT4 #(
		.INIT('h7d00)
	) name12225 (
		_w4700_,
		_w11256_,
		_w11258_,
		_w12258_,
		_w12259_
	);
	LUT4 #(
		.INIT('h7d00)
	) name12226 (
		_w4459_,
		_w11459_,
		_w11461_,
		_w12259_,
		_w12260_
	);
	LUT2 #(
		.INIT('h9)
	) name12227 (
		_w12098_,
		_w12100_,
		_w12261_
	);
	LUT3 #(
		.INIT('h90)
	) name12228 (
		\a[11] ,
		_w12260_,
		_w12261_,
		_w12262_
	);
	LUT3 #(
		.INIT('h82)
	) name12229 (
		_w4458_,
		_w10599_,
		_w11253_,
		_w12263_
	);
	LUT4 #(
		.INIT('h007d)
	) name12230 (
		_w4684_,
		_w10580_,
		_w11254_,
		_w12263_,
		_w12264_
	);
	LUT4 #(
		.INIT('h7d00)
	) name12231 (
		_w4700_,
		_w10268_,
		_w11255_,
		_w12264_,
		_w12265_
	);
	LUT4 #(
		.INIT('h7d00)
	) name12232 (
		_w4459_,
		_w11456_,
		_w11458_,
		_w12265_,
		_w12266_
	);
	LUT2 #(
		.INIT('h9)
	) name12233 (
		_w12095_,
		_w12097_,
		_w12267_
	);
	LUT3 #(
		.INIT('h90)
	) name12234 (
		\a[11] ,
		_w12266_,
		_w12267_,
		_w12268_
	);
	LUT2 #(
		.INIT('h8)
	) name12235 (
		_w4458_,
		_w11415_,
		_w12269_
	);
	LUT4 #(
		.INIT('h007d)
	) name12236 (
		_w4684_,
		_w10599_,
		_w11253_,
		_w12269_,
		_w12270_
	);
	LUT4 #(
		.INIT('h7d00)
	) name12237 (
		_w4700_,
		_w10580_,
		_w11254_,
		_w12270_,
		_w12271_
	);
	LUT4 #(
		.INIT('h7d00)
	) name12238 (
		_w4459_,
		_w11453_,
		_w11455_,
		_w12271_,
		_w12272_
	);
	LUT3 #(
		.INIT('h1e)
	) name12239 (
		_w12039_,
		_w12093_,
		_w12094_,
		_w12273_
	);
	LUT3 #(
		.INIT('h90)
	) name12240 (
		\a[11] ,
		_w12272_,
		_w12273_,
		_w12274_
	);
	LUT4 #(
		.INIT('h54ab)
	) name12241 (
		_w12045_,
		_w12089_,
		_w12090_,
		_w12092_,
		_w12275_
	);
	LUT3 #(
		.INIT('h82)
	) name12242 (
		_w4458_,
		_w11249_,
		_w11251_,
		_w12276_
	);
	LUT3 #(
		.INIT('h07)
	) name12243 (
		_w4684_,
		_w11415_,
		_w12276_,
		_w12277_
	);
	LUT4 #(
		.INIT('h7d00)
	) name12244 (
		_w4700_,
		_w10599_,
		_w11253_,
		_w12277_,
		_w12278_
	);
	LUT4 #(
		.INIT('h7d00)
	) name12245 (
		_w4459_,
		_w11450_,
		_w11452_,
		_w12278_,
		_w12279_
	);
	LUT3 #(
		.INIT('h84)
	) name12246 (
		\a[11] ,
		_w12275_,
		_w12279_,
		_w12280_
	);
	LUT2 #(
		.INIT('h9)
	) name12247 (
		_w12089_,
		_w12091_,
		_w12281_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12248 (
		_w4458_,
		_w10945_,
		_w11246_,
		_w11248_,
		_w12282_
	);
	LUT4 #(
		.INIT('h007d)
	) name12249 (
		_w4684_,
		_w11249_,
		_w11251_,
		_w12282_,
		_w12283_
	);
	LUT3 #(
		.INIT('h70)
	) name12250 (
		_w4700_,
		_w11415_,
		_w12283_,
		_w12284_
	);
	LUT4 #(
		.INIT('h95aa)
	) name12251 (
		\a[11] ,
		_w4459_,
		_w11675_,
		_w12284_,
		_w12285_
	);
	LUT2 #(
		.INIT('h2)
	) name12252 (
		_w12281_,
		_w12285_,
		_w12286_
	);
	LUT2 #(
		.INIT('h9)
	) name12253 (
		_w12086_,
		_w12088_,
		_w12287_
	);
	LUT3 #(
		.INIT('h82)
	) name12254 (
		_w4459_,
		_w11445_,
		_w11447_,
		_w12288_
	);
	LUT3 #(
		.INIT('h82)
	) name12255 (
		_w4700_,
		_w11249_,
		_w11251_,
		_w12289_
	);
	LUT2 #(
		.INIT('h8)
	) name12256 (
		_w4458_,
		_w11421_,
		_w12290_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12257 (
		_w4684_,
		_w10945_,
		_w11246_,
		_w11248_,
		_w12291_
	);
	LUT2 #(
		.INIT('h1)
	) name12258 (
		_w12290_,
		_w12291_,
		_w12292_
	);
	LUT2 #(
		.INIT('h4)
	) name12259 (
		_w12289_,
		_w12292_,
		_w12293_
	);
	LUT4 #(
		.INIT('h4844)
	) name12260 (
		\a[11] ,
		_w12287_,
		_w12288_,
		_w12293_,
		_w12294_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12261 (
		_w4459_,
		_w11423_,
		_w11443_,
		_w11444_,
		_w12295_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12262 (
		_w4700_,
		_w10945_,
		_w11246_,
		_w11248_,
		_w12296_
	);
	LUT3 #(
		.INIT('h82)
	) name12263 (
		_w4458_,
		_w11241_,
		_w11243_,
		_w12297_
	);
	LUT3 #(
		.INIT('h07)
	) name12264 (
		_w4684_,
		_w11421_,
		_w12297_,
		_w12298_
	);
	LUT2 #(
		.INIT('h4)
	) name12265 (
		_w12296_,
		_w12298_,
		_w12299_
	);
	LUT2 #(
		.INIT('h9)
	) name12266 (
		_w12083_,
		_w12085_,
		_w12300_
	);
	LUT4 #(
		.INIT('h6500)
	) name12267 (
		\a[11] ,
		_w12295_,
		_w12299_,
		_w12300_,
		_w12301_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12268 (
		_w4458_,
		_w10968_,
		_w11238_,
		_w11240_,
		_w12302_
	);
	LUT4 #(
		.INIT('h007d)
	) name12269 (
		_w4684_,
		_w11241_,
		_w11243_,
		_w12302_,
		_w12303_
	);
	LUT3 #(
		.INIT('h70)
	) name12270 (
		_w4700_,
		_w11421_,
		_w12303_,
		_w12304_
	);
	LUT4 #(
		.INIT('h95aa)
	) name12271 (
		\a[11] ,
		_w4459_,
		_w11569_,
		_w12304_,
		_w12305_
	);
	LUT2 #(
		.INIT('h9)
	) name12272 (
		_w12080_,
		_w12082_,
		_w12306_
	);
	LUT2 #(
		.INIT('h4)
	) name12273 (
		_w12305_,
		_w12306_,
		_w12307_
	);
	LUT3 #(
		.INIT('h82)
	) name12274 (
		_w4459_,
		_w11439_,
		_w11441_,
		_w12308_
	);
	LUT3 #(
		.INIT('h82)
	) name12275 (
		_w4700_,
		_w11241_,
		_w11243_,
		_w12309_
	);
	LUT2 #(
		.INIT('h8)
	) name12276 (
		_w4458_,
		_w11427_,
		_w12310_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12277 (
		_w4684_,
		_w10968_,
		_w11238_,
		_w11240_,
		_w12311_
	);
	LUT2 #(
		.INIT('h1)
	) name12278 (
		_w12310_,
		_w12311_,
		_w12312_
	);
	LUT2 #(
		.INIT('h4)
	) name12279 (
		_w12309_,
		_w12312_,
		_w12313_
	);
	LUT3 #(
		.INIT('h8a)
	) name12280 (
		\a[14] ,
		_w12066_,
		_w12065_,
		_w12314_
	);
	LUT2 #(
		.INIT('h9)
	) name12281 (
		_w12074_,
		_w12314_,
		_w12315_
	);
	LUT4 #(
		.INIT('h6500)
	) name12282 (
		\a[11] ,
		_w12308_,
		_w12313_,
		_w12315_,
		_w12316_
	);
	LUT3 #(
		.INIT('h82)
	) name12283 (
		_w4459_,
		_w11436_,
		_w11438_,
		_w12317_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12284 (
		_w4700_,
		_w10968_,
		_w11238_,
		_w11240_,
		_w12318_
	);
	LUT3 #(
		.INIT('h82)
	) name12285 (
		_w4458_,
		_w11233_,
		_w11235_,
		_w12319_
	);
	LUT3 #(
		.INIT('h07)
	) name12286 (
		_w4684_,
		_w11427_,
		_w12319_,
		_w12320_
	);
	LUT2 #(
		.INIT('h4)
	) name12287 (
		_w12318_,
		_w12320_,
		_w12321_
	);
	LUT3 #(
		.INIT('h20)
	) name12288 (
		\a[14] ,
		_w4032_,
		_w11434_,
		_w12322_
	);
	LUT2 #(
		.INIT('h9)
	) name12289 (
		_w12065_,
		_w12322_,
		_w12323_
	);
	LUT4 #(
		.INIT('h6500)
	) name12290 (
		\a[11] ,
		_w12317_,
		_w12321_,
		_w12323_,
		_w12324_
	);
	LUT2 #(
		.INIT('h8)
	) name12291 (
		_w4684_,
		_w11434_,
		_w12325_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12292 (
		_w4700_,
		_w10991_,
		_w11230_,
		_w11232_,
		_w12326_
	);
	LUT4 #(
		.INIT('h000d)
	) name12293 (
		_w4459_,
		_w11581_,
		_w12325_,
		_w12326_,
		_w12327_
	);
	LUT2 #(
		.INIT('h4)
	) name12294 (
		_w4457_,
		_w11434_,
		_w12328_
	);
	LUT3 #(
		.INIT('h8a)
	) name12295 (
		\a[11] ,
		_w4457_,
		_w11434_,
		_w12329_
	);
	LUT2 #(
		.INIT('h8)
	) name12296 (
		_w12327_,
		_w12329_,
		_w12330_
	);
	LUT4 #(
		.INIT('h2882)
	) name12297 (
		_w4459_,
		_w11233_,
		_w11235_,
		_w11580_,
		_w12331_
	);
	LUT3 #(
		.INIT('h82)
	) name12298 (
		_w4700_,
		_w11233_,
		_w11235_,
		_w12332_
	);
	LUT2 #(
		.INIT('h8)
	) name12299 (
		_w4458_,
		_w11434_,
		_w12333_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12300 (
		_w4684_,
		_w10991_,
		_w11230_,
		_w11232_,
		_w12334_
	);
	LUT2 #(
		.INIT('h1)
	) name12301 (
		_w12333_,
		_w12334_,
		_w12335_
	);
	LUT3 #(
		.INIT('h10)
	) name12302 (
		_w12332_,
		_w12331_,
		_w12335_,
		_w12336_
	);
	LUT3 #(
		.INIT('h80)
	) name12303 (
		_w12066_,
		_w12330_,
		_w12336_,
		_w12337_
	);
	LUT3 #(
		.INIT('h28)
	) name12304 (
		_w4459_,
		_w11431_,
		_w11435_,
		_w12338_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12305 (
		_w4458_,
		_w10991_,
		_w11230_,
		_w11232_,
		_w12339_
	);
	LUT4 #(
		.INIT('h007d)
	) name12306 (
		_w4684_,
		_w11233_,
		_w11235_,
		_w12339_,
		_w12340_
	);
	LUT3 #(
		.INIT('h70)
	) name12307 (
		_w4700_,
		_w11427_,
		_w12340_,
		_w12341_
	);
	LUT3 #(
		.INIT('h9a)
	) name12308 (
		\a[11] ,
		_w12338_,
		_w12341_,
		_w12342_
	);
	LUT3 #(
		.INIT('h15)
	) name12309 (
		_w12066_,
		_w12330_,
		_w12336_,
		_w12343_
	);
	LUT3 #(
		.INIT('h6a)
	) name12310 (
		_w12066_,
		_w12330_,
		_w12336_,
		_w12344_
	);
	LUT3 #(
		.INIT('h54)
	) name12311 (
		_w12337_,
		_w12342_,
		_w12343_,
		_w12345_
	);
	LUT4 #(
		.INIT('h009a)
	) name12312 (
		\a[11] ,
		_w12317_,
		_w12321_,
		_w12323_,
		_w12346_
	);
	LUT4 #(
		.INIT('h9a65)
	) name12313 (
		\a[11] ,
		_w12317_,
		_w12321_,
		_w12323_,
		_w12347_
	);
	LUT3 #(
		.INIT('h54)
	) name12314 (
		_w12324_,
		_w12345_,
		_w12346_,
		_w12348_
	);
	LUT4 #(
		.INIT('h009a)
	) name12315 (
		\a[11] ,
		_w12308_,
		_w12313_,
		_w12315_,
		_w12349_
	);
	LUT4 #(
		.INIT('h9a65)
	) name12316 (
		\a[11] ,
		_w12308_,
		_w12313_,
		_w12315_,
		_w12350_
	);
	LUT3 #(
		.INIT('h54)
	) name12317 (
		_w12316_,
		_w12348_,
		_w12349_,
		_w12351_
	);
	LUT2 #(
		.INIT('h2)
	) name12318 (
		_w12305_,
		_w12306_,
		_w12352_
	);
	LUT2 #(
		.INIT('h9)
	) name12319 (
		_w12305_,
		_w12306_,
		_w12353_
	);
	LUT4 #(
		.INIT('h9a65)
	) name12320 (
		\a[11] ,
		_w12295_,
		_w12299_,
		_w12300_,
		_w12354_
	);
	LUT4 #(
		.INIT('h4d00)
	) name12321 (
		_w12305_,
		_w12306_,
		_w12351_,
		_w12354_,
		_w12355_
	);
	LUT4 #(
		.INIT('h9699)
	) name12322 (
		\a[11] ,
		_w12287_,
		_w12288_,
		_w12293_,
		_w12356_
	);
	LUT4 #(
		.INIT('h0155)
	) name12323 (
		_w12294_,
		_w12301_,
		_w12355_,
		_w12356_,
		_w12357_
	);
	LUT2 #(
		.INIT('h4)
	) name12324 (
		_w12281_,
		_w12285_,
		_w12358_
	);
	LUT2 #(
		.INIT('h9)
	) name12325 (
		_w12281_,
		_w12285_,
		_w12359_
	);
	LUT3 #(
		.INIT('h54)
	) name12326 (
		_w12286_,
		_w12357_,
		_w12358_,
		_w12360_
	);
	LUT3 #(
		.INIT('h12)
	) name12327 (
		\a[11] ,
		_w12275_,
		_w12279_,
		_w12361_
	);
	LUT3 #(
		.INIT('h69)
	) name12328 (
		\a[11] ,
		_w12275_,
		_w12279_,
		_w12362_
	);
	LUT3 #(
		.INIT('h54)
	) name12329 (
		_w12280_,
		_w12360_,
		_w12361_,
		_w12363_
	);
	LUT3 #(
		.INIT('h06)
	) name12330 (
		\a[11] ,
		_w12272_,
		_w12273_,
		_w12364_
	);
	LUT3 #(
		.INIT('h69)
	) name12331 (
		\a[11] ,
		_w12272_,
		_w12273_,
		_w12365_
	);
	LUT3 #(
		.INIT('h54)
	) name12332 (
		_w12274_,
		_w12363_,
		_w12364_,
		_w12366_
	);
	LUT3 #(
		.INIT('h06)
	) name12333 (
		\a[11] ,
		_w12266_,
		_w12267_,
		_w12367_
	);
	LUT3 #(
		.INIT('h69)
	) name12334 (
		\a[11] ,
		_w12266_,
		_w12267_,
		_w12368_
	);
	LUT3 #(
		.INIT('h54)
	) name12335 (
		_w12268_,
		_w12366_,
		_w12367_,
		_w12369_
	);
	LUT3 #(
		.INIT('h06)
	) name12336 (
		\a[11] ,
		_w12260_,
		_w12261_,
		_w12370_
	);
	LUT3 #(
		.INIT('h69)
	) name12337 (
		\a[11] ,
		_w12260_,
		_w12261_,
		_w12371_
	);
	LUT3 #(
		.INIT('h54)
	) name12338 (
		_w12262_,
		_w12369_,
		_w12370_,
		_w12372_
	);
	LUT2 #(
		.INIT('h4)
	) name12339 (
		_w12251_,
		_w12255_,
		_w12373_
	);
	LUT2 #(
		.INIT('h9)
	) name12340 (
		_w12251_,
		_w12255_,
		_w12374_
	);
	LUT4 #(
		.INIT('h9699)
	) name12341 (
		\a[11] ,
		_w12244_,
		_w12245_,
		_w12249_,
		_w12375_
	);
	LUT4 #(
		.INIT('h2b00)
	) name12342 (
		_w12251_,
		_w12255_,
		_w12372_,
		_w12375_,
		_w12376_
	);
	LUT4 #(
		.INIT('h9699)
	) name12343 (
		\a[11] ,
		_w12236_,
		_w12237_,
		_w12242_,
		_w12377_
	);
	LUT4 #(
		.INIT('h0155)
	) name12344 (
		_w12243_,
		_w12250_,
		_w12376_,
		_w12377_,
		_w12378_
	);
	LUT2 #(
		.INIT('h2)
	) name12345 (
		_w12233_,
		_w12234_,
		_w12379_
	);
	LUT2 #(
		.INIT('h9)
	) name12346 (
		_w12233_,
		_w12234_,
		_w12380_
	);
	LUT4 #(
		.INIT('h9a65)
	) name12347 (
		\a[11] ,
		_w12223_,
		_w12227_,
		_w12228_,
		_w12381_
	);
	LUT4 #(
		.INIT('h4d00)
	) name12348 (
		_w12233_,
		_w12234_,
		_w12378_,
		_w12381_,
		_w12382_
	);
	LUT4 #(
		.INIT('h9a65)
	) name12349 (
		\a[11] ,
		_w12215_,
		_w12220_,
		_w12221_,
		_w12383_
	);
	LUT4 #(
		.INIT('h0155)
	) name12350 (
		_w12222_,
		_w12229_,
		_w12382_,
		_w12383_,
		_w12384_
	);
	LUT2 #(
		.INIT('h4)
	) name12351 (
		_w12208_,
		_w12213_,
		_w12385_
	);
	LUT2 #(
		.INIT('h9)
	) name12352 (
		_w12208_,
		_w12213_,
		_w12386_
	);
	LUT4 #(
		.INIT('h9699)
	) name12353 (
		\a[11] ,
		_w12201_,
		_w12202_,
		_w12206_,
		_w12387_
	);
	LUT4 #(
		.INIT('h2b00)
	) name12354 (
		_w12208_,
		_w12213_,
		_w12384_,
		_w12387_,
		_w12388_
	);
	LUT4 #(
		.INIT('h9a65)
	) name12355 (
		\a[11] ,
		_w11558_,
		_w11563_,
		_w12199_,
		_w12389_
	);
	LUT4 #(
		.INIT('h0155)
	) name12356 (
		_w12200_,
		_w12207_,
		_w12388_,
		_w12389_,
		_w12390_
	);
	LUT4 #(
		.INIT('h54ab)
	) name12357 (
		_w11392_,
		_w11478_,
		_w11479_,
		_w11481_,
		_w12391_
	);
	LUT4 #(
		.INIT('h2228)
	) name12358 (
		_w4458_,
		_w8466_,
		_w8541_,
		_w11273_,
		_w12392_
	);
	LUT4 #(
		.INIT('h007d)
	) name12359 (
		_w4684_,
		_w11274_,
		_w11276_,
		_w12392_,
		_w12393_
	);
	LUT3 #(
		.INIT('h70)
	) name12360 (
		_w4700_,
		_w11388_,
		_w12393_,
		_w12394_
	);
	LUT4 #(
		.INIT('h95aa)
	) name12361 (
		\a[11] ,
		_w4459_,
		_w12391_,
		_w12394_,
		_w12395_
	);
	LUT4 #(
		.INIT('h010f)
	) name12362 (
		_w11966_,
		_w12120_,
		_w12197_,
		_w12198_,
		_w12396_
	);
	LUT4 #(
		.INIT('h010f)
	) name12363 (
		_w11962_,
		_w11964_,
		_w12188_,
		_w12189_,
		_w12397_
	);
	LUT4 #(
		.INIT('h2228)
	) name12364 (
		_w3709_,
		_w9446_,
		_w9702_,
		_w11261_,
		_w12398_
	);
	LUT4 #(
		.INIT('h007d)
	) name12365 (
		_w3877_,
		_w11262_,
		_w11264_,
		_w12398_,
		_w12399_
	);
	LUT3 #(
		.INIT('h70)
	) name12366 (
		_w3886_,
		_w11400_,
		_w12399_,
		_w12400_
	);
	LUT4 #(
		.INIT('h95aa)
	) name12367 (
		\a[17] ,
		_w3710_,
		_w11967_,
		_w12400_,
		_w12401_
	);
	LUT3 #(
		.INIT('h32)
	) name12368 (
		_w12127_,
		_w12184_,
		_w12185_,
		_w12402_
	);
	LUT3 #(
		.INIT('h32)
	) name12369 (
		_w12128_,
		_w12176_,
		_w12177_,
		_w12403_
	);
	LUT2 #(
		.INIT('h8)
	) name12370 (
		_w3214_,
		_w11415_,
		_w12404_
	);
	LUT4 #(
		.INIT('h007d)
	) name12371 (
		_w3249_,
		_w10599_,
		_w11253_,
		_w12404_,
		_w12405_
	);
	LUT4 #(
		.INIT('h7d00)
	) name12372 (
		_w3262_,
		_w10580_,
		_w11254_,
		_w12405_,
		_w12406_
	);
	LUT4 #(
		.INIT('h7d00)
	) name12373 (
		_w37_,
		_w11453_,
		_w11455_,
		_w12406_,
		_w12407_
	);
	LUT3 #(
		.INIT('h32)
	) name12374 (
		_w12138_,
		_w12168_,
		_w12169_,
		_w12408_
	);
	LUT3 #(
		.INIT('h82)
	) name12375 (
		_w2550_,
		_w11439_,
		_w11441_,
		_w12409_
	);
	LUT3 #(
		.INIT('h82)
	) name12376 (
		_w2854_,
		_w11241_,
		_w11243_,
		_w12410_
	);
	LUT2 #(
		.INIT('h8)
	) name12377 (
		_w2549_,
		_w11427_,
		_w12411_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12378 (
		_w2617_,
		_w10968_,
		_w11238_,
		_w11240_,
		_w12412_
	);
	LUT2 #(
		.INIT('h1)
	) name12379 (
		_w12411_,
		_w12412_,
		_w12413_
	);
	LUT2 #(
		.INIT('h4)
	) name12380 (
		_w12410_,
		_w12413_,
		_w12414_
	);
	LUT3 #(
		.INIT('h80)
	) name12381 (
		_w2039_,
		_w3144_,
		_w7297_,
		_w12415_
	);
	LUT4 #(
		.INIT('h8000)
	) name12382 (
		_w1277_,
		_w2688_,
		_w2896_,
		_w12415_,
		_w12416_
	);
	LUT4 #(
		.INIT('h8000)
	) name12383 (
		_w518_,
		_w964_,
		_w1360_,
		_w1438_,
		_w12417_
	);
	LUT4 #(
		.INIT('h153f)
	) name12384 (
		_w90_,
		_w41_,
		_w72_,
		_w39_,
		_w12418_
	);
	LUT2 #(
		.INIT('h4)
	) name12385 (
		_w186_,
		_w12418_,
		_w12419_
	);
	LUT4 #(
		.INIT('h153f)
	) name12386 (
		_w110_,
		_w78_,
		_w90_,
		_w158_,
		_w12420_
	);
	LUT4 #(
		.INIT('h2000)
	) name12387 (
		_w42_,
		_w186_,
		_w12418_,
		_w12420_,
		_w12421_
	);
	LUT4 #(
		.INIT('h8000)
	) name12388 (
		_w2670_,
		_w3546_,
		_w12417_,
		_w12421_,
		_w12422_
	);
	LUT4 #(
		.INIT('h8000)
	) name12389 (
		_w4199_,
		_w4206_,
		_w12416_,
		_w12422_,
		_w12423_
	);
	LUT2 #(
		.INIT('h8)
	) name12390 (
		_w8268_,
		_w12423_,
		_w12424_
	);
	LUT3 #(
		.INIT('h01)
	) name12391 (
		_w12163_,
		_w12166_,
		_w12424_,
		_w12425_
	);
	LUT3 #(
		.INIT('he0)
	) name12392 (
		_w12163_,
		_w12166_,
		_w12424_,
		_w12426_
	);
	LUT3 #(
		.INIT('h1e)
	) name12393 (
		_w12163_,
		_w12166_,
		_w12424_,
		_w12427_
	);
	LUT4 #(
		.INIT('h2882)
	) name12394 (
		_w377_,
		_w11233_,
		_w11235_,
		_w11580_,
		_w12428_
	);
	LUT3 #(
		.INIT('h82)
	) name12395 (
		_w2527_,
		_w11233_,
		_w11235_,
		_w12429_
	);
	LUT2 #(
		.INIT('h8)
	) name12396 (
		_w376_,
		_w11434_,
		_w12430_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12397 (
		_w2407_,
		_w10991_,
		_w11230_,
		_w11232_,
		_w12431_
	);
	LUT2 #(
		.INIT('h1)
	) name12398 (
		_w12430_,
		_w12431_,
		_w12432_
	);
	LUT3 #(
		.INIT('h10)
	) name12399 (
		_w12429_,
		_w12428_,
		_w12432_,
		_w12433_
	);
	LUT2 #(
		.INIT('h9)
	) name12400 (
		_w12427_,
		_w12433_,
		_w12434_
	);
	LUT4 #(
		.INIT('h6500)
	) name12401 (
		\a[29] ,
		_w12409_,
		_w12414_,
		_w12434_,
		_w12435_
	);
	LUT4 #(
		.INIT('h009a)
	) name12402 (
		\a[29] ,
		_w12409_,
		_w12414_,
		_w12434_,
		_w12436_
	);
	LUT4 #(
		.INIT('h9a65)
	) name12403 (
		\a[29] ,
		_w12409_,
		_w12414_,
		_w12434_,
		_w12437_
	);
	LUT2 #(
		.INIT('h9)
	) name12404 (
		_w12408_,
		_w12437_,
		_w12438_
	);
	LUT3 #(
		.INIT('h82)
	) name12405 (
		_w2875_,
		_w11445_,
		_w11447_,
		_w12439_
	);
	LUT3 #(
		.INIT('h82)
	) name12406 (
		_w2986_,
		_w11249_,
		_w11251_,
		_w12440_
	);
	LUT2 #(
		.INIT('h8)
	) name12407 (
		_w2874_,
		_w11421_,
		_w12441_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12408 (
		_w2975_,
		_w10945_,
		_w11246_,
		_w11248_,
		_w12442_
	);
	LUT2 #(
		.INIT('h1)
	) name12409 (
		_w12441_,
		_w12442_,
		_w12443_
	);
	LUT2 #(
		.INIT('h4)
	) name12410 (
		_w12440_,
		_w12443_,
		_w12444_
	);
	LUT4 #(
		.INIT('h4844)
	) name12411 (
		\a[26] ,
		_w12438_,
		_w12439_,
		_w12444_,
		_w12445_
	);
	LUT4 #(
		.INIT('h9699)
	) name12412 (
		\a[26] ,
		_w12438_,
		_w12439_,
		_w12444_,
		_w12446_
	);
	LUT3 #(
		.INIT('h1e)
	) name12413 (
		_w12172_,
		_w12174_,
		_w12446_,
		_w12447_
	);
	LUT3 #(
		.INIT('h90)
	) name12414 (
		\a[23] ,
		_w12407_,
		_w12447_,
		_w12448_
	);
	LUT3 #(
		.INIT('h06)
	) name12415 (
		\a[23] ,
		_w12407_,
		_w12447_,
		_w12449_
	);
	LUT3 #(
		.INIT('h69)
	) name12416 (
		\a[23] ,
		_w12407_,
		_w12447_,
		_w12450_
	);
	LUT2 #(
		.INIT('h9)
	) name12417 (
		_w12403_,
		_w12450_,
		_w12451_
	);
	LUT3 #(
		.INIT('h82)
	) name12418 (
		_w3311_,
		_w10268_,
		_w11255_,
		_w12452_
	);
	LUT4 #(
		.INIT('h007d)
	) name12419 (
		_w3645_,
		_w11256_,
		_w11258_,
		_w12452_,
		_w12453_
	);
	LUT3 #(
		.INIT('h70)
	) name12420 (
		_w3654_,
		_w11406_,
		_w12453_,
		_w12454_
	);
	LUT4 #(
		.INIT('h95aa)
	) name12421 (
		\a[20] ,
		_w3312_,
		_w11796_,
		_w12454_,
		_w12455_
	);
	LUT2 #(
		.INIT('h2)
	) name12422 (
		_w12451_,
		_w12455_,
		_w12456_
	);
	LUT2 #(
		.INIT('h4)
	) name12423 (
		_w12451_,
		_w12455_,
		_w12457_
	);
	LUT2 #(
		.INIT('h9)
	) name12424 (
		_w12451_,
		_w12455_,
		_w12458_
	);
	LUT2 #(
		.INIT('h9)
	) name12425 (
		_w12402_,
		_w12458_,
		_w12459_
	);
	LUT2 #(
		.INIT('h4)
	) name12426 (
		_w12401_,
		_w12459_,
		_w12460_
	);
	LUT2 #(
		.INIT('h2)
	) name12427 (
		_w12401_,
		_w12459_,
		_w12461_
	);
	LUT2 #(
		.INIT('h9)
	) name12428 (
		_w12401_,
		_w12459_,
		_w12462_
	);
	LUT2 #(
		.INIT('h9)
	) name12429 (
		_w12397_,
		_w12462_,
		_w12463_
	);
	LUT4 #(
		.INIT('h2228)
	) name12430 (
		_w4033_,
		_w8794_,
		_w8994_,
		_w11267_,
		_w12464_
	);
	LUT4 #(
		.INIT('h007d)
	) name12431 (
		_w4367_,
		_w11268_,
		_w11270_,
		_w12464_,
		_w12465_
	);
	LUT3 #(
		.INIT('h70)
	) name12432 (
		_w4382_,
		_w11394_,
		_w12465_,
		_w12466_
	);
	LUT4 #(
		.INIT('h95aa)
	) name12433 (
		\a[14] ,
		_w4034_,
		_w12209_,
		_w12466_,
		_w12467_
	);
	LUT2 #(
		.INIT('h2)
	) name12434 (
		_w12463_,
		_w12467_,
		_w12468_
	);
	LUT2 #(
		.INIT('h4)
	) name12435 (
		_w12463_,
		_w12467_,
		_w12469_
	);
	LUT2 #(
		.INIT('h9)
	) name12436 (
		_w12463_,
		_w12467_,
		_w12470_
	);
	LUT2 #(
		.INIT('h9)
	) name12437 (
		_w12396_,
		_w12470_,
		_w12471_
	);
	LUT2 #(
		.INIT('h4)
	) name12438 (
		_w12395_,
		_w12471_,
		_w12472_
	);
	LUT2 #(
		.INIT('h2)
	) name12439 (
		_w12395_,
		_w12471_,
		_w12473_
	);
	LUT2 #(
		.INIT('h9)
	) name12440 (
		_w12395_,
		_w12471_,
		_w12474_
	);
	LUT2 #(
		.INIT('h9)
	) name12441 (
		_w12390_,
		_w12474_,
		_w12475_
	);
	LUT4 #(
		.INIT('h54ab)
	) name12442 (
		_w11386_,
		_w11484_,
		_w11485_,
		_w11487_,
		_w12476_
	);
	LUT4 #(
		.INIT('h2228)
	) name12443 (
		_w4875_,
		_w7935_,
		_w8077_,
		_w11279_,
		_w12477_
	);
	LUT4 #(
		.INIT('h007d)
	) name12444 (
		_w5271_,
		_w11280_,
		_w11282_,
		_w12477_,
		_w12478_
	);
	LUT3 #(
		.INIT('h70)
	) name12445 (
		_w5286_,
		_w11382_,
		_w12478_,
		_w12479_
	);
	LUT4 #(
		.INIT('h95aa)
	) name12446 (
		\a[8] ,
		_w4876_,
		_w12476_,
		_w12479_,
		_w12480_
	);
	LUT2 #(
		.INIT('h2)
	) name12447 (
		_w12475_,
		_w12480_,
		_w12481_
	);
	LUT3 #(
		.INIT('h1e)
	) name12448 (
		_w12207_,
		_w12388_,
		_w12389_,
		_w12482_
	);
	LUT3 #(
		.INIT('h82)
	) name12449 (
		_w4876_,
		_w11484_,
		_w11486_,
		_w12483_
	);
	LUT3 #(
		.INIT('h82)
	) name12450 (
		_w5286_,
		_w11280_,
		_w11282_,
		_w12484_
	);
	LUT2 #(
		.INIT('h8)
	) name12451 (
		_w4875_,
		_w11388_,
		_w12485_
	);
	LUT4 #(
		.INIT('h2228)
	) name12452 (
		_w5271_,
		_w7935_,
		_w8077_,
		_w11279_,
		_w12486_
	);
	LUT2 #(
		.INIT('h1)
	) name12453 (
		_w12485_,
		_w12486_,
		_w12487_
	);
	LUT2 #(
		.INIT('h4)
	) name12454 (
		_w12484_,
		_w12487_,
		_w12488_
	);
	LUT4 #(
		.INIT('h4844)
	) name12455 (
		\a[8] ,
		_w12482_,
		_w12483_,
		_w12488_,
		_w12489_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12456 (
		_w4876_,
		_w11390_,
		_w11482_,
		_w11483_,
		_w12490_
	);
	LUT4 #(
		.INIT('h2228)
	) name12457 (
		_w5286_,
		_w7935_,
		_w8077_,
		_w11279_,
		_w12491_
	);
	LUT3 #(
		.INIT('h82)
	) name12458 (
		_w4875_,
		_w11274_,
		_w11276_,
		_w12492_
	);
	LUT3 #(
		.INIT('h07)
	) name12459 (
		_w5271_,
		_w11388_,
		_w12492_,
		_w12493_
	);
	LUT2 #(
		.INIT('h4)
	) name12460 (
		_w12491_,
		_w12493_,
		_w12494_
	);
	LUT4 #(
		.INIT('h54ab)
	) name12461 (
		_w12214_,
		_w12384_,
		_w12385_,
		_w12387_,
		_w12495_
	);
	LUT4 #(
		.INIT('h6500)
	) name12462 (
		\a[8] ,
		_w12490_,
		_w12494_,
		_w12495_,
		_w12496_
	);
	LUT4 #(
		.INIT('h2228)
	) name12463 (
		_w4875_,
		_w8466_,
		_w8541_,
		_w11273_,
		_w12497_
	);
	LUT4 #(
		.INIT('h007d)
	) name12464 (
		_w5271_,
		_w11274_,
		_w11276_,
		_w12497_,
		_w12498_
	);
	LUT3 #(
		.INIT('h70)
	) name12465 (
		_w5286_,
		_w11388_,
		_w12498_,
		_w12499_
	);
	LUT4 #(
		.INIT('h95aa)
	) name12466 (
		\a[8] ,
		_w4876_,
		_w12391_,
		_w12499_,
		_w12500_
	);
	LUT2 #(
		.INIT('h9)
	) name12467 (
		_w12384_,
		_w12386_,
		_w12501_
	);
	LUT2 #(
		.INIT('h4)
	) name12468 (
		_w12500_,
		_w12501_,
		_w12502_
	);
	LUT3 #(
		.INIT('h1e)
	) name12469 (
		_w12229_,
		_w12382_,
		_w12383_,
		_w12503_
	);
	LUT3 #(
		.INIT('h82)
	) name12470 (
		_w4876_,
		_w11478_,
		_w11480_,
		_w12504_
	);
	LUT3 #(
		.INIT('h82)
	) name12471 (
		_w5286_,
		_w11274_,
		_w11276_,
		_w12505_
	);
	LUT2 #(
		.INIT('h8)
	) name12472 (
		_w4875_,
		_w11394_,
		_w12506_
	);
	LUT4 #(
		.INIT('h2228)
	) name12473 (
		_w5271_,
		_w8466_,
		_w8541_,
		_w11273_,
		_w12507_
	);
	LUT2 #(
		.INIT('h1)
	) name12474 (
		_w12506_,
		_w12507_,
		_w12508_
	);
	LUT2 #(
		.INIT('h4)
	) name12475 (
		_w12505_,
		_w12508_,
		_w12509_
	);
	LUT4 #(
		.INIT('h4844)
	) name12476 (
		\a[8] ,
		_w12503_,
		_w12504_,
		_w12509_,
		_w12510_
	);
	LUT4 #(
		.INIT('h54ab)
	) name12477 (
		_w12235_,
		_w12378_,
		_w12379_,
		_w12381_,
		_w12511_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12478 (
		_w4876_,
		_w11396_,
		_w11476_,
		_w11477_,
		_w12512_
	);
	LUT4 #(
		.INIT('h2228)
	) name12479 (
		_w5286_,
		_w8466_,
		_w8541_,
		_w11273_,
		_w12513_
	);
	LUT3 #(
		.INIT('h82)
	) name12480 (
		_w4875_,
		_w11268_,
		_w11270_,
		_w12514_
	);
	LUT3 #(
		.INIT('h07)
	) name12481 (
		_w5271_,
		_w11394_,
		_w12514_,
		_w12515_
	);
	LUT2 #(
		.INIT('h4)
	) name12482 (
		_w12513_,
		_w12515_,
		_w12516_
	);
	LUT4 #(
		.INIT('h4844)
	) name12483 (
		\a[8] ,
		_w12511_,
		_w12512_,
		_w12516_,
		_w12517_
	);
	LUT2 #(
		.INIT('h9)
	) name12484 (
		_w12378_,
		_w12380_,
		_w12518_
	);
	LUT4 #(
		.INIT('h2228)
	) name12485 (
		_w4875_,
		_w8794_,
		_w8994_,
		_w11267_,
		_w12519_
	);
	LUT4 #(
		.INIT('h007d)
	) name12486 (
		_w5271_,
		_w11268_,
		_w11270_,
		_w12519_,
		_w12520_
	);
	LUT3 #(
		.INIT('h70)
	) name12487 (
		_w5286_,
		_w11394_,
		_w12520_,
		_w12521_
	);
	LUT4 #(
		.INIT('h95aa)
	) name12488 (
		\a[8] ,
		_w4876_,
		_w12209_,
		_w12521_,
		_w12522_
	);
	LUT2 #(
		.INIT('h2)
	) name12489 (
		_w12518_,
		_w12522_,
		_w12523_
	);
	LUT3 #(
		.INIT('h82)
	) name12490 (
		_w4876_,
		_w11472_,
		_w11474_,
		_w12524_
	);
	LUT3 #(
		.INIT('h82)
	) name12491 (
		_w5286_,
		_w11268_,
		_w11270_,
		_w12525_
	);
	LUT2 #(
		.INIT('h8)
	) name12492 (
		_w4875_,
		_w11400_,
		_w12526_
	);
	LUT4 #(
		.INIT('h2228)
	) name12493 (
		_w5271_,
		_w8794_,
		_w8994_,
		_w11267_,
		_w12527_
	);
	LUT2 #(
		.INIT('h1)
	) name12494 (
		_w12526_,
		_w12527_,
		_w12528_
	);
	LUT2 #(
		.INIT('h4)
	) name12495 (
		_w12525_,
		_w12528_,
		_w12529_
	);
	LUT3 #(
		.INIT('h1e)
	) name12496 (
		_w12250_,
		_w12376_,
		_w12377_,
		_w12530_
	);
	LUT4 #(
		.INIT('h6500)
	) name12497 (
		\a[8] ,
		_w12524_,
		_w12529_,
		_w12530_,
		_w12531_
	);
	LUT3 #(
		.INIT('h82)
	) name12498 (
		_w4876_,
		_w11469_,
		_w11471_,
		_w12532_
	);
	LUT4 #(
		.INIT('h2228)
	) name12499 (
		_w5286_,
		_w8794_,
		_w8994_,
		_w11267_,
		_w12533_
	);
	LUT3 #(
		.INIT('h82)
	) name12500 (
		_w4875_,
		_w11262_,
		_w11264_,
		_w12534_
	);
	LUT3 #(
		.INIT('h07)
	) name12501 (
		_w5271_,
		_w11400_,
		_w12534_,
		_w12535_
	);
	LUT2 #(
		.INIT('h4)
	) name12502 (
		_w12533_,
		_w12535_,
		_w12536_
	);
	LUT4 #(
		.INIT('h54ab)
	) name12503 (
		_w12256_,
		_w12372_,
		_w12373_,
		_w12375_,
		_w12537_
	);
	LUT4 #(
		.INIT('h6500)
	) name12504 (
		\a[8] ,
		_w12532_,
		_w12536_,
		_w12537_,
		_w12538_
	);
	LUT4 #(
		.INIT('h2228)
	) name12505 (
		_w4875_,
		_w9446_,
		_w9702_,
		_w11261_,
		_w12539_
	);
	LUT4 #(
		.INIT('h007d)
	) name12506 (
		_w5271_,
		_w11262_,
		_w11264_,
		_w12539_,
		_w12540_
	);
	LUT3 #(
		.INIT('h70)
	) name12507 (
		_w5286_,
		_w11400_,
		_w12540_,
		_w12541_
	);
	LUT4 #(
		.INIT('h95aa)
	) name12508 (
		\a[8] ,
		_w4876_,
		_w11967_,
		_w12541_,
		_w12542_
	);
	LUT2 #(
		.INIT('h9)
	) name12509 (
		_w12372_,
		_w12374_,
		_w12543_
	);
	LUT2 #(
		.INIT('h4)
	) name12510 (
		_w12542_,
		_w12543_,
		_w12544_
	);
	LUT2 #(
		.INIT('h9)
	) name12511 (
		_w12369_,
		_w12371_,
		_w12545_
	);
	LUT3 #(
		.INIT('h82)
	) name12512 (
		_w4876_,
		_w11465_,
		_w11467_,
		_w12546_
	);
	LUT3 #(
		.INIT('h82)
	) name12513 (
		_w5286_,
		_w11262_,
		_w11264_,
		_w12547_
	);
	LUT2 #(
		.INIT('h8)
	) name12514 (
		_w4875_,
		_w11406_,
		_w12548_
	);
	LUT4 #(
		.INIT('h2228)
	) name12515 (
		_w5271_,
		_w9446_,
		_w9702_,
		_w11261_,
		_w12549_
	);
	LUT2 #(
		.INIT('h1)
	) name12516 (
		_w12548_,
		_w12549_,
		_w12550_
	);
	LUT2 #(
		.INIT('h4)
	) name12517 (
		_w12547_,
		_w12550_,
		_w12551_
	);
	LUT4 #(
		.INIT('h4844)
	) name12518 (
		\a[8] ,
		_w12545_,
		_w12546_,
		_w12551_,
		_w12552_
	);
	LUT2 #(
		.INIT('h9)
	) name12519 (
		_w12366_,
		_w12368_,
		_w12553_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12520 (
		_w4876_,
		_w11408_,
		_w11463_,
		_w11464_,
		_w12554_
	);
	LUT4 #(
		.INIT('h2228)
	) name12521 (
		_w5286_,
		_w9446_,
		_w9702_,
		_w11261_,
		_w12555_
	);
	LUT3 #(
		.INIT('h82)
	) name12522 (
		_w4875_,
		_w11256_,
		_w11258_,
		_w12556_
	);
	LUT3 #(
		.INIT('h07)
	) name12523 (
		_w5271_,
		_w11406_,
		_w12556_,
		_w12557_
	);
	LUT2 #(
		.INIT('h4)
	) name12524 (
		_w12555_,
		_w12557_,
		_w12558_
	);
	LUT4 #(
		.INIT('h4844)
	) name12525 (
		\a[8] ,
		_w12553_,
		_w12554_,
		_w12558_,
		_w12559_
	);
	LUT2 #(
		.INIT('h9)
	) name12526 (
		_w12363_,
		_w12365_,
		_w12560_
	);
	LUT3 #(
		.INIT('h82)
	) name12527 (
		_w4875_,
		_w10268_,
		_w11255_,
		_w12561_
	);
	LUT4 #(
		.INIT('h007d)
	) name12528 (
		_w5271_,
		_w11256_,
		_w11258_,
		_w12561_,
		_w12562_
	);
	LUT3 #(
		.INIT('h70)
	) name12529 (
		_w5286_,
		_w11406_,
		_w12562_,
		_w12563_
	);
	LUT4 #(
		.INIT('h95aa)
	) name12530 (
		\a[8] ,
		_w4876_,
		_w11796_,
		_w12563_,
		_w12564_
	);
	LUT2 #(
		.INIT('h2)
	) name12531 (
		_w12560_,
		_w12564_,
		_w12565_
	);
	LUT3 #(
		.INIT('h82)
	) name12532 (
		_w4875_,
		_w10580_,
		_w11254_,
		_w12566_
	);
	LUT4 #(
		.INIT('h007d)
	) name12533 (
		_w5271_,
		_w10268_,
		_w11255_,
		_w12566_,
		_w12567_
	);
	LUT4 #(
		.INIT('h7d00)
	) name12534 (
		_w5286_,
		_w11256_,
		_w11258_,
		_w12567_,
		_w12568_
	);
	LUT4 #(
		.INIT('h7d00)
	) name12535 (
		_w4876_,
		_w11459_,
		_w11461_,
		_w12568_,
		_w12569_
	);
	LUT2 #(
		.INIT('h9)
	) name12536 (
		_w12360_,
		_w12362_,
		_w12570_
	);
	LUT3 #(
		.INIT('h90)
	) name12537 (
		\a[8] ,
		_w12569_,
		_w12570_,
		_w12571_
	);
	LUT3 #(
		.INIT('h82)
	) name12538 (
		_w4875_,
		_w10599_,
		_w11253_,
		_w12572_
	);
	LUT4 #(
		.INIT('h007d)
	) name12539 (
		_w5271_,
		_w10580_,
		_w11254_,
		_w12572_,
		_w12573_
	);
	LUT4 #(
		.INIT('h7d00)
	) name12540 (
		_w5286_,
		_w10268_,
		_w11255_,
		_w12573_,
		_w12574_
	);
	LUT4 #(
		.INIT('h7d00)
	) name12541 (
		_w4876_,
		_w11456_,
		_w11458_,
		_w12574_,
		_w12575_
	);
	LUT2 #(
		.INIT('h9)
	) name12542 (
		_w12357_,
		_w12359_,
		_w12576_
	);
	LUT3 #(
		.INIT('h90)
	) name12543 (
		\a[8] ,
		_w12575_,
		_w12576_,
		_w12577_
	);
	LUT2 #(
		.INIT('h8)
	) name12544 (
		_w4875_,
		_w11415_,
		_w12578_
	);
	LUT4 #(
		.INIT('h007d)
	) name12545 (
		_w5271_,
		_w10599_,
		_w11253_,
		_w12578_,
		_w12579_
	);
	LUT4 #(
		.INIT('h7d00)
	) name12546 (
		_w5286_,
		_w10580_,
		_w11254_,
		_w12579_,
		_w12580_
	);
	LUT4 #(
		.INIT('h7d00)
	) name12547 (
		_w4876_,
		_w11453_,
		_w11455_,
		_w12580_,
		_w12581_
	);
	LUT3 #(
		.INIT('h1e)
	) name12548 (
		_w12301_,
		_w12355_,
		_w12356_,
		_w12582_
	);
	LUT3 #(
		.INIT('h90)
	) name12549 (
		\a[8] ,
		_w12581_,
		_w12582_,
		_w12583_
	);
	LUT4 #(
		.INIT('h54ab)
	) name12550 (
		_w12307_,
		_w12351_,
		_w12352_,
		_w12354_,
		_w12584_
	);
	LUT3 #(
		.INIT('h82)
	) name12551 (
		_w4875_,
		_w11249_,
		_w11251_,
		_w12585_
	);
	LUT3 #(
		.INIT('h07)
	) name12552 (
		_w5271_,
		_w11415_,
		_w12585_,
		_w12586_
	);
	LUT4 #(
		.INIT('h7d00)
	) name12553 (
		_w5286_,
		_w10599_,
		_w11253_,
		_w12586_,
		_w12587_
	);
	LUT4 #(
		.INIT('h7d00)
	) name12554 (
		_w4876_,
		_w11450_,
		_w11452_,
		_w12587_,
		_w12588_
	);
	LUT3 #(
		.INIT('h84)
	) name12555 (
		\a[8] ,
		_w12584_,
		_w12588_,
		_w12589_
	);
	LUT2 #(
		.INIT('h9)
	) name12556 (
		_w12351_,
		_w12353_,
		_w12590_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12557 (
		_w4875_,
		_w10945_,
		_w11246_,
		_w11248_,
		_w12591_
	);
	LUT4 #(
		.INIT('h007d)
	) name12558 (
		_w5271_,
		_w11249_,
		_w11251_,
		_w12591_,
		_w12592_
	);
	LUT3 #(
		.INIT('h70)
	) name12559 (
		_w5286_,
		_w11415_,
		_w12592_,
		_w12593_
	);
	LUT4 #(
		.INIT('h95aa)
	) name12560 (
		\a[8] ,
		_w4876_,
		_w11675_,
		_w12593_,
		_w12594_
	);
	LUT2 #(
		.INIT('h2)
	) name12561 (
		_w12590_,
		_w12594_,
		_w12595_
	);
	LUT2 #(
		.INIT('h9)
	) name12562 (
		_w12348_,
		_w12350_,
		_w12596_
	);
	LUT3 #(
		.INIT('h82)
	) name12563 (
		_w4876_,
		_w11445_,
		_w11447_,
		_w12597_
	);
	LUT3 #(
		.INIT('h82)
	) name12564 (
		_w5286_,
		_w11249_,
		_w11251_,
		_w12598_
	);
	LUT2 #(
		.INIT('h8)
	) name12565 (
		_w4875_,
		_w11421_,
		_w12599_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12566 (
		_w5271_,
		_w10945_,
		_w11246_,
		_w11248_,
		_w12600_
	);
	LUT2 #(
		.INIT('h1)
	) name12567 (
		_w12599_,
		_w12600_,
		_w12601_
	);
	LUT2 #(
		.INIT('h4)
	) name12568 (
		_w12598_,
		_w12601_,
		_w12602_
	);
	LUT4 #(
		.INIT('h4844)
	) name12569 (
		\a[8] ,
		_w12596_,
		_w12597_,
		_w12602_,
		_w12603_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12570 (
		_w4876_,
		_w11423_,
		_w11443_,
		_w11444_,
		_w12604_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12571 (
		_w5286_,
		_w10945_,
		_w11246_,
		_w11248_,
		_w12605_
	);
	LUT3 #(
		.INIT('h82)
	) name12572 (
		_w4875_,
		_w11241_,
		_w11243_,
		_w12606_
	);
	LUT3 #(
		.INIT('h07)
	) name12573 (
		_w5271_,
		_w11421_,
		_w12606_,
		_w12607_
	);
	LUT2 #(
		.INIT('h4)
	) name12574 (
		_w12605_,
		_w12607_,
		_w12608_
	);
	LUT2 #(
		.INIT('h9)
	) name12575 (
		_w12345_,
		_w12347_,
		_w12609_
	);
	LUT4 #(
		.INIT('h6500)
	) name12576 (
		\a[8] ,
		_w12604_,
		_w12608_,
		_w12609_,
		_w12610_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12577 (
		_w4875_,
		_w10968_,
		_w11238_,
		_w11240_,
		_w12611_
	);
	LUT4 #(
		.INIT('h007d)
	) name12578 (
		_w5271_,
		_w11241_,
		_w11243_,
		_w12611_,
		_w12612_
	);
	LUT3 #(
		.INIT('h70)
	) name12579 (
		_w5286_,
		_w11421_,
		_w12612_,
		_w12613_
	);
	LUT4 #(
		.INIT('h95aa)
	) name12580 (
		\a[8] ,
		_w4876_,
		_w11569_,
		_w12613_,
		_w12614_
	);
	LUT2 #(
		.INIT('h9)
	) name12581 (
		_w12342_,
		_w12344_,
		_w12615_
	);
	LUT2 #(
		.INIT('h4)
	) name12582 (
		_w12614_,
		_w12615_,
		_w12616_
	);
	LUT3 #(
		.INIT('h82)
	) name12583 (
		_w4876_,
		_w11439_,
		_w11441_,
		_w12617_
	);
	LUT3 #(
		.INIT('h82)
	) name12584 (
		_w5286_,
		_w11241_,
		_w11243_,
		_w12618_
	);
	LUT2 #(
		.INIT('h8)
	) name12585 (
		_w4875_,
		_w11427_,
		_w12619_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12586 (
		_w5271_,
		_w10968_,
		_w11238_,
		_w11240_,
		_w12620_
	);
	LUT2 #(
		.INIT('h1)
	) name12587 (
		_w12619_,
		_w12620_,
		_w12621_
	);
	LUT2 #(
		.INIT('h4)
	) name12588 (
		_w12618_,
		_w12621_,
		_w12622_
	);
	LUT3 #(
		.INIT('h8a)
	) name12589 (
		\a[11] ,
		_w12328_,
		_w12327_,
		_w12623_
	);
	LUT2 #(
		.INIT('h9)
	) name12590 (
		_w12336_,
		_w12623_,
		_w12624_
	);
	LUT4 #(
		.INIT('h6500)
	) name12591 (
		\a[8] ,
		_w12617_,
		_w12622_,
		_w12624_,
		_w12625_
	);
	LUT3 #(
		.INIT('h82)
	) name12592 (
		_w4876_,
		_w11436_,
		_w11438_,
		_w12626_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12593 (
		_w5286_,
		_w10968_,
		_w11238_,
		_w11240_,
		_w12627_
	);
	LUT3 #(
		.INIT('h82)
	) name12594 (
		_w4875_,
		_w11233_,
		_w11235_,
		_w12628_
	);
	LUT3 #(
		.INIT('h07)
	) name12595 (
		_w5271_,
		_w11427_,
		_w12628_,
		_w12629_
	);
	LUT2 #(
		.INIT('h4)
	) name12596 (
		_w12627_,
		_w12629_,
		_w12630_
	);
	LUT3 #(
		.INIT('h20)
	) name12597 (
		\a[11] ,
		_w4457_,
		_w11434_,
		_w12631_
	);
	LUT2 #(
		.INIT('h9)
	) name12598 (
		_w12327_,
		_w12631_,
		_w12632_
	);
	LUT4 #(
		.INIT('h6500)
	) name12599 (
		\a[8] ,
		_w12626_,
		_w12630_,
		_w12632_,
		_w12633_
	);
	LUT2 #(
		.INIT('h8)
	) name12600 (
		_w5271_,
		_w11434_,
		_w12634_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12601 (
		_w5286_,
		_w10991_,
		_w11230_,
		_w11232_,
		_w12635_
	);
	LUT4 #(
		.INIT('h000d)
	) name12602 (
		_w4876_,
		_w11581_,
		_w12634_,
		_w12635_,
		_w12636_
	);
	LUT2 #(
		.INIT('h4)
	) name12603 (
		_w4874_,
		_w11434_,
		_w12637_
	);
	LUT3 #(
		.INIT('h8a)
	) name12604 (
		\a[8] ,
		_w4874_,
		_w11434_,
		_w12638_
	);
	LUT2 #(
		.INIT('h8)
	) name12605 (
		_w12636_,
		_w12638_,
		_w12639_
	);
	LUT4 #(
		.INIT('h2882)
	) name12606 (
		_w4876_,
		_w11233_,
		_w11235_,
		_w11580_,
		_w12640_
	);
	LUT3 #(
		.INIT('h82)
	) name12607 (
		_w5286_,
		_w11233_,
		_w11235_,
		_w12641_
	);
	LUT2 #(
		.INIT('h8)
	) name12608 (
		_w4875_,
		_w11434_,
		_w12642_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12609 (
		_w5271_,
		_w10991_,
		_w11230_,
		_w11232_,
		_w12643_
	);
	LUT2 #(
		.INIT('h1)
	) name12610 (
		_w12642_,
		_w12643_,
		_w12644_
	);
	LUT3 #(
		.INIT('h10)
	) name12611 (
		_w12641_,
		_w12640_,
		_w12644_,
		_w12645_
	);
	LUT3 #(
		.INIT('h80)
	) name12612 (
		_w12328_,
		_w12639_,
		_w12645_,
		_w12646_
	);
	LUT3 #(
		.INIT('h28)
	) name12613 (
		_w4876_,
		_w11431_,
		_w11435_,
		_w12647_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12614 (
		_w4875_,
		_w10991_,
		_w11230_,
		_w11232_,
		_w12648_
	);
	LUT4 #(
		.INIT('h007d)
	) name12615 (
		_w5271_,
		_w11233_,
		_w11235_,
		_w12648_,
		_w12649_
	);
	LUT3 #(
		.INIT('h70)
	) name12616 (
		_w5286_,
		_w11427_,
		_w12649_,
		_w12650_
	);
	LUT3 #(
		.INIT('h9a)
	) name12617 (
		\a[8] ,
		_w12647_,
		_w12650_,
		_w12651_
	);
	LUT3 #(
		.INIT('h15)
	) name12618 (
		_w12328_,
		_w12639_,
		_w12645_,
		_w12652_
	);
	LUT3 #(
		.INIT('h6a)
	) name12619 (
		_w12328_,
		_w12639_,
		_w12645_,
		_w12653_
	);
	LUT3 #(
		.INIT('h54)
	) name12620 (
		_w12646_,
		_w12651_,
		_w12652_,
		_w12654_
	);
	LUT4 #(
		.INIT('h009a)
	) name12621 (
		\a[8] ,
		_w12626_,
		_w12630_,
		_w12632_,
		_w12655_
	);
	LUT4 #(
		.INIT('h9a65)
	) name12622 (
		\a[8] ,
		_w12626_,
		_w12630_,
		_w12632_,
		_w12656_
	);
	LUT3 #(
		.INIT('h54)
	) name12623 (
		_w12633_,
		_w12654_,
		_w12655_,
		_w12657_
	);
	LUT4 #(
		.INIT('h009a)
	) name12624 (
		\a[8] ,
		_w12617_,
		_w12622_,
		_w12624_,
		_w12658_
	);
	LUT4 #(
		.INIT('h9a65)
	) name12625 (
		\a[8] ,
		_w12617_,
		_w12622_,
		_w12624_,
		_w12659_
	);
	LUT3 #(
		.INIT('h54)
	) name12626 (
		_w12625_,
		_w12657_,
		_w12658_,
		_w12660_
	);
	LUT2 #(
		.INIT('h2)
	) name12627 (
		_w12614_,
		_w12615_,
		_w12661_
	);
	LUT2 #(
		.INIT('h9)
	) name12628 (
		_w12614_,
		_w12615_,
		_w12662_
	);
	LUT4 #(
		.INIT('h9a65)
	) name12629 (
		\a[8] ,
		_w12604_,
		_w12608_,
		_w12609_,
		_w12663_
	);
	LUT4 #(
		.INIT('h4d00)
	) name12630 (
		_w12614_,
		_w12615_,
		_w12660_,
		_w12663_,
		_w12664_
	);
	LUT4 #(
		.INIT('h9699)
	) name12631 (
		\a[8] ,
		_w12596_,
		_w12597_,
		_w12602_,
		_w12665_
	);
	LUT4 #(
		.INIT('h0155)
	) name12632 (
		_w12603_,
		_w12610_,
		_w12664_,
		_w12665_,
		_w12666_
	);
	LUT2 #(
		.INIT('h4)
	) name12633 (
		_w12590_,
		_w12594_,
		_w12667_
	);
	LUT2 #(
		.INIT('h9)
	) name12634 (
		_w12590_,
		_w12594_,
		_w12668_
	);
	LUT3 #(
		.INIT('h54)
	) name12635 (
		_w12595_,
		_w12666_,
		_w12667_,
		_w12669_
	);
	LUT3 #(
		.INIT('h12)
	) name12636 (
		\a[8] ,
		_w12584_,
		_w12588_,
		_w12670_
	);
	LUT3 #(
		.INIT('h69)
	) name12637 (
		\a[8] ,
		_w12584_,
		_w12588_,
		_w12671_
	);
	LUT3 #(
		.INIT('h54)
	) name12638 (
		_w12589_,
		_w12669_,
		_w12670_,
		_w12672_
	);
	LUT3 #(
		.INIT('h06)
	) name12639 (
		\a[8] ,
		_w12581_,
		_w12582_,
		_w12673_
	);
	LUT3 #(
		.INIT('h69)
	) name12640 (
		\a[8] ,
		_w12581_,
		_w12582_,
		_w12674_
	);
	LUT3 #(
		.INIT('h54)
	) name12641 (
		_w12583_,
		_w12672_,
		_w12673_,
		_w12675_
	);
	LUT3 #(
		.INIT('h06)
	) name12642 (
		\a[8] ,
		_w12575_,
		_w12576_,
		_w12676_
	);
	LUT3 #(
		.INIT('h69)
	) name12643 (
		\a[8] ,
		_w12575_,
		_w12576_,
		_w12677_
	);
	LUT3 #(
		.INIT('h54)
	) name12644 (
		_w12577_,
		_w12675_,
		_w12676_,
		_w12678_
	);
	LUT3 #(
		.INIT('h06)
	) name12645 (
		\a[8] ,
		_w12569_,
		_w12570_,
		_w12679_
	);
	LUT3 #(
		.INIT('h69)
	) name12646 (
		\a[8] ,
		_w12569_,
		_w12570_,
		_w12680_
	);
	LUT3 #(
		.INIT('h54)
	) name12647 (
		_w12571_,
		_w12678_,
		_w12679_,
		_w12681_
	);
	LUT2 #(
		.INIT('h4)
	) name12648 (
		_w12560_,
		_w12564_,
		_w12682_
	);
	LUT2 #(
		.INIT('h9)
	) name12649 (
		_w12560_,
		_w12564_,
		_w12683_
	);
	LUT4 #(
		.INIT('h9699)
	) name12650 (
		\a[8] ,
		_w12553_,
		_w12554_,
		_w12558_,
		_w12684_
	);
	LUT4 #(
		.INIT('h2b00)
	) name12651 (
		_w12560_,
		_w12564_,
		_w12681_,
		_w12684_,
		_w12685_
	);
	LUT4 #(
		.INIT('h9699)
	) name12652 (
		\a[8] ,
		_w12545_,
		_w12546_,
		_w12551_,
		_w12686_
	);
	LUT4 #(
		.INIT('h0155)
	) name12653 (
		_w12552_,
		_w12559_,
		_w12685_,
		_w12686_,
		_w12687_
	);
	LUT2 #(
		.INIT('h2)
	) name12654 (
		_w12542_,
		_w12543_,
		_w12688_
	);
	LUT2 #(
		.INIT('h9)
	) name12655 (
		_w12542_,
		_w12543_,
		_w12689_
	);
	LUT4 #(
		.INIT('h9a65)
	) name12656 (
		\a[8] ,
		_w12532_,
		_w12536_,
		_w12537_,
		_w12690_
	);
	LUT4 #(
		.INIT('h4d00)
	) name12657 (
		_w12542_,
		_w12543_,
		_w12687_,
		_w12690_,
		_w12691_
	);
	LUT4 #(
		.INIT('h9a65)
	) name12658 (
		\a[8] ,
		_w12524_,
		_w12529_,
		_w12530_,
		_w12692_
	);
	LUT4 #(
		.INIT('h0155)
	) name12659 (
		_w12531_,
		_w12538_,
		_w12691_,
		_w12692_,
		_w12693_
	);
	LUT2 #(
		.INIT('h4)
	) name12660 (
		_w12518_,
		_w12522_,
		_w12694_
	);
	LUT2 #(
		.INIT('h9)
	) name12661 (
		_w12518_,
		_w12522_,
		_w12695_
	);
	LUT4 #(
		.INIT('h9699)
	) name12662 (
		\a[8] ,
		_w12511_,
		_w12512_,
		_w12516_,
		_w12696_
	);
	LUT4 #(
		.INIT('h2b00)
	) name12663 (
		_w12518_,
		_w12522_,
		_w12693_,
		_w12696_,
		_w12697_
	);
	LUT4 #(
		.INIT('h9699)
	) name12664 (
		\a[8] ,
		_w12503_,
		_w12504_,
		_w12509_,
		_w12698_
	);
	LUT4 #(
		.INIT('h0155)
	) name12665 (
		_w12510_,
		_w12517_,
		_w12697_,
		_w12698_,
		_w12699_
	);
	LUT2 #(
		.INIT('h2)
	) name12666 (
		_w12500_,
		_w12501_,
		_w12700_
	);
	LUT2 #(
		.INIT('h9)
	) name12667 (
		_w12500_,
		_w12501_,
		_w12701_
	);
	LUT4 #(
		.INIT('h9a65)
	) name12668 (
		\a[8] ,
		_w12490_,
		_w12494_,
		_w12495_,
		_w12702_
	);
	LUT4 #(
		.INIT('h4d00)
	) name12669 (
		_w12500_,
		_w12501_,
		_w12699_,
		_w12702_,
		_w12703_
	);
	LUT4 #(
		.INIT('h9699)
	) name12670 (
		\a[8] ,
		_w12482_,
		_w12483_,
		_w12488_,
		_w12704_
	);
	LUT4 #(
		.INIT('h0155)
	) name12671 (
		_w12489_,
		_w12496_,
		_w12703_,
		_w12704_,
		_w12705_
	);
	LUT2 #(
		.INIT('h4)
	) name12672 (
		_w12475_,
		_w12480_,
		_w12706_
	);
	LUT2 #(
		.INIT('h9)
	) name12673 (
		_w12475_,
		_w12480_,
		_w12707_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12674 (
		_w4459_,
		_w11390_,
		_w11482_,
		_w11483_,
		_w12708_
	);
	LUT4 #(
		.INIT('h2228)
	) name12675 (
		_w4700_,
		_w7935_,
		_w8077_,
		_w11279_,
		_w12709_
	);
	LUT3 #(
		.INIT('h82)
	) name12676 (
		_w4458_,
		_w11274_,
		_w11276_,
		_w12710_
	);
	LUT3 #(
		.INIT('h07)
	) name12677 (
		_w4684_,
		_w11388_,
		_w12710_,
		_w12711_
	);
	LUT2 #(
		.INIT('h4)
	) name12678 (
		_w12709_,
		_w12711_,
		_w12712_
	);
	LUT3 #(
		.INIT('h82)
	) name12679 (
		_w3710_,
		_w11469_,
		_w11471_,
		_w12713_
	);
	LUT4 #(
		.INIT('h2228)
	) name12680 (
		_w3886_,
		_w8794_,
		_w8994_,
		_w11267_,
		_w12714_
	);
	LUT3 #(
		.INIT('h82)
	) name12681 (
		_w3709_,
		_w11262_,
		_w11264_,
		_w12715_
	);
	LUT3 #(
		.INIT('h07)
	) name12682 (
		_w3877_,
		_w11400_,
		_w12715_,
		_w12716_
	);
	LUT2 #(
		.INIT('h4)
	) name12683 (
		_w12714_,
		_w12716_,
		_w12717_
	);
	LUT3 #(
		.INIT('h32)
	) name12684 (
		_w12403_,
		_w12448_,
		_w12449_,
		_w12718_
	);
	LUT3 #(
		.INIT('h82)
	) name12685 (
		_w3214_,
		_w10599_,
		_w11253_,
		_w12719_
	);
	LUT4 #(
		.INIT('h007d)
	) name12686 (
		_w3249_,
		_w10580_,
		_w11254_,
		_w12719_,
		_w12720_
	);
	LUT4 #(
		.INIT('h7d00)
	) name12687 (
		_w3262_,
		_w10268_,
		_w11255_,
		_w12720_,
		_w12721_
	);
	LUT4 #(
		.INIT('h7d00)
	) name12688 (
		_w37_,
		_w11456_,
		_w11458_,
		_w12721_,
		_w12722_
	);
	LUT4 #(
		.INIT('h010f)
	) name12689 (
		_w12172_,
		_w12174_,
		_w12445_,
		_w12446_,
		_w12723_
	);
	LUT3 #(
		.INIT('h32)
	) name12690 (
		_w12408_,
		_w12435_,
		_w12436_,
		_w12724_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12691 (
		_w2549_,
		_w10968_,
		_w11238_,
		_w11240_,
		_w12725_
	);
	LUT4 #(
		.INIT('h007d)
	) name12692 (
		_w2617_,
		_w11241_,
		_w11243_,
		_w12725_,
		_w12726_
	);
	LUT3 #(
		.INIT('h70)
	) name12693 (
		_w2854_,
		_w11421_,
		_w12726_,
		_w12727_
	);
	LUT4 #(
		.INIT('h95aa)
	) name12694 (
		\a[29] ,
		_w2550_,
		_w11569_,
		_w12727_,
		_w12728_
	);
	LUT3 #(
		.INIT('h54)
	) name12695 (
		_w12425_,
		_w12426_,
		_w12433_,
		_w12729_
	);
	LUT4 #(
		.INIT('h153f)
	) name12696 (
		_w38_,
		_w43_,
		_w65_,
		_w158_,
		_w12730_
	);
	LUT4 #(
		.INIT('h8000)
	) name12697 (
		_w555_,
		_w772_,
		_w790_,
		_w12730_,
		_w12731_
	);
	LUT3 #(
		.INIT('h57)
	) name12698 (
		_w90_,
		_w166_,
		_w419_,
		_w12732_
	);
	LUT4 #(
		.INIT('h8000)
	) name12699 (
		_w116_,
		_w343_,
		_w663_,
		_w12732_,
		_w12733_
	);
	LUT3 #(
		.INIT('h80)
	) name12700 (
		_w1450_,
		_w1811_,
		_w7445_,
		_w12734_
	);
	LUT4 #(
		.INIT('h8000)
	) name12701 (
		_w1640_,
		_w12734_,
		_w12731_,
		_w12733_,
		_w12735_
	);
	LUT4 #(
		.INIT('h8000)
	) name12702 (
		_w2912_,
		_w2915_,
		_w3588_,
		_w3591_,
		_w12736_
	);
	LUT2 #(
		.INIT('h8)
	) name12703 (
		_w12735_,
		_w12736_,
		_w12737_
	);
	LUT3 #(
		.INIT('h80)
	) name12704 (
		_w1202_,
		_w1799_,
		_w12737_,
		_w12738_
	);
	LUT3 #(
		.INIT('h28)
	) name12705 (
		_w377_,
		_w11431_,
		_w11435_,
		_w12739_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12706 (
		_w376_,
		_w10991_,
		_w11230_,
		_w11232_,
		_w12740_
	);
	LUT4 #(
		.INIT('h007d)
	) name12707 (
		_w2407_,
		_w11233_,
		_w11235_,
		_w12740_,
		_w12741_
	);
	LUT3 #(
		.INIT('h70)
	) name12708 (
		_w2527_,
		_w11427_,
		_w12741_,
		_w12742_
	);
	LUT3 #(
		.INIT('h45)
	) name12709 (
		_w12738_,
		_w12739_,
		_w12742_,
		_w12743_
	);
	LUT3 #(
		.INIT('h20)
	) name12710 (
		_w12738_,
		_w12739_,
		_w12742_,
		_w12744_
	);
	LUT3 #(
		.INIT('h9a)
	) name12711 (
		_w12738_,
		_w12739_,
		_w12742_,
		_w12745_
	);
	LUT2 #(
		.INIT('h9)
	) name12712 (
		_w12729_,
		_w12745_,
		_w12746_
	);
	LUT2 #(
		.INIT('h4)
	) name12713 (
		_w12728_,
		_w12746_,
		_w12747_
	);
	LUT2 #(
		.INIT('h2)
	) name12714 (
		_w12728_,
		_w12746_,
		_w12748_
	);
	LUT2 #(
		.INIT('h9)
	) name12715 (
		_w12728_,
		_w12746_,
		_w12749_
	);
	LUT2 #(
		.INIT('h9)
	) name12716 (
		_w12724_,
		_w12749_,
		_w12750_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12717 (
		_w2874_,
		_w10945_,
		_w11246_,
		_w11248_,
		_w12751_
	);
	LUT4 #(
		.INIT('h007d)
	) name12718 (
		_w2975_,
		_w11249_,
		_w11251_,
		_w12751_,
		_w12752_
	);
	LUT3 #(
		.INIT('h70)
	) name12719 (
		_w2986_,
		_w11415_,
		_w12752_,
		_w12753_
	);
	LUT4 #(
		.INIT('h95aa)
	) name12720 (
		\a[26] ,
		_w2875_,
		_w11675_,
		_w12753_,
		_w12754_
	);
	LUT2 #(
		.INIT('h2)
	) name12721 (
		_w12750_,
		_w12754_,
		_w12755_
	);
	LUT2 #(
		.INIT('h4)
	) name12722 (
		_w12750_,
		_w12754_,
		_w12756_
	);
	LUT2 #(
		.INIT('h9)
	) name12723 (
		_w12750_,
		_w12754_,
		_w12757_
	);
	LUT2 #(
		.INIT('h9)
	) name12724 (
		_w12723_,
		_w12757_,
		_w12758_
	);
	LUT3 #(
		.INIT('h90)
	) name12725 (
		\a[23] ,
		_w12722_,
		_w12758_,
		_w12759_
	);
	LUT3 #(
		.INIT('h06)
	) name12726 (
		\a[23] ,
		_w12722_,
		_w12758_,
		_w12760_
	);
	LUT3 #(
		.INIT('h69)
	) name12727 (
		\a[23] ,
		_w12722_,
		_w12758_,
		_w12761_
	);
	LUT2 #(
		.INIT('h9)
	) name12728 (
		_w12718_,
		_w12761_,
		_w12762_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12729 (
		_w3312_,
		_w11408_,
		_w11463_,
		_w11464_,
		_w12763_
	);
	LUT4 #(
		.INIT('h2228)
	) name12730 (
		_w3654_,
		_w9446_,
		_w9702_,
		_w11261_,
		_w12764_
	);
	LUT3 #(
		.INIT('h82)
	) name12731 (
		_w3311_,
		_w11256_,
		_w11258_,
		_w12765_
	);
	LUT3 #(
		.INIT('h07)
	) name12732 (
		_w3645_,
		_w11406_,
		_w12765_,
		_w12766_
	);
	LUT2 #(
		.INIT('h4)
	) name12733 (
		_w12764_,
		_w12766_,
		_w12767_
	);
	LUT4 #(
		.INIT('h4844)
	) name12734 (
		\a[20] ,
		_w12762_,
		_w12763_,
		_w12767_,
		_w12768_
	);
	LUT4 #(
		.INIT('h9699)
	) name12735 (
		\a[20] ,
		_w12762_,
		_w12763_,
		_w12767_,
		_w12769_
	);
	LUT4 #(
		.INIT('h4d00)
	) name12736 (
		_w12402_,
		_w12451_,
		_w12455_,
		_w12769_,
		_w12770_
	);
	LUT4 #(
		.INIT('h32cd)
	) name12737 (
		_w12402_,
		_w12456_,
		_w12457_,
		_w12769_,
		_w12771_
	);
	LUT4 #(
		.INIT('h6500)
	) name12738 (
		\a[17] ,
		_w12713_,
		_w12717_,
		_w12771_,
		_w12772_
	);
	LUT4 #(
		.INIT('h9a65)
	) name12739 (
		\a[17] ,
		_w12713_,
		_w12717_,
		_w12771_,
		_w12773_
	);
	LUT4 #(
		.INIT('h7100)
	) name12740 (
		_w12397_,
		_w12401_,
		_w12459_,
		_w12773_,
		_w12774_
	);
	LUT4 #(
		.INIT('h32cd)
	) name12741 (
		_w12397_,
		_w12460_,
		_w12461_,
		_w12773_,
		_w12775_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12742 (
		_w4034_,
		_w11396_,
		_w11476_,
		_w11477_,
		_w12776_
	);
	LUT4 #(
		.INIT('h2228)
	) name12743 (
		_w4382_,
		_w8466_,
		_w8541_,
		_w11273_,
		_w12777_
	);
	LUT3 #(
		.INIT('h82)
	) name12744 (
		_w4033_,
		_w11268_,
		_w11270_,
		_w12778_
	);
	LUT3 #(
		.INIT('h07)
	) name12745 (
		_w4367_,
		_w11394_,
		_w12778_,
		_w12779_
	);
	LUT2 #(
		.INIT('h4)
	) name12746 (
		_w12777_,
		_w12779_,
		_w12780_
	);
	LUT4 #(
		.INIT('h4844)
	) name12747 (
		\a[14] ,
		_w12775_,
		_w12776_,
		_w12780_,
		_w12781_
	);
	LUT4 #(
		.INIT('h9699)
	) name12748 (
		\a[14] ,
		_w12775_,
		_w12776_,
		_w12780_,
		_w12782_
	);
	LUT4 #(
		.INIT('h4d00)
	) name12749 (
		_w12396_,
		_w12463_,
		_w12467_,
		_w12782_,
		_w12783_
	);
	LUT4 #(
		.INIT('h32cd)
	) name12750 (
		_w12396_,
		_w12468_,
		_w12469_,
		_w12782_,
		_w12784_
	);
	LUT4 #(
		.INIT('h6500)
	) name12751 (
		\a[11] ,
		_w12708_,
		_w12712_,
		_w12784_,
		_w12785_
	);
	LUT4 #(
		.INIT('h9a65)
	) name12752 (
		\a[11] ,
		_w12708_,
		_w12712_,
		_w12784_,
		_w12786_
	);
	LUT4 #(
		.INIT('h7100)
	) name12753 (
		_w12390_,
		_w12395_,
		_w12471_,
		_w12786_,
		_w12787_
	);
	LUT4 #(
		.INIT('h32cd)
	) name12754 (
		_w12390_,
		_w12472_,
		_w12473_,
		_w12786_,
		_w12788_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12755 (
		_w4876_,
		_w11384_,
		_w11488_,
		_w11489_,
		_w12789_
	);
	LUT4 #(
		.INIT('h2228)
	) name12756 (
		_w5286_,
		_w7695_,
		_w7750_,
		_w11285_,
		_w12790_
	);
	LUT3 #(
		.INIT('h82)
	) name12757 (
		_w4875_,
		_w11280_,
		_w11282_,
		_w12791_
	);
	LUT3 #(
		.INIT('h07)
	) name12758 (
		_w5271_,
		_w11382_,
		_w12791_,
		_w12792_
	);
	LUT2 #(
		.INIT('h4)
	) name12759 (
		_w12790_,
		_w12792_,
		_w12793_
	);
	LUT4 #(
		.INIT('h4844)
	) name12760 (
		\a[8] ,
		_w12788_,
		_w12789_,
		_w12793_,
		_w12794_
	);
	LUT4 #(
		.INIT('h9699)
	) name12761 (
		\a[8] ,
		_w12788_,
		_w12789_,
		_w12793_,
		_w12795_
	);
	LUT4 #(
		.INIT('h2b00)
	) name12762 (
		_w12475_,
		_w12480_,
		_w12705_,
		_w12795_,
		_w12796_
	);
	LUT4 #(
		.INIT('h54ab)
	) name12763 (
		_w12481_,
		_w12705_,
		_w12706_,
		_w12795_,
		_w12797_
	);
	LUT4 #(
		.INIT('h6500)
	) name12764 (
		\a[5] ,
		_w11553_,
		_w11557_,
		_w12797_,
		_w12798_
	);
	LUT4 #(
		.INIT('h54ab)
	) name12765 (
		_w11380_,
		_w11490_,
		_w11491_,
		_w11493_,
		_w12799_
	);
	LUT4 #(
		.INIT('h2228)
	) name12766 (
		_w5524_,
		_w7695_,
		_w7750_,
		_w11285_,
		_w12800_
	);
	LUT4 #(
		.INIT('h007d)
	) name12767 (
		_w6031_,
		_w11286_,
		_w11335_,
		_w12800_,
		_w12801_
	);
	LUT3 #(
		.INIT('h70)
	) name12768 (
		_w6324_,
		_w11377_,
		_w12801_,
		_w12802_
	);
	LUT4 #(
		.INIT('h95aa)
	) name12769 (
		\a[5] ,
		_w35_,
		_w12799_,
		_w12802_,
		_w12803_
	);
	LUT2 #(
		.INIT('h9)
	) name12770 (
		_w12705_,
		_w12707_,
		_w12804_
	);
	LUT2 #(
		.INIT('h4)
	) name12771 (
		_w12803_,
		_w12804_,
		_w12805_
	);
	LUT3 #(
		.INIT('h82)
	) name12772 (
		_w35_,
		_w11490_,
		_w11492_,
		_w12806_
	);
	LUT3 #(
		.INIT('h82)
	) name12773 (
		_w6324_,
		_w11286_,
		_w11335_,
		_w12807_
	);
	LUT2 #(
		.INIT('h8)
	) name12774 (
		_w5524_,
		_w11382_,
		_w12808_
	);
	LUT4 #(
		.INIT('h2228)
	) name12775 (
		_w6031_,
		_w7695_,
		_w7750_,
		_w11285_,
		_w12809_
	);
	LUT2 #(
		.INIT('h1)
	) name12776 (
		_w12808_,
		_w12809_,
		_w12810_
	);
	LUT2 #(
		.INIT('h4)
	) name12777 (
		_w12807_,
		_w12810_,
		_w12811_
	);
	LUT3 #(
		.INIT('h1e)
	) name12778 (
		_w12496_,
		_w12703_,
		_w12704_,
		_w12812_
	);
	LUT4 #(
		.INIT('h6500)
	) name12779 (
		\a[5] ,
		_w12806_,
		_w12811_,
		_w12812_,
		_w12813_
	);
	LUT4 #(
		.INIT('h54ab)
	) name12780 (
		_w12502_,
		_w12699_,
		_w12700_,
		_w12702_,
		_w12814_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12781 (
		_w35_,
		_w11384_,
		_w11488_,
		_w11489_,
		_w12815_
	);
	LUT4 #(
		.INIT('h2228)
	) name12782 (
		_w6324_,
		_w7695_,
		_w7750_,
		_w11285_,
		_w12816_
	);
	LUT3 #(
		.INIT('h82)
	) name12783 (
		_w5524_,
		_w11280_,
		_w11282_,
		_w12817_
	);
	LUT3 #(
		.INIT('h07)
	) name12784 (
		_w6031_,
		_w11382_,
		_w12817_,
		_w12818_
	);
	LUT2 #(
		.INIT('h4)
	) name12785 (
		_w12816_,
		_w12818_,
		_w12819_
	);
	LUT4 #(
		.INIT('h4844)
	) name12786 (
		\a[5] ,
		_w12814_,
		_w12815_,
		_w12819_,
		_w12820_
	);
	LUT2 #(
		.INIT('h9)
	) name12787 (
		_w12699_,
		_w12701_,
		_w12821_
	);
	LUT4 #(
		.INIT('h2228)
	) name12788 (
		_w5524_,
		_w7935_,
		_w8077_,
		_w11279_,
		_w12822_
	);
	LUT4 #(
		.INIT('h007d)
	) name12789 (
		_w6031_,
		_w11280_,
		_w11282_,
		_w12822_,
		_w12823_
	);
	LUT3 #(
		.INIT('h70)
	) name12790 (
		_w6324_,
		_w11382_,
		_w12823_,
		_w12824_
	);
	LUT4 #(
		.INIT('h95aa)
	) name12791 (
		\a[5] ,
		_w35_,
		_w12476_,
		_w12824_,
		_w12825_
	);
	LUT2 #(
		.INIT('h2)
	) name12792 (
		_w12821_,
		_w12825_,
		_w12826_
	);
	LUT3 #(
		.INIT('h82)
	) name12793 (
		_w35_,
		_w11484_,
		_w11486_,
		_w12827_
	);
	LUT3 #(
		.INIT('h82)
	) name12794 (
		_w6324_,
		_w11280_,
		_w11282_,
		_w12828_
	);
	LUT2 #(
		.INIT('h8)
	) name12795 (
		_w5524_,
		_w11388_,
		_w12829_
	);
	LUT4 #(
		.INIT('h2228)
	) name12796 (
		_w6031_,
		_w7935_,
		_w8077_,
		_w11279_,
		_w12830_
	);
	LUT2 #(
		.INIT('h1)
	) name12797 (
		_w12829_,
		_w12830_,
		_w12831_
	);
	LUT2 #(
		.INIT('h4)
	) name12798 (
		_w12828_,
		_w12831_,
		_w12832_
	);
	LUT3 #(
		.INIT('h1e)
	) name12799 (
		_w12517_,
		_w12697_,
		_w12698_,
		_w12833_
	);
	LUT4 #(
		.INIT('h6500)
	) name12800 (
		\a[5] ,
		_w12827_,
		_w12832_,
		_w12833_,
		_w12834_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12801 (
		_w35_,
		_w11390_,
		_w11482_,
		_w11483_,
		_w12835_
	);
	LUT4 #(
		.INIT('h2228)
	) name12802 (
		_w6324_,
		_w7935_,
		_w8077_,
		_w11279_,
		_w12836_
	);
	LUT3 #(
		.INIT('h82)
	) name12803 (
		_w5524_,
		_w11274_,
		_w11276_,
		_w12837_
	);
	LUT3 #(
		.INIT('h07)
	) name12804 (
		_w6031_,
		_w11388_,
		_w12837_,
		_w12838_
	);
	LUT2 #(
		.INIT('h4)
	) name12805 (
		_w12836_,
		_w12838_,
		_w12839_
	);
	LUT4 #(
		.INIT('h54ab)
	) name12806 (
		_w12523_,
		_w12693_,
		_w12694_,
		_w12696_,
		_w12840_
	);
	LUT4 #(
		.INIT('h6500)
	) name12807 (
		\a[5] ,
		_w12835_,
		_w12839_,
		_w12840_,
		_w12841_
	);
	LUT4 #(
		.INIT('h2228)
	) name12808 (
		_w5524_,
		_w8466_,
		_w8541_,
		_w11273_,
		_w12842_
	);
	LUT4 #(
		.INIT('h007d)
	) name12809 (
		_w6031_,
		_w11274_,
		_w11276_,
		_w12842_,
		_w12843_
	);
	LUT3 #(
		.INIT('h70)
	) name12810 (
		_w6324_,
		_w11388_,
		_w12843_,
		_w12844_
	);
	LUT4 #(
		.INIT('h95aa)
	) name12811 (
		\a[5] ,
		_w35_,
		_w12391_,
		_w12844_,
		_w12845_
	);
	LUT2 #(
		.INIT('h9)
	) name12812 (
		_w12693_,
		_w12695_,
		_w12846_
	);
	LUT2 #(
		.INIT('h4)
	) name12813 (
		_w12845_,
		_w12846_,
		_w12847_
	);
	LUT3 #(
		.INIT('h1e)
	) name12814 (
		_w12538_,
		_w12691_,
		_w12692_,
		_w12848_
	);
	LUT3 #(
		.INIT('h82)
	) name12815 (
		_w35_,
		_w11478_,
		_w11480_,
		_w12849_
	);
	LUT3 #(
		.INIT('h82)
	) name12816 (
		_w6324_,
		_w11274_,
		_w11276_,
		_w12850_
	);
	LUT2 #(
		.INIT('h8)
	) name12817 (
		_w5524_,
		_w11394_,
		_w12851_
	);
	LUT4 #(
		.INIT('h2228)
	) name12818 (
		_w6031_,
		_w8466_,
		_w8541_,
		_w11273_,
		_w12852_
	);
	LUT2 #(
		.INIT('h1)
	) name12819 (
		_w12851_,
		_w12852_,
		_w12853_
	);
	LUT2 #(
		.INIT('h4)
	) name12820 (
		_w12850_,
		_w12853_,
		_w12854_
	);
	LUT4 #(
		.INIT('h4844)
	) name12821 (
		\a[5] ,
		_w12848_,
		_w12849_,
		_w12854_,
		_w12855_
	);
	LUT4 #(
		.INIT('h54ab)
	) name12822 (
		_w12544_,
		_w12687_,
		_w12688_,
		_w12690_,
		_w12856_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12823 (
		_w35_,
		_w11396_,
		_w11476_,
		_w11477_,
		_w12857_
	);
	LUT4 #(
		.INIT('h2228)
	) name12824 (
		_w6324_,
		_w8466_,
		_w8541_,
		_w11273_,
		_w12858_
	);
	LUT3 #(
		.INIT('h82)
	) name12825 (
		_w5524_,
		_w11268_,
		_w11270_,
		_w12859_
	);
	LUT3 #(
		.INIT('h07)
	) name12826 (
		_w6031_,
		_w11394_,
		_w12859_,
		_w12860_
	);
	LUT2 #(
		.INIT('h4)
	) name12827 (
		_w12858_,
		_w12860_,
		_w12861_
	);
	LUT4 #(
		.INIT('h4844)
	) name12828 (
		\a[5] ,
		_w12856_,
		_w12857_,
		_w12861_,
		_w12862_
	);
	LUT2 #(
		.INIT('h9)
	) name12829 (
		_w12687_,
		_w12689_,
		_w12863_
	);
	LUT4 #(
		.INIT('h2228)
	) name12830 (
		_w5524_,
		_w8794_,
		_w8994_,
		_w11267_,
		_w12864_
	);
	LUT4 #(
		.INIT('h007d)
	) name12831 (
		_w6031_,
		_w11268_,
		_w11270_,
		_w12864_,
		_w12865_
	);
	LUT3 #(
		.INIT('h70)
	) name12832 (
		_w6324_,
		_w11394_,
		_w12865_,
		_w12866_
	);
	LUT4 #(
		.INIT('h95aa)
	) name12833 (
		\a[5] ,
		_w35_,
		_w12209_,
		_w12866_,
		_w12867_
	);
	LUT2 #(
		.INIT('h2)
	) name12834 (
		_w12863_,
		_w12867_,
		_w12868_
	);
	LUT3 #(
		.INIT('h82)
	) name12835 (
		_w35_,
		_w11472_,
		_w11474_,
		_w12869_
	);
	LUT3 #(
		.INIT('h82)
	) name12836 (
		_w6324_,
		_w11268_,
		_w11270_,
		_w12870_
	);
	LUT2 #(
		.INIT('h8)
	) name12837 (
		_w5524_,
		_w11400_,
		_w12871_
	);
	LUT4 #(
		.INIT('h2228)
	) name12838 (
		_w6031_,
		_w8794_,
		_w8994_,
		_w11267_,
		_w12872_
	);
	LUT2 #(
		.INIT('h1)
	) name12839 (
		_w12871_,
		_w12872_,
		_w12873_
	);
	LUT2 #(
		.INIT('h4)
	) name12840 (
		_w12870_,
		_w12873_,
		_w12874_
	);
	LUT3 #(
		.INIT('h1e)
	) name12841 (
		_w12559_,
		_w12685_,
		_w12686_,
		_w12875_
	);
	LUT4 #(
		.INIT('h6500)
	) name12842 (
		\a[5] ,
		_w12869_,
		_w12874_,
		_w12875_,
		_w12876_
	);
	LUT3 #(
		.INIT('h82)
	) name12843 (
		_w35_,
		_w11469_,
		_w11471_,
		_w12877_
	);
	LUT4 #(
		.INIT('h2228)
	) name12844 (
		_w6324_,
		_w8794_,
		_w8994_,
		_w11267_,
		_w12878_
	);
	LUT3 #(
		.INIT('h82)
	) name12845 (
		_w5524_,
		_w11262_,
		_w11264_,
		_w12879_
	);
	LUT3 #(
		.INIT('h07)
	) name12846 (
		_w6031_,
		_w11400_,
		_w12879_,
		_w12880_
	);
	LUT2 #(
		.INIT('h4)
	) name12847 (
		_w12878_,
		_w12880_,
		_w12881_
	);
	LUT4 #(
		.INIT('h54ab)
	) name12848 (
		_w12565_,
		_w12681_,
		_w12682_,
		_w12684_,
		_w12882_
	);
	LUT4 #(
		.INIT('h6500)
	) name12849 (
		\a[5] ,
		_w12877_,
		_w12881_,
		_w12882_,
		_w12883_
	);
	LUT4 #(
		.INIT('h2228)
	) name12850 (
		_w5524_,
		_w9446_,
		_w9702_,
		_w11261_,
		_w12884_
	);
	LUT4 #(
		.INIT('h007d)
	) name12851 (
		_w6031_,
		_w11262_,
		_w11264_,
		_w12884_,
		_w12885_
	);
	LUT3 #(
		.INIT('h70)
	) name12852 (
		_w6324_,
		_w11400_,
		_w12885_,
		_w12886_
	);
	LUT4 #(
		.INIT('h95aa)
	) name12853 (
		\a[5] ,
		_w35_,
		_w11967_,
		_w12886_,
		_w12887_
	);
	LUT2 #(
		.INIT('h9)
	) name12854 (
		_w12681_,
		_w12683_,
		_w12888_
	);
	LUT2 #(
		.INIT('h4)
	) name12855 (
		_w12887_,
		_w12888_,
		_w12889_
	);
	LUT2 #(
		.INIT('h9)
	) name12856 (
		_w12678_,
		_w12680_,
		_w12890_
	);
	LUT3 #(
		.INIT('h82)
	) name12857 (
		_w35_,
		_w11465_,
		_w11467_,
		_w12891_
	);
	LUT3 #(
		.INIT('h82)
	) name12858 (
		_w6324_,
		_w11262_,
		_w11264_,
		_w12892_
	);
	LUT2 #(
		.INIT('h8)
	) name12859 (
		_w5524_,
		_w11406_,
		_w12893_
	);
	LUT4 #(
		.INIT('h2228)
	) name12860 (
		_w6031_,
		_w9446_,
		_w9702_,
		_w11261_,
		_w12894_
	);
	LUT2 #(
		.INIT('h1)
	) name12861 (
		_w12893_,
		_w12894_,
		_w12895_
	);
	LUT2 #(
		.INIT('h4)
	) name12862 (
		_w12892_,
		_w12895_,
		_w12896_
	);
	LUT4 #(
		.INIT('h4844)
	) name12863 (
		\a[5] ,
		_w12890_,
		_w12891_,
		_w12896_,
		_w12897_
	);
	LUT2 #(
		.INIT('h9)
	) name12864 (
		_w12675_,
		_w12677_,
		_w12898_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12865 (
		_w35_,
		_w11408_,
		_w11463_,
		_w11464_,
		_w12899_
	);
	LUT4 #(
		.INIT('h2228)
	) name12866 (
		_w6324_,
		_w9446_,
		_w9702_,
		_w11261_,
		_w12900_
	);
	LUT3 #(
		.INIT('h82)
	) name12867 (
		_w5524_,
		_w11256_,
		_w11258_,
		_w12901_
	);
	LUT3 #(
		.INIT('h07)
	) name12868 (
		_w6031_,
		_w11406_,
		_w12901_,
		_w12902_
	);
	LUT2 #(
		.INIT('h4)
	) name12869 (
		_w12900_,
		_w12902_,
		_w12903_
	);
	LUT4 #(
		.INIT('h4844)
	) name12870 (
		\a[5] ,
		_w12898_,
		_w12899_,
		_w12903_,
		_w12904_
	);
	LUT2 #(
		.INIT('h9)
	) name12871 (
		_w12672_,
		_w12674_,
		_w12905_
	);
	LUT3 #(
		.INIT('h82)
	) name12872 (
		_w5524_,
		_w10268_,
		_w11255_,
		_w12906_
	);
	LUT4 #(
		.INIT('h007d)
	) name12873 (
		_w6031_,
		_w11256_,
		_w11258_,
		_w12906_,
		_w12907_
	);
	LUT3 #(
		.INIT('h70)
	) name12874 (
		_w6324_,
		_w11406_,
		_w12907_,
		_w12908_
	);
	LUT4 #(
		.INIT('h95aa)
	) name12875 (
		\a[5] ,
		_w35_,
		_w11796_,
		_w12908_,
		_w12909_
	);
	LUT2 #(
		.INIT('h2)
	) name12876 (
		_w12905_,
		_w12909_,
		_w12910_
	);
	LUT3 #(
		.INIT('h82)
	) name12877 (
		_w5524_,
		_w10580_,
		_w11254_,
		_w12911_
	);
	LUT4 #(
		.INIT('h007d)
	) name12878 (
		_w6031_,
		_w10268_,
		_w11255_,
		_w12911_,
		_w12912_
	);
	LUT4 #(
		.INIT('h7d00)
	) name12879 (
		_w6324_,
		_w11256_,
		_w11258_,
		_w12912_,
		_w12913_
	);
	LUT4 #(
		.INIT('h7d00)
	) name12880 (
		_w35_,
		_w11459_,
		_w11461_,
		_w12913_,
		_w12914_
	);
	LUT2 #(
		.INIT('h9)
	) name12881 (
		_w12669_,
		_w12671_,
		_w12915_
	);
	LUT3 #(
		.INIT('h90)
	) name12882 (
		\a[5] ,
		_w12914_,
		_w12915_,
		_w12916_
	);
	LUT3 #(
		.INIT('h82)
	) name12883 (
		_w5524_,
		_w10599_,
		_w11253_,
		_w12917_
	);
	LUT4 #(
		.INIT('h007d)
	) name12884 (
		_w6031_,
		_w10580_,
		_w11254_,
		_w12917_,
		_w12918_
	);
	LUT4 #(
		.INIT('h7d00)
	) name12885 (
		_w6324_,
		_w10268_,
		_w11255_,
		_w12918_,
		_w12919_
	);
	LUT4 #(
		.INIT('h7d00)
	) name12886 (
		_w35_,
		_w11456_,
		_w11458_,
		_w12919_,
		_w12920_
	);
	LUT2 #(
		.INIT('h9)
	) name12887 (
		_w12666_,
		_w12668_,
		_w12921_
	);
	LUT3 #(
		.INIT('h90)
	) name12888 (
		\a[5] ,
		_w12920_,
		_w12921_,
		_w12922_
	);
	LUT2 #(
		.INIT('h8)
	) name12889 (
		_w5524_,
		_w11415_,
		_w12923_
	);
	LUT4 #(
		.INIT('h007d)
	) name12890 (
		_w6031_,
		_w10599_,
		_w11253_,
		_w12923_,
		_w12924_
	);
	LUT4 #(
		.INIT('h7d00)
	) name12891 (
		_w6324_,
		_w10580_,
		_w11254_,
		_w12924_,
		_w12925_
	);
	LUT4 #(
		.INIT('h7d00)
	) name12892 (
		_w35_,
		_w11453_,
		_w11455_,
		_w12925_,
		_w12926_
	);
	LUT3 #(
		.INIT('h1e)
	) name12893 (
		_w12610_,
		_w12664_,
		_w12665_,
		_w12927_
	);
	LUT3 #(
		.INIT('h90)
	) name12894 (
		\a[5] ,
		_w12926_,
		_w12927_,
		_w12928_
	);
	LUT4 #(
		.INIT('h54ab)
	) name12895 (
		_w12616_,
		_w12660_,
		_w12661_,
		_w12663_,
		_w12929_
	);
	LUT3 #(
		.INIT('h82)
	) name12896 (
		_w5524_,
		_w11249_,
		_w11251_,
		_w12930_
	);
	LUT3 #(
		.INIT('h07)
	) name12897 (
		_w6031_,
		_w11415_,
		_w12930_,
		_w12931_
	);
	LUT4 #(
		.INIT('h7d00)
	) name12898 (
		_w6324_,
		_w10599_,
		_w11253_,
		_w12931_,
		_w12932_
	);
	LUT4 #(
		.INIT('h7d00)
	) name12899 (
		_w35_,
		_w11450_,
		_w11452_,
		_w12932_,
		_w12933_
	);
	LUT3 #(
		.INIT('h84)
	) name12900 (
		\a[5] ,
		_w12929_,
		_w12933_,
		_w12934_
	);
	LUT2 #(
		.INIT('h9)
	) name12901 (
		_w12660_,
		_w12662_,
		_w12935_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12902 (
		_w5524_,
		_w10945_,
		_w11246_,
		_w11248_,
		_w12936_
	);
	LUT4 #(
		.INIT('h007d)
	) name12903 (
		_w6031_,
		_w11249_,
		_w11251_,
		_w12936_,
		_w12937_
	);
	LUT3 #(
		.INIT('h70)
	) name12904 (
		_w6324_,
		_w11415_,
		_w12937_,
		_w12938_
	);
	LUT4 #(
		.INIT('h95aa)
	) name12905 (
		\a[5] ,
		_w35_,
		_w11675_,
		_w12938_,
		_w12939_
	);
	LUT2 #(
		.INIT('h2)
	) name12906 (
		_w12935_,
		_w12939_,
		_w12940_
	);
	LUT2 #(
		.INIT('h9)
	) name12907 (
		_w12657_,
		_w12659_,
		_w12941_
	);
	LUT3 #(
		.INIT('h82)
	) name12908 (
		_w35_,
		_w11445_,
		_w11447_,
		_w12942_
	);
	LUT3 #(
		.INIT('h82)
	) name12909 (
		_w6324_,
		_w11249_,
		_w11251_,
		_w12943_
	);
	LUT2 #(
		.INIT('h8)
	) name12910 (
		_w5524_,
		_w11421_,
		_w12944_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12911 (
		_w6031_,
		_w10945_,
		_w11246_,
		_w11248_,
		_w12945_
	);
	LUT2 #(
		.INIT('h1)
	) name12912 (
		_w12944_,
		_w12945_,
		_w12946_
	);
	LUT2 #(
		.INIT('h4)
	) name12913 (
		_w12943_,
		_w12946_,
		_w12947_
	);
	LUT4 #(
		.INIT('h4844)
	) name12914 (
		\a[5] ,
		_w12941_,
		_w12942_,
		_w12947_,
		_w12948_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12915 (
		_w35_,
		_w11423_,
		_w11443_,
		_w11444_,
		_w12949_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12916 (
		_w6324_,
		_w10945_,
		_w11246_,
		_w11248_,
		_w12950_
	);
	LUT3 #(
		.INIT('h82)
	) name12917 (
		_w5524_,
		_w11241_,
		_w11243_,
		_w12951_
	);
	LUT3 #(
		.INIT('h07)
	) name12918 (
		_w6031_,
		_w11421_,
		_w12951_,
		_w12952_
	);
	LUT2 #(
		.INIT('h4)
	) name12919 (
		_w12950_,
		_w12952_,
		_w12953_
	);
	LUT2 #(
		.INIT('h9)
	) name12920 (
		_w12654_,
		_w12656_,
		_w12954_
	);
	LUT4 #(
		.INIT('h6500)
	) name12921 (
		\a[5] ,
		_w12949_,
		_w12953_,
		_w12954_,
		_w12955_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12922 (
		_w5524_,
		_w10968_,
		_w11238_,
		_w11240_,
		_w12956_
	);
	LUT4 #(
		.INIT('h007d)
	) name12923 (
		_w6031_,
		_w11241_,
		_w11243_,
		_w12956_,
		_w12957_
	);
	LUT3 #(
		.INIT('h70)
	) name12924 (
		_w6324_,
		_w11421_,
		_w12957_,
		_w12958_
	);
	LUT4 #(
		.INIT('h95aa)
	) name12925 (
		\a[5] ,
		_w35_,
		_w11569_,
		_w12958_,
		_w12959_
	);
	LUT2 #(
		.INIT('h9)
	) name12926 (
		_w12651_,
		_w12653_,
		_w12960_
	);
	LUT2 #(
		.INIT('h4)
	) name12927 (
		_w12959_,
		_w12960_,
		_w12961_
	);
	LUT3 #(
		.INIT('h82)
	) name12928 (
		_w35_,
		_w11439_,
		_w11441_,
		_w12962_
	);
	LUT3 #(
		.INIT('h82)
	) name12929 (
		_w6324_,
		_w11241_,
		_w11243_,
		_w12963_
	);
	LUT2 #(
		.INIT('h8)
	) name12930 (
		_w5524_,
		_w11427_,
		_w12964_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12931 (
		_w6031_,
		_w10968_,
		_w11238_,
		_w11240_,
		_w12965_
	);
	LUT2 #(
		.INIT('h1)
	) name12932 (
		_w12964_,
		_w12965_,
		_w12966_
	);
	LUT2 #(
		.INIT('h4)
	) name12933 (
		_w12963_,
		_w12966_,
		_w12967_
	);
	LUT3 #(
		.INIT('h8a)
	) name12934 (
		\a[8] ,
		_w12637_,
		_w12636_,
		_w12968_
	);
	LUT2 #(
		.INIT('h9)
	) name12935 (
		_w12645_,
		_w12968_,
		_w12969_
	);
	LUT4 #(
		.INIT('h6500)
	) name12936 (
		\a[5] ,
		_w12962_,
		_w12967_,
		_w12969_,
		_w12970_
	);
	LUT3 #(
		.INIT('h82)
	) name12937 (
		_w35_,
		_w11436_,
		_w11438_,
		_w12971_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12938 (
		_w6324_,
		_w10968_,
		_w11238_,
		_w11240_,
		_w12972_
	);
	LUT3 #(
		.INIT('h82)
	) name12939 (
		_w5524_,
		_w11233_,
		_w11235_,
		_w12973_
	);
	LUT3 #(
		.INIT('h07)
	) name12940 (
		_w6031_,
		_w11427_,
		_w12973_,
		_w12974_
	);
	LUT2 #(
		.INIT('h4)
	) name12941 (
		_w12972_,
		_w12974_,
		_w12975_
	);
	LUT3 #(
		.INIT('h20)
	) name12942 (
		\a[8] ,
		_w4874_,
		_w11434_,
		_w12976_
	);
	LUT2 #(
		.INIT('h9)
	) name12943 (
		_w12636_,
		_w12976_,
		_w12977_
	);
	LUT4 #(
		.INIT('h6500)
	) name12944 (
		\a[5] ,
		_w12971_,
		_w12975_,
		_w12977_,
		_w12978_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12945 (
		_w6324_,
		_w10991_,
		_w11230_,
		_w11232_,
		_w12979_
	);
	LUT2 #(
		.INIT('h8)
	) name12946 (
		_w6031_,
		_w11434_,
		_w12980_
	);
	LUT4 #(
		.INIT('h000d)
	) name12947 (
		_w35_,
		_w11581_,
		_w12979_,
		_w12980_,
		_w12981_
	);
	LUT2 #(
		.INIT('h4)
	) name12948 (
		_w34_,
		_w11434_,
		_w12982_
	);
	LUT3 #(
		.INIT('h8a)
	) name12949 (
		\a[5] ,
		_w34_,
		_w11434_,
		_w12983_
	);
	LUT2 #(
		.INIT('h8)
	) name12950 (
		_w12981_,
		_w12983_,
		_w12984_
	);
	LUT4 #(
		.INIT('h2882)
	) name12951 (
		_w35_,
		_w11233_,
		_w11235_,
		_w11580_,
		_w12985_
	);
	LUT3 #(
		.INIT('h82)
	) name12952 (
		_w6324_,
		_w11233_,
		_w11235_,
		_w12986_
	);
	LUT2 #(
		.INIT('h8)
	) name12953 (
		_w5524_,
		_w11434_,
		_w12987_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12954 (
		_w6031_,
		_w10991_,
		_w11230_,
		_w11232_,
		_w12988_
	);
	LUT2 #(
		.INIT('h1)
	) name12955 (
		_w12987_,
		_w12988_,
		_w12989_
	);
	LUT3 #(
		.INIT('h10)
	) name12956 (
		_w12986_,
		_w12985_,
		_w12989_,
		_w12990_
	);
	LUT3 #(
		.INIT('h80)
	) name12957 (
		_w12637_,
		_w12984_,
		_w12990_,
		_w12991_
	);
	LUT3 #(
		.INIT('h28)
	) name12958 (
		_w35_,
		_w11431_,
		_w11435_,
		_w12992_
	);
	LUT4 #(
		.INIT('h02a8)
	) name12959 (
		_w5524_,
		_w10991_,
		_w11230_,
		_w11232_,
		_w12993_
	);
	LUT4 #(
		.INIT('h007d)
	) name12960 (
		_w6031_,
		_w11233_,
		_w11235_,
		_w12993_,
		_w12994_
	);
	LUT3 #(
		.INIT('h70)
	) name12961 (
		_w6324_,
		_w11427_,
		_w12994_,
		_w12995_
	);
	LUT3 #(
		.INIT('h9a)
	) name12962 (
		\a[5] ,
		_w12992_,
		_w12995_,
		_w12996_
	);
	LUT3 #(
		.INIT('h15)
	) name12963 (
		_w12637_,
		_w12984_,
		_w12990_,
		_w12997_
	);
	LUT3 #(
		.INIT('h6a)
	) name12964 (
		_w12637_,
		_w12984_,
		_w12990_,
		_w12998_
	);
	LUT3 #(
		.INIT('h54)
	) name12965 (
		_w12991_,
		_w12996_,
		_w12997_,
		_w12999_
	);
	LUT4 #(
		.INIT('h009a)
	) name12966 (
		\a[5] ,
		_w12971_,
		_w12975_,
		_w12977_,
		_w13000_
	);
	LUT4 #(
		.INIT('h9a65)
	) name12967 (
		\a[5] ,
		_w12971_,
		_w12975_,
		_w12977_,
		_w13001_
	);
	LUT3 #(
		.INIT('h54)
	) name12968 (
		_w12978_,
		_w12999_,
		_w13000_,
		_w13002_
	);
	LUT4 #(
		.INIT('h009a)
	) name12969 (
		\a[5] ,
		_w12962_,
		_w12967_,
		_w12969_,
		_w13003_
	);
	LUT4 #(
		.INIT('h9a65)
	) name12970 (
		\a[5] ,
		_w12962_,
		_w12967_,
		_w12969_,
		_w13004_
	);
	LUT3 #(
		.INIT('h54)
	) name12971 (
		_w12970_,
		_w13002_,
		_w13003_,
		_w13005_
	);
	LUT2 #(
		.INIT('h2)
	) name12972 (
		_w12959_,
		_w12960_,
		_w13006_
	);
	LUT2 #(
		.INIT('h9)
	) name12973 (
		_w12959_,
		_w12960_,
		_w13007_
	);
	LUT4 #(
		.INIT('h9a65)
	) name12974 (
		\a[5] ,
		_w12949_,
		_w12953_,
		_w12954_,
		_w13008_
	);
	LUT4 #(
		.INIT('h4d00)
	) name12975 (
		_w12959_,
		_w12960_,
		_w13005_,
		_w13008_,
		_w13009_
	);
	LUT4 #(
		.INIT('h9699)
	) name12976 (
		\a[5] ,
		_w12941_,
		_w12942_,
		_w12947_,
		_w13010_
	);
	LUT4 #(
		.INIT('h0155)
	) name12977 (
		_w12948_,
		_w12955_,
		_w13009_,
		_w13010_,
		_w13011_
	);
	LUT2 #(
		.INIT('h4)
	) name12978 (
		_w12935_,
		_w12939_,
		_w13012_
	);
	LUT2 #(
		.INIT('h9)
	) name12979 (
		_w12935_,
		_w12939_,
		_w13013_
	);
	LUT3 #(
		.INIT('h54)
	) name12980 (
		_w12940_,
		_w13011_,
		_w13012_,
		_w13014_
	);
	LUT3 #(
		.INIT('h12)
	) name12981 (
		\a[5] ,
		_w12929_,
		_w12933_,
		_w13015_
	);
	LUT3 #(
		.INIT('h69)
	) name12982 (
		\a[5] ,
		_w12929_,
		_w12933_,
		_w13016_
	);
	LUT3 #(
		.INIT('h54)
	) name12983 (
		_w12934_,
		_w13014_,
		_w13015_,
		_w13017_
	);
	LUT3 #(
		.INIT('h06)
	) name12984 (
		\a[5] ,
		_w12926_,
		_w12927_,
		_w13018_
	);
	LUT3 #(
		.INIT('h69)
	) name12985 (
		\a[5] ,
		_w12926_,
		_w12927_,
		_w13019_
	);
	LUT3 #(
		.INIT('h54)
	) name12986 (
		_w12928_,
		_w13017_,
		_w13018_,
		_w13020_
	);
	LUT3 #(
		.INIT('h06)
	) name12987 (
		\a[5] ,
		_w12920_,
		_w12921_,
		_w13021_
	);
	LUT3 #(
		.INIT('h69)
	) name12988 (
		\a[5] ,
		_w12920_,
		_w12921_,
		_w13022_
	);
	LUT3 #(
		.INIT('h54)
	) name12989 (
		_w12922_,
		_w13020_,
		_w13021_,
		_w13023_
	);
	LUT3 #(
		.INIT('h06)
	) name12990 (
		\a[5] ,
		_w12914_,
		_w12915_,
		_w13024_
	);
	LUT3 #(
		.INIT('h69)
	) name12991 (
		\a[5] ,
		_w12914_,
		_w12915_,
		_w13025_
	);
	LUT3 #(
		.INIT('h54)
	) name12992 (
		_w12916_,
		_w13023_,
		_w13024_,
		_w13026_
	);
	LUT2 #(
		.INIT('h4)
	) name12993 (
		_w12905_,
		_w12909_,
		_w13027_
	);
	LUT2 #(
		.INIT('h9)
	) name12994 (
		_w12905_,
		_w12909_,
		_w13028_
	);
	LUT4 #(
		.INIT('h9699)
	) name12995 (
		\a[5] ,
		_w12898_,
		_w12899_,
		_w12903_,
		_w13029_
	);
	LUT4 #(
		.INIT('h2b00)
	) name12996 (
		_w12905_,
		_w12909_,
		_w13026_,
		_w13029_,
		_w13030_
	);
	LUT4 #(
		.INIT('h9699)
	) name12997 (
		\a[5] ,
		_w12890_,
		_w12891_,
		_w12896_,
		_w13031_
	);
	LUT4 #(
		.INIT('h0155)
	) name12998 (
		_w12897_,
		_w12904_,
		_w13030_,
		_w13031_,
		_w13032_
	);
	LUT2 #(
		.INIT('h2)
	) name12999 (
		_w12887_,
		_w12888_,
		_w13033_
	);
	LUT2 #(
		.INIT('h9)
	) name13000 (
		_w12887_,
		_w12888_,
		_w13034_
	);
	LUT4 #(
		.INIT('h9a65)
	) name13001 (
		\a[5] ,
		_w12877_,
		_w12881_,
		_w12882_,
		_w13035_
	);
	LUT4 #(
		.INIT('h4d00)
	) name13002 (
		_w12887_,
		_w12888_,
		_w13032_,
		_w13035_,
		_w13036_
	);
	LUT4 #(
		.INIT('h9a65)
	) name13003 (
		\a[5] ,
		_w12869_,
		_w12874_,
		_w12875_,
		_w13037_
	);
	LUT4 #(
		.INIT('h0155)
	) name13004 (
		_w12876_,
		_w12883_,
		_w13036_,
		_w13037_,
		_w13038_
	);
	LUT2 #(
		.INIT('h4)
	) name13005 (
		_w12863_,
		_w12867_,
		_w13039_
	);
	LUT2 #(
		.INIT('h9)
	) name13006 (
		_w12863_,
		_w12867_,
		_w13040_
	);
	LUT4 #(
		.INIT('h9699)
	) name13007 (
		\a[5] ,
		_w12856_,
		_w12857_,
		_w12861_,
		_w13041_
	);
	LUT4 #(
		.INIT('h2b00)
	) name13008 (
		_w12863_,
		_w12867_,
		_w13038_,
		_w13041_,
		_w13042_
	);
	LUT4 #(
		.INIT('h9699)
	) name13009 (
		\a[5] ,
		_w12848_,
		_w12849_,
		_w12854_,
		_w13043_
	);
	LUT4 #(
		.INIT('h0155)
	) name13010 (
		_w12855_,
		_w12862_,
		_w13042_,
		_w13043_,
		_w13044_
	);
	LUT2 #(
		.INIT('h2)
	) name13011 (
		_w12845_,
		_w12846_,
		_w13045_
	);
	LUT2 #(
		.INIT('h9)
	) name13012 (
		_w12845_,
		_w12846_,
		_w13046_
	);
	LUT4 #(
		.INIT('h9a65)
	) name13013 (
		\a[5] ,
		_w12835_,
		_w12839_,
		_w12840_,
		_w13047_
	);
	LUT4 #(
		.INIT('h4d00)
	) name13014 (
		_w12845_,
		_w12846_,
		_w13044_,
		_w13047_,
		_w13048_
	);
	LUT4 #(
		.INIT('h9a65)
	) name13015 (
		\a[5] ,
		_w12827_,
		_w12832_,
		_w12833_,
		_w13049_
	);
	LUT4 #(
		.INIT('h0155)
	) name13016 (
		_w12834_,
		_w12841_,
		_w13048_,
		_w13049_,
		_w13050_
	);
	LUT2 #(
		.INIT('h4)
	) name13017 (
		_w12821_,
		_w12825_,
		_w13051_
	);
	LUT2 #(
		.INIT('h9)
	) name13018 (
		_w12821_,
		_w12825_,
		_w13052_
	);
	LUT4 #(
		.INIT('h9699)
	) name13019 (
		\a[5] ,
		_w12814_,
		_w12815_,
		_w12819_,
		_w13053_
	);
	LUT4 #(
		.INIT('h2b00)
	) name13020 (
		_w12821_,
		_w12825_,
		_w13050_,
		_w13053_,
		_w13054_
	);
	LUT4 #(
		.INIT('h9a65)
	) name13021 (
		\a[5] ,
		_w12806_,
		_w12811_,
		_w12812_,
		_w13055_
	);
	LUT4 #(
		.INIT('h0155)
	) name13022 (
		_w12813_,
		_w12820_,
		_w13054_,
		_w13055_,
		_w13056_
	);
	LUT2 #(
		.INIT('h2)
	) name13023 (
		_w12803_,
		_w12804_,
		_w13057_
	);
	LUT2 #(
		.INIT('h9)
	) name13024 (
		_w12803_,
		_w12804_,
		_w13058_
	);
	LUT4 #(
		.INIT('h9a65)
	) name13025 (
		\a[5] ,
		_w11553_,
		_w11557_,
		_w12797_,
		_w13059_
	);
	LUT4 #(
		.INIT('h4d00)
	) name13026 (
		_w12803_,
		_w12804_,
		_w13056_,
		_w13059_,
		_w13060_
	);
	LUT4 #(
		.INIT('h010f)
	) name13027 (
		_w11378_,
		_w11494_,
		_w11551_,
		_w11552_,
		_w13061_
	);
	LUT4 #(
		.INIT('h4445)
	) name13028 (
		_w11547_,
		_w11548_,
		_w11373_,
		_w11375_,
		_w13062_
	);
	LUT3 #(
		.INIT('h28)
	) name13029 (
		_w2975_,
		_w7136_,
		_w7168_,
		_w13063_
	);
	LUT4 #(
		.INIT('h028a)
	) name13030 (
		_w2986_,
		_w7136_,
		_w7166_,
		_w7167_,
		_w13064_
	);
	LUT4 #(
		.INIT('h04c8)
	) name13031 (
		_w2411_,
		_w2874_,
		_w6983_,
		_w6993_,
		_w13065_
	);
	LUT3 #(
		.INIT('h01)
	) name13032 (
		_w13064_,
		_w13065_,
		_w13063_,
		_w13066_
	);
	LUT4 #(
		.INIT('h95aa)
	) name13033 (
		\a[26] ,
		_w2875_,
		_w7696_,
		_w13066_,
		_w13067_
	);
	LUT4 #(
		.INIT('h004d)
	) name13034 (
		_w11503_,
		_w11533_,
		_w11543_,
		_w13067_,
		_w13068_
	);
	LUT4 #(
		.INIT('hb200)
	) name13035 (
		_w11503_,
		_w11533_,
		_w11543_,
		_w13067_,
		_w13069_
	);
	LUT4 #(
		.INIT('h23dc)
	) name13036 (
		_w11534_,
		_w11535_,
		_w11543_,
		_w13067_,
		_w13070_
	);
	LUT3 #(
		.INIT('hb2)
	) name13037 (
		_w11510_,
		_w11525_,
		_w11532_,
		_w13071_
	);
	LUT4 #(
		.INIT('h80fe)
	) name13038 (
		_w7148_,
		_w11352_,
		_w11361_,
		_w11523_,
		_w13072_
	);
	LUT4 #(
		.INIT('h8001)
	) name13039 (
		\a[20] ,
		\a[21] ,
		\a[22] ,
		\a[23] ,
		_w13073_
	);
	LUT4 #(
		.INIT('h559a)
	) name13040 (
		\a[23] ,
		_w7136_,
		_w7166_,
		_w13073_,
		_w13074_
	);
	LUT4 #(
		.INIT('h135f)
	) name13041 (
		_w106_,
		_w55_,
		_w90_,
		_w184_,
		_w13075_
	);
	LUT4 #(
		.INIT('h8000)
	) name13042 (
		_w116_,
		_w710_,
		_w777_,
		_w13075_,
		_w13076_
	);
	LUT4 #(
		.INIT('h8000)
	) name13043 (
		_w1180_,
		_w2365_,
		_w2744_,
		_w4230_,
		_w13077_
	);
	LUT4 #(
		.INIT('h8000)
	) name13044 (
		_w576_,
		_w4166_,
		_w13077_,
		_w13076_,
		_w13078_
	);
	LUT4 #(
		.INIT('h8000)
	) name13045 (
		_w3327_,
		_w7606_,
		_w8370_,
		_w13078_,
		_w13079_
	);
	LUT2 #(
		.INIT('h8)
	) name13046 (
		_w7306_,
		_w13079_,
		_w13080_
	);
	LUT2 #(
		.INIT('h8)
	) name13047 (
		_w11523_,
		_w13080_,
		_w13081_
	);
	LUT2 #(
		.INIT('h1)
	) name13048 (
		_w11523_,
		_w13080_,
		_w13082_
	);
	LUT2 #(
		.INIT('h6)
	) name13049 (
		_w11523_,
		_w13080_,
		_w13083_
	);
	LUT2 #(
		.INIT('h6)
	) name13050 (
		_w13074_,
		_w13083_,
		_w13084_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13051 (
		_w376_,
		_w2983_,
		_w6972_,
		_w6974_,
		_w13085_
	);
	LUT4 #(
		.INIT('h007d)
	) name13052 (
		_w2407_,
		_w2872_,
		_w6975_,
		_w13085_,
		_w13086_
	);
	LUT3 #(
		.INIT('h70)
	) name13053 (
		_w2527_,
		_w7002_,
		_w13086_,
		_w13087_
	);
	LUT3 #(
		.INIT('h70)
	) name13054 (
		_w377_,
		_w7426_,
		_w13087_,
		_w13088_
	);
	LUT3 #(
		.INIT('h96)
	) name13055 (
		_w13072_,
		_w13084_,
		_w13088_,
		_w13089_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13056 (
		_w2549_,
		_w2622_,
		_w6978_,
		_w6980_,
		_w13090_
	);
	LUT4 #(
		.INIT('h007b)
	) name13057 (
		_w2546_,
		_w2617_,
		_w6981_,
		_w13090_,
		_w13091_
	);
	LUT3 #(
		.INIT('h70)
	) name13058 (
		_w2854_,
		_w6996_,
		_w13091_,
		_w13092_
	);
	LUT4 #(
		.INIT('h95aa)
	) name13059 (
		\a[29] ,
		_w2550_,
		_w7500_,
		_w13092_,
		_w13093_
	);
	LUT3 #(
		.INIT('h96)
	) name13060 (
		_w13071_,
		_w13089_,
		_w13093_,
		_w13094_
	);
	LUT2 #(
		.INIT('h6)
	) name13061 (
		_w13070_,
		_w13094_,
		_w13095_
	);
	LUT3 #(
		.INIT('h32)
	) name13062 (
		_w11500_,
		_w11501_,
		_w11544_,
		_w13096_
	);
	LUT4 #(
		.INIT('h7100)
	) name13063 (
		_w11498_,
		_w11499_,
		_w11544_,
		_w13095_,
		_w13097_
	);
	LUT4 #(
		.INIT('h008e)
	) name13064 (
		_w11498_,
		_w11499_,
		_w11544_,
		_w13095_,
		_w13098_
	);
	LUT4 #(
		.INIT('hcd32)
	) name13065 (
		_w11500_,
		_w11501_,
		_w11544_,
		_w13095_,
		_w13099_
	);
	LUT3 #(
		.INIT('h82)
	) name13066 (
		_w11550_,
		_w13062_,
		_w13099_,
		_w13100_
	);
	LUT3 #(
		.INIT('h14)
	) name13067 (
		_w11550_,
		_w13062_,
		_w13099_,
		_w13101_
	);
	LUT3 #(
		.INIT('h69)
	) name13068 (
		_w11550_,
		_w13062_,
		_w13099_,
		_w13102_
	);
	LUT3 #(
		.INIT('h82)
	) name13069 (
		_w35_,
		_w13061_,
		_w13102_,
		_w13103_
	);
	LUT3 #(
		.INIT('h82)
	) name13070 (
		_w6324_,
		_w13062_,
		_w13099_,
		_w13104_
	);
	LUT2 #(
		.INIT('h8)
	) name13071 (
		_w5524_,
		_w11377_,
		_w13105_
	);
	LUT4 #(
		.INIT('h2228)
	) name13072 (
		_w6031_,
		_w11549_,
		_w11373_,
		_w11375_,
		_w13106_
	);
	LUT2 #(
		.INIT('h1)
	) name13073 (
		_w13105_,
		_w13106_,
		_w13107_
	);
	LUT2 #(
		.INIT('h4)
	) name13074 (
		_w13104_,
		_w13107_,
		_w13108_
	);
	LUT3 #(
		.INIT('h82)
	) name13075 (
		_w4459_,
		_w11484_,
		_w11486_,
		_w13109_
	);
	LUT3 #(
		.INIT('h82)
	) name13076 (
		_w4700_,
		_w11280_,
		_w11282_,
		_w13110_
	);
	LUT2 #(
		.INIT('h8)
	) name13077 (
		_w4458_,
		_w11388_,
		_w13111_
	);
	LUT4 #(
		.INIT('h2228)
	) name13078 (
		_w4684_,
		_w7935_,
		_w8077_,
		_w11279_,
		_w13112_
	);
	LUT2 #(
		.INIT('h1)
	) name13079 (
		_w13111_,
		_w13112_,
		_w13113_
	);
	LUT2 #(
		.INIT('h4)
	) name13080 (
		_w13110_,
		_w13113_,
		_w13114_
	);
	LUT3 #(
		.INIT('h82)
	) name13081 (
		_w3710_,
		_w11472_,
		_w11474_,
		_w13115_
	);
	LUT3 #(
		.INIT('h82)
	) name13082 (
		_w3886_,
		_w11268_,
		_w11270_,
		_w13116_
	);
	LUT2 #(
		.INIT('h8)
	) name13083 (
		_w3709_,
		_w11400_,
		_w13117_
	);
	LUT4 #(
		.INIT('h2228)
	) name13084 (
		_w3877_,
		_w8794_,
		_w8994_,
		_w11267_,
		_w13118_
	);
	LUT2 #(
		.INIT('h1)
	) name13085 (
		_w13117_,
		_w13118_,
		_w13119_
	);
	LUT2 #(
		.INIT('h4)
	) name13086 (
		_w13116_,
		_w13119_,
		_w13120_
	);
	LUT3 #(
		.INIT('h32)
	) name13087 (
		_w12718_,
		_w12759_,
		_w12760_,
		_w13121_
	);
	LUT3 #(
		.INIT('h82)
	) name13088 (
		_w3214_,
		_w10580_,
		_w11254_,
		_w13122_
	);
	LUT4 #(
		.INIT('h007d)
	) name13089 (
		_w3249_,
		_w10268_,
		_w11255_,
		_w13122_,
		_w13123_
	);
	LUT4 #(
		.INIT('h7d00)
	) name13090 (
		_w3262_,
		_w11256_,
		_w11258_,
		_w13123_,
		_w13124_
	);
	LUT4 #(
		.INIT('h7d00)
	) name13091 (
		_w37_,
		_w11459_,
		_w11461_,
		_w13124_,
		_w13125_
	);
	LUT3 #(
		.INIT('h32)
	) name13092 (
		_w12723_,
		_w12755_,
		_w12756_,
		_w13126_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13093 (
		_w2550_,
		_w11423_,
		_w11443_,
		_w11444_,
		_w13127_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13094 (
		_w2854_,
		_w10945_,
		_w11246_,
		_w11248_,
		_w13128_
	);
	LUT3 #(
		.INIT('h82)
	) name13095 (
		_w2549_,
		_w11241_,
		_w11243_,
		_w13129_
	);
	LUT3 #(
		.INIT('h07)
	) name13096 (
		_w2617_,
		_w11421_,
		_w13129_,
		_w13130_
	);
	LUT2 #(
		.INIT('h4)
	) name13097 (
		_w13128_,
		_w13130_,
		_w13131_
	);
	LUT3 #(
		.INIT('h32)
	) name13098 (
		_w12729_,
		_w12743_,
		_w12744_,
		_w13132_
	);
	LUT3 #(
		.INIT('h40)
	) name13099 (
		_w324_,
		_w752_,
		_w1235_,
		_w13133_
	);
	LUT4 #(
		.INIT('h1000)
	) name13100 (
		_w227_,
		_w462_,
		_w1635_,
		_w3791_,
		_w13134_
	);
	LUT3 #(
		.INIT('h1f)
	) name13101 (
		_w59_,
		_w67_,
		_w378_,
		_w13135_
	);
	LUT3 #(
		.INIT('h1f)
	) name13102 (
		_w110_,
		_w46_,
		_w259_,
		_w13136_
	);
	LUT4 #(
		.INIT('h4000)
	) name13103 (
		_w426_,
		_w7516_,
		_w13136_,
		_w13135_,
		_w13137_
	);
	LUT4 #(
		.INIT('h8000)
	) name13104 (
		_w7213_,
		_w13137_,
		_w13133_,
		_w13134_,
		_w13138_
	);
	LUT3 #(
		.INIT('h80)
	) name13105 (
		_w7190_,
		_w11515_,
		_w13138_,
		_w13139_
	);
	LUT2 #(
		.INIT('h8)
	) name13106 (
		_w8291_,
		_w13139_,
		_w13140_
	);
	LUT3 #(
		.INIT('h82)
	) name13107 (
		_w377_,
		_w11436_,
		_w11438_,
		_w13141_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13108 (
		_w2527_,
		_w10968_,
		_w11238_,
		_w11240_,
		_w13142_
	);
	LUT3 #(
		.INIT('h82)
	) name13109 (
		_w376_,
		_w11233_,
		_w11235_,
		_w13143_
	);
	LUT3 #(
		.INIT('h07)
	) name13110 (
		_w2407_,
		_w11427_,
		_w13143_,
		_w13144_
	);
	LUT2 #(
		.INIT('h4)
	) name13111 (
		_w13142_,
		_w13144_,
		_w13145_
	);
	LUT3 #(
		.INIT('h45)
	) name13112 (
		_w13140_,
		_w13141_,
		_w13145_,
		_w13146_
	);
	LUT3 #(
		.INIT('h20)
	) name13113 (
		_w13140_,
		_w13141_,
		_w13145_,
		_w13147_
	);
	LUT3 #(
		.INIT('h9a)
	) name13114 (
		_w13140_,
		_w13141_,
		_w13145_,
		_w13148_
	);
	LUT2 #(
		.INIT('h9)
	) name13115 (
		_w13132_,
		_w13148_,
		_w13149_
	);
	LUT4 #(
		.INIT('h6500)
	) name13116 (
		\a[29] ,
		_w13127_,
		_w13131_,
		_w13149_,
		_w13150_
	);
	LUT4 #(
		.INIT('h9a65)
	) name13117 (
		\a[29] ,
		_w13127_,
		_w13131_,
		_w13149_,
		_w13151_
	);
	LUT4 #(
		.INIT('h7100)
	) name13118 (
		_w12724_,
		_w12728_,
		_w12746_,
		_w13151_,
		_w13152_
	);
	LUT4 #(
		.INIT('h32cd)
	) name13119 (
		_w12724_,
		_w12747_,
		_w12748_,
		_w13151_,
		_w13153_
	);
	LUT3 #(
		.INIT('h82)
	) name13120 (
		_w2874_,
		_w11249_,
		_w11251_,
		_w13154_
	);
	LUT3 #(
		.INIT('h07)
	) name13121 (
		_w2975_,
		_w11415_,
		_w13154_,
		_w13155_
	);
	LUT4 #(
		.INIT('h7d00)
	) name13122 (
		_w2986_,
		_w10599_,
		_w11253_,
		_w13155_,
		_w13156_
	);
	LUT4 #(
		.INIT('h7d00)
	) name13123 (
		_w2875_,
		_w11450_,
		_w11452_,
		_w13156_,
		_w13157_
	);
	LUT3 #(
		.INIT('h84)
	) name13124 (
		\a[26] ,
		_w13153_,
		_w13157_,
		_w13158_
	);
	LUT3 #(
		.INIT('h12)
	) name13125 (
		\a[26] ,
		_w13153_,
		_w13157_,
		_w13159_
	);
	LUT3 #(
		.INIT('h69)
	) name13126 (
		\a[26] ,
		_w13153_,
		_w13157_,
		_w13160_
	);
	LUT2 #(
		.INIT('h9)
	) name13127 (
		_w13126_,
		_w13160_,
		_w13161_
	);
	LUT3 #(
		.INIT('h90)
	) name13128 (
		\a[23] ,
		_w13125_,
		_w13161_,
		_w13162_
	);
	LUT3 #(
		.INIT('h06)
	) name13129 (
		\a[23] ,
		_w13125_,
		_w13161_,
		_w13163_
	);
	LUT3 #(
		.INIT('h69)
	) name13130 (
		\a[23] ,
		_w13125_,
		_w13161_,
		_w13164_
	);
	LUT2 #(
		.INIT('h9)
	) name13131 (
		_w13121_,
		_w13164_,
		_w13165_
	);
	LUT3 #(
		.INIT('h82)
	) name13132 (
		_w3312_,
		_w11465_,
		_w11467_,
		_w13166_
	);
	LUT3 #(
		.INIT('h82)
	) name13133 (
		_w3654_,
		_w11262_,
		_w11264_,
		_w13167_
	);
	LUT2 #(
		.INIT('h8)
	) name13134 (
		_w3311_,
		_w11406_,
		_w13168_
	);
	LUT4 #(
		.INIT('h2228)
	) name13135 (
		_w3645_,
		_w9446_,
		_w9702_,
		_w11261_,
		_w13169_
	);
	LUT2 #(
		.INIT('h1)
	) name13136 (
		_w13168_,
		_w13169_,
		_w13170_
	);
	LUT2 #(
		.INIT('h4)
	) name13137 (
		_w13167_,
		_w13170_,
		_w13171_
	);
	LUT4 #(
		.INIT('h4844)
	) name13138 (
		\a[20] ,
		_w13165_,
		_w13166_,
		_w13171_,
		_w13172_
	);
	LUT4 #(
		.INIT('h9699)
	) name13139 (
		\a[20] ,
		_w13165_,
		_w13166_,
		_w13171_,
		_w13173_
	);
	LUT3 #(
		.INIT('h1e)
	) name13140 (
		_w12768_,
		_w12770_,
		_w13173_,
		_w13174_
	);
	LUT4 #(
		.INIT('h6500)
	) name13141 (
		\a[17] ,
		_w13115_,
		_w13120_,
		_w13174_,
		_w13175_
	);
	LUT4 #(
		.INIT('h9a65)
	) name13142 (
		\a[17] ,
		_w13115_,
		_w13120_,
		_w13174_,
		_w13176_
	);
	LUT3 #(
		.INIT('h1e)
	) name13143 (
		_w12772_,
		_w12774_,
		_w13176_,
		_w13177_
	);
	LUT3 #(
		.INIT('h82)
	) name13144 (
		_w4034_,
		_w11478_,
		_w11480_,
		_w13178_
	);
	LUT3 #(
		.INIT('h82)
	) name13145 (
		_w4382_,
		_w11274_,
		_w11276_,
		_w13179_
	);
	LUT2 #(
		.INIT('h8)
	) name13146 (
		_w4033_,
		_w11394_,
		_w13180_
	);
	LUT4 #(
		.INIT('h2228)
	) name13147 (
		_w4367_,
		_w8466_,
		_w8541_,
		_w11273_,
		_w13181_
	);
	LUT2 #(
		.INIT('h1)
	) name13148 (
		_w13180_,
		_w13181_,
		_w13182_
	);
	LUT2 #(
		.INIT('h4)
	) name13149 (
		_w13179_,
		_w13182_,
		_w13183_
	);
	LUT4 #(
		.INIT('h4844)
	) name13150 (
		\a[14] ,
		_w13177_,
		_w13178_,
		_w13183_,
		_w13184_
	);
	LUT4 #(
		.INIT('h9699)
	) name13151 (
		\a[14] ,
		_w13177_,
		_w13178_,
		_w13183_,
		_w13185_
	);
	LUT3 #(
		.INIT('h1e)
	) name13152 (
		_w12781_,
		_w12783_,
		_w13185_,
		_w13186_
	);
	LUT4 #(
		.INIT('h6500)
	) name13153 (
		\a[11] ,
		_w13109_,
		_w13114_,
		_w13186_,
		_w13187_
	);
	LUT4 #(
		.INIT('h9a65)
	) name13154 (
		\a[11] ,
		_w13109_,
		_w13114_,
		_w13186_,
		_w13188_
	);
	LUT3 #(
		.INIT('h1e)
	) name13155 (
		_w12785_,
		_w12787_,
		_w13188_,
		_w13189_
	);
	LUT3 #(
		.INIT('h82)
	) name13156 (
		_w4876_,
		_w11490_,
		_w11492_,
		_w13190_
	);
	LUT3 #(
		.INIT('h82)
	) name13157 (
		_w5286_,
		_w11286_,
		_w11335_,
		_w13191_
	);
	LUT2 #(
		.INIT('h8)
	) name13158 (
		_w4875_,
		_w11382_,
		_w13192_
	);
	LUT4 #(
		.INIT('h2228)
	) name13159 (
		_w5271_,
		_w7695_,
		_w7750_,
		_w11285_,
		_w13193_
	);
	LUT2 #(
		.INIT('h1)
	) name13160 (
		_w13192_,
		_w13193_,
		_w13194_
	);
	LUT2 #(
		.INIT('h4)
	) name13161 (
		_w13191_,
		_w13194_,
		_w13195_
	);
	LUT4 #(
		.INIT('h4844)
	) name13162 (
		\a[8] ,
		_w13189_,
		_w13190_,
		_w13195_,
		_w13196_
	);
	LUT4 #(
		.INIT('h9699)
	) name13163 (
		\a[8] ,
		_w13189_,
		_w13190_,
		_w13195_,
		_w13197_
	);
	LUT3 #(
		.INIT('h1e)
	) name13164 (
		_w12794_,
		_w12796_,
		_w13197_,
		_w13198_
	);
	LUT4 #(
		.INIT('h6500)
	) name13165 (
		\a[5] ,
		_w13103_,
		_w13108_,
		_w13198_,
		_w13199_
	);
	LUT4 #(
		.INIT('h9a65)
	) name13166 (
		\a[5] ,
		_w13103_,
		_w13108_,
		_w13198_,
		_w13200_
	);
	LUT3 #(
		.INIT('h1e)
	) name13167 (
		_w12798_,
		_w13060_,
		_w13200_,
		_w13201_
	);
	LUT3 #(
		.INIT('h45)
	) name13168 (
		_w13068_,
		_w13069_,
		_w13094_,
		_w13202_
	);
	LUT4 #(
		.INIT('h0a02)
	) name13169 (
		_w2875_,
		_w7169_,
		_w7419_,
		_w7686_,
		_w13203_
	);
	LUT3 #(
		.INIT('h28)
	) name13170 (
		_w2874_,
		_w7136_,
		_w7168_,
		_w13204_
	);
	LUT4 #(
		.INIT('h87e1)
	) name13171 (
		\a[23] ,
		\a[24] ,
		\a[25] ,
		\a[26] ,
		_w13205_
	);
	LUT3 #(
		.INIT('h0b)
	) name13172 (
		_w7136_,
		_w7166_,
		_w13205_,
		_w13206_
	);
	LUT3 #(
		.INIT('h40)
	) name13173 (
		_w2986_,
		_w7136_,
		_w7167_,
		_w13207_
	);
	LUT3 #(
		.INIT('h31)
	) name13174 (
		_w13206_,
		_w13204_,
		_w13207_,
		_w13208_
	);
	LUT3 #(
		.INIT('h9a)
	) name13175 (
		\a[26] ,
		_w13203_,
		_w13208_,
		_w13209_
	);
	LUT3 #(
		.INIT('h0d)
	) name13176 (
		_w13074_,
		_w13081_,
		_w13082_,
		_w13210_
	);
	LUT4 #(
		.INIT('h135f)
	) name13177 (
		_w122_,
		_w110_,
		_w41_,
		_w176_,
		_w13211_
	);
	LUT3 #(
		.INIT('h80)
	) name13178 (
		_w503_,
		_w1180_,
		_w13211_,
		_w13212_
	);
	LUT4 #(
		.INIT('h8000)
	) name13179 (
		_w521_,
		_w522_,
		_w720_,
		_w4282_,
		_w13213_
	);
	LUT2 #(
		.INIT('h8)
	) name13180 (
		_w13212_,
		_w13213_,
		_w13214_
	);
	LUT2 #(
		.INIT('h2)
	) name13181 (
		_w287_,
		_w462_,
		_w13215_
	);
	LUT4 #(
		.INIT('h8000)
	) name13182 (
		_w804_,
		_w816_,
		_w1402_,
		_w1982_,
		_w13216_
	);
	LUT3 #(
		.INIT('h80)
	) name13183 (
		_w622_,
		_w13215_,
		_w13216_,
		_w13217_
	);
	LUT4 #(
		.INIT('h8000)
	) name13184 (
		_w175_,
		_w178_,
		_w13214_,
		_w13217_,
		_w13218_
	);
	LUT2 #(
		.INIT('h8)
	) name13185 (
		_w666_,
		_w13218_,
		_w13219_
	);
	LUT4 #(
		.INIT('h4d00)
	) name13186 (
		_w11523_,
		_w13074_,
		_w13080_,
		_w13219_,
		_w13220_
	);
	LUT4 #(
		.INIT('h00b2)
	) name13187 (
		_w11523_,
		_w13074_,
		_w13080_,
		_w13219_,
		_w13221_
	);
	LUT4 #(
		.INIT('h0df2)
	) name13188 (
		_w13074_,
		_w13081_,
		_w13082_,
		_w13219_,
		_w13222_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13189 (
		_w377_,
		_w7004_,
		_w7127_,
		_w7128_,
		_w13223_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13190 (
		_w2527_,
		_w2622_,
		_w6978_,
		_w6980_,
		_w13224_
	);
	LUT3 #(
		.INIT('h82)
	) name13191 (
		_w376_,
		_w2872_,
		_w6975_,
		_w13225_
	);
	LUT3 #(
		.INIT('h07)
	) name13192 (
		_w2407_,
		_w7002_,
		_w13225_,
		_w13226_
	);
	LUT2 #(
		.INIT('h4)
	) name13193 (
		_w13224_,
		_w13226_,
		_w13227_
	);
	LUT2 #(
		.INIT('h4)
	) name13194 (
		_w13223_,
		_w13227_,
		_w13228_
	);
	LUT2 #(
		.INIT('h9)
	) name13195 (
		_w13222_,
		_w13228_,
		_w13229_
	);
	LUT3 #(
		.INIT('h4d)
	) name13196 (
		_w13072_,
		_w13084_,
		_w13088_,
		_w13230_
	);
	LUT4 #(
		.INIT('h4d00)
	) name13197 (
		_w13072_,
		_w13084_,
		_w13088_,
		_w13229_,
		_w13231_
	);
	LUT4 #(
		.INIT('h00b2)
	) name13198 (
		_w13072_,
		_w13084_,
		_w13088_,
		_w13229_,
		_w13232_
	);
	LUT4 #(
		.INIT('hb24d)
	) name13199 (
		_w13072_,
		_w13084_,
		_w13088_,
		_w13229_,
		_w13233_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13200 (
		_w2550_,
		_w6998_,
		_w7133_,
		_w7134_,
		_w13234_
	);
	LUT4 #(
		.INIT('h04c8)
	) name13201 (
		_w2411_,
		_w2854_,
		_w6983_,
		_w6993_,
		_w13235_
	);
	LUT3 #(
		.INIT('h84)
	) name13202 (
		_w2546_,
		_w2549_,
		_w6981_,
		_w13236_
	);
	LUT3 #(
		.INIT('h07)
	) name13203 (
		_w2617_,
		_w6996_,
		_w13236_,
		_w13237_
	);
	LUT2 #(
		.INIT('h4)
	) name13204 (
		_w13235_,
		_w13237_,
		_w13238_
	);
	LUT3 #(
		.INIT('h9a)
	) name13205 (
		\a[29] ,
		_w13234_,
		_w13238_,
		_w13239_
	);
	LUT2 #(
		.INIT('h9)
	) name13206 (
		_w13233_,
		_w13239_,
		_w13240_
	);
	LUT3 #(
		.INIT('h4d)
	) name13207 (
		_w13071_,
		_w13089_,
		_w13093_,
		_w13241_
	);
	LUT3 #(
		.INIT('h69)
	) name13208 (
		_w13240_,
		_w13241_,
		_w13209_,
		_w13242_
	);
	LUT2 #(
		.INIT('h4)
	) name13209 (
		_w13202_,
		_w13242_,
		_w13243_
	);
	LUT2 #(
		.INIT('h9)
	) name13210 (
		_w13202_,
		_w13242_,
		_w13244_
	);
	LUT4 #(
		.INIT('hd400)
	) name13211 (
		_w13062_,
		_w13095_,
		_w13096_,
		_w13244_,
		_w13245_
	);
	LUT4 #(
		.INIT('h002b)
	) name13212 (
		_w13062_,
		_w13095_,
		_w13096_,
		_w13244_,
		_w13246_
	);
	LUT4 #(
		.INIT('h32cd)
	) name13213 (
		_w13062_,
		_w13097_,
		_w13098_,
		_w13244_,
		_w13247_
	);
	LUT4 #(
		.INIT('h135f)
	) name13214 (
		_w122_,
		_w55_,
		_w50_,
		_w259_,
		_w13248_
	);
	LUT4 #(
		.INIT('h8000)
	) name13215 (
		_w260_,
		_w3796_,
		_w7993_,
		_w13248_,
		_w13249_
	);
	LUT4 #(
		.INIT('h2000)
	) name13216 (
		_w116_,
		_w273_,
		_w348_,
		_w995_,
		_w13250_
	);
	LUT3 #(
		.INIT('h80)
	) name13217 (
		_w532_,
		_w13249_,
		_w13250_,
		_w13251_
	);
	LUT4 #(
		.INIT('h8000)
	) name13218 (
		_w175_,
		_w178_,
		_w505_,
		_w13251_,
		_w13252_
	);
	LUT3 #(
		.INIT('h80)
	) name13219 (
		_w587_,
		_w608_,
		_w13252_,
		_w13253_
	);
	LUT2 #(
		.INIT('h4)
	) name13220 (
		_w13219_,
		_w13253_,
		_w13254_
	);
	LUT2 #(
		.INIT('h2)
	) name13221 (
		_w13219_,
		_w13253_,
		_w13255_
	);
	LUT2 #(
		.INIT('h9)
	) name13222 (
		_w13219_,
		_w13253_,
		_w13256_
	);
	LUT3 #(
		.INIT('h82)
	) name13223 (
		_w377_,
		_w7129_,
		_w7131_,
		_w13257_
	);
	LUT3 #(
		.INIT('h82)
	) name13224 (
		_w2527_,
		_w2546_,
		_w6981_,
		_w13258_
	);
	LUT2 #(
		.INIT('h8)
	) name13225 (
		_w376_,
		_w7002_,
		_w13259_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13226 (
		_w2407_,
		_w2622_,
		_w6978_,
		_w6980_,
		_w13260_
	);
	LUT2 #(
		.INIT('h1)
	) name13227 (
		_w13259_,
		_w13260_,
		_w13261_
	);
	LUT2 #(
		.INIT('h4)
	) name13228 (
		_w13258_,
		_w13261_,
		_w13262_
	);
	LUT3 #(
		.INIT('h65)
	) name13229 (
		_w13256_,
		_w13257_,
		_w13262_,
		_w13263_
	);
	LUT4 #(
		.INIT('h4d00)
	) name13230 (
		_w13210_,
		_w13219_,
		_w13228_,
		_w13263_,
		_w13264_
	);
	LUT4 #(
		.INIT('h54ab)
	) name13231 (
		_w13220_,
		_w13221_,
		_w13228_,
		_w13263_,
		_w13265_
	);
	LUT4 #(
		.INIT('h80a8)
	) name13232 (
		_w13265_,
		_w13229_,
		_w13230_,
		_w13239_,
		_w13266_
	);
	LUT4 #(
		.INIT('h6665)
	) name13233 (
		_w13265_,
		_w13231_,
		_w13232_,
		_w13239_,
		_w13267_
	);
	LUT4 #(
		.INIT('h028a)
	) name13234 (
		_w2874_,
		_w7136_,
		_w7166_,
		_w7167_,
		_w13268_
	);
	LUT2 #(
		.INIT('h1)
	) name13235 (
		_w13268_,
		_w13206_,
		_w13269_
	);
	LUT4 #(
		.INIT('h5700)
	) name13236 (
		_w2875_,
		_w7418_,
		_w7419_,
		_w13269_,
		_w13270_
	);
	LUT3 #(
		.INIT('h82)
	) name13237 (
		_w2550_,
		_w7135_,
		_w7172_,
		_w13271_
	);
	LUT3 #(
		.INIT('h28)
	) name13238 (
		_w2854_,
		_w7136_,
		_w7168_,
		_w13272_
	);
	LUT2 #(
		.INIT('h8)
	) name13239 (
		_w2549_,
		_w6996_,
		_w13273_
	);
	LUT4 #(
		.INIT('h04c8)
	) name13240 (
		_w2411_,
		_w2617_,
		_w6983_,
		_w6993_,
		_w13274_
	);
	LUT2 #(
		.INIT('h1)
	) name13241 (
		_w13273_,
		_w13274_,
		_w13275_
	);
	LUT2 #(
		.INIT('h4)
	) name13242 (
		_w13272_,
		_w13275_,
		_w13276_
	);
	LUT3 #(
		.INIT('h9a)
	) name13243 (
		\a[29] ,
		_w13271_,
		_w13276_,
		_w13277_
	);
	LUT3 #(
		.INIT('h09)
	) name13244 (
		\a[26] ,
		_w13270_,
		_w13277_,
		_w13278_
	);
	LUT3 #(
		.INIT('h60)
	) name13245 (
		\a[26] ,
		_w13270_,
		_w13277_,
		_w13279_
	);
	LUT3 #(
		.INIT('h96)
	) name13246 (
		\a[26] ,
		_w13270_,
		_w13277_,
		_w13280_
	);
	LUT2 #(
		.INIT('h6)
	) name13247 (
		_w13267_,
		_w13280_,
		_w13281_
	);
	LUT3 #(
		.INIT('h8e)
	) name13248 (
		_w13240_,
		_w13241_,
		_w13209_,
		_w13282_
	);
	LUT2 #(
		.INIT('h8)
	) name13249 (
		_w13281_,
		_w13282_,
		_w13283_
	);
	LUT2 #(
		.INIT('h1)
	) name13250 (
		_w13281_,
		_w13282_,
		_w13284_
	);
	LUT2 #(
		.INIT('h6)
	) name13251 (
		_w13281_,
		_w13282_,
		_w13285_
	);
	LUT3 #(
		.INIT('h1e)
	) name13252 (
		_w13243_,
		_w13245_,
		_w13285_,
		_w13286_
	);
	LUT4 #(
		.INIT('h1e00)
	) name13253 (
		_w13243_,
		_w13245_,
		_w13285_,
		_w13247_,
		_w13287_
	);
	LUT4 #(
		.INIT('h2940)
	) name13254 (
		_w13062_,
		_w13095_,
		_w13096_,
		_w13244_,
		_w13288_
	);
	LUT4 #(
		.INIT('h8679)
	) name13255 (
		_w13062_,
		_w13097_,
		_w13099_,
		_w13244_,
		_w13289_
	);
	LUT4 #(
		.INIT('hdc00)
	) name13256 (
		_w13061_,
		_w13100_,
		_w13102_,
		_w13289_,
		_w13290_
	);
	LUT4 #(
		.INIT('h1e2d)
	) name13257 (
		_w13243_,
		_w13245_,
		_w13285_,
		_w13246_,
		_w13291_
	);
	LUT4 #(
		.INIT('h0155)
	) name13258 (
		_w13287_,
		_w13288_,
		_w13290_,
		_w13291_,
		_w13292_
	);
	LUT4 #(
		.INIT('h5501)
	) name13259 (
		_w13283_,
		_w13243_,
		_w13245_,
		_w13284_,
		_w13293_
	);
	LUT3 #(
		.INIT('h28)
	) name13260 (
		_w2617_,
		_w7136_,
		_w7168_,
		_w13294_
	);
	LUT4 #(
		.INIT('h028a)
	) name13261 (
		_w2854_,
		_w7136_,
		_w7166_,
		_w7167_,
		_w13295_
	);
	LUT4 #(
		.INIT('h04c8)
	) name13262 (
		_w2411_,
		_w2549_,
		_w6983_,
		_w6993_,
		_w13296_
	);
	LUT3 #(
		.INIT('h01)
	) name13263 (
		_w13295_,
		_w13296_,
		_w13294_,
		_w13297_
	);
	LUT4 #(
		.INIT('h95aa)
	) name13264 (
		\a[29] ,
		_w2550_,
		_w7696_,
		_w13297_,
		_w13298_
	);
	LUT4 #(
		.INIT('h2322)
	) name13265 (
		_w13254_,
		_w13255_,
		_w13257_,
		_w13262_,
		_w13299_
	);
	LUT4 #(
		.INIT('h8001)
	) name13266 (
		\a[23] ,
		\a[24] ,
		\a[25] ,
		\a[26] ,
		_w13300_
	);
	LUT4 #(
		.INIT('h559a)
	) name13267 (
		\a[26] ,
		_w7136_,
		_w7166_,
		_w13300_,
		_w13301_
	);
	LUT3 #(
		.INIT('h80)
	) name13268 (
		_w341_,
		_w416_,
		_w417_,
		_w13302_
	);
	LUT4 #(
		.INIT('h0777)
	) name13269 (
		_w78_,
		_w56_,
		_w65_,
		_w419_,
		_w13303_
	);
	LUT2 #(
		.INIT('h8)
	) name13270 (
		_w553_,
		_w13303_,
		_w13304_
	);
	LUT3 #(
		.INIT('h80)
	) name13271 (
		_w100_,
		_w499_,
		_w13304_,
		_w13305_
	);
	LUT3 #(
		.INIT('h80)
	) name13272 (
		_w257_,
		_w13302_,
		_w13305_,
		_w13306_
	);
	LUT2 #(
		.INIT('h8)
	) name13273 (
		_w13219_,
		_w13306_,
		_w13307_
	);
	LUT2 #(
		.INIT('h1)
	) name13274 (
		_w13219_,
		_w13306_,
		_w13308_
	);
	LUT2 #(
		.INIT('h6)
	) name13275 (
		_w13219_,
		_w13306_,
		_w13309_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13276 (
		_w376_,
		_w2622_,
		_w6978_,
		_w6980_,
		_w13310_
	);
	LUT4 #(
		.INIT('h007d)
	) name13277 (
		_w2407_,
		_w2546_,
		_w6981_,
		_w13310_,
		_w13311_
	);
	LUT3 #(
		.INIT('h70)
	) name13278 (
		_w2527_,
		_w6996_,
		_w13311_,
		_w13312_
	);
	LUT3 #(
		.INIT('h70)
	) name13279 (
		_w377_,
		_w7500_,
		_w13312_,
		_w13313_
	);
	LUT4 #(
		.INIT('h6996)
	) name13280 (
		_w13299_,
		_w13301_,
		_w13309_,
		_w13313_,
		_w13314_
	);
	LUT2 #(
		.INIT('h4)
	) name13281 (
		_w13298_,
		_w13314_,
		_w13315_
	);
	LUT2 #(
		.INIT('h2)
	) name13282 (
		_w13298_,
		_w13314_,
		_w13316_
	);
	LUT2 #(
		.INIT('h9)
	) name13283 (
		_w13298_,
		_w13314_,
		_w13317_
	);
	LUT3 #(
		.INIT('h1e)
	) name13284 (
		_w13264_,
		_w13266_,
		_w13317_,
		_w13318_
	);
	LUT3 #(
		.INIT('h31)
	) name13285 (
		_w13267_,
		_w13278_,
		_w13279_,
		_w13319_
	);
	LUT2 #(
		.INIT('h2)
	) name13286 (
		_w13318_,
		_w13319_,
		_w13320_
	);
	LUT2 #(
		.INIT('h4)
	) name13287 (
		_w13318_,
		_w13319_,
		_w13321_
	);
	LUT2 #(
		.INIT('h9)
	) name13288 (
		_w13318_,
		_w13319_,
		_w13322_
	);
	LUT3 #(
		.INIT('h90)
	) name13289 (
		_w13293_,
		_w13322_,
		_w13286_,
		_w13323_
	);
	LUT3 #(
		.INIT('h06)
	) name13290 (
		_w13293_,
		_w13322_,
		_w13286_,
		_w13324_
	);
	LUT3 #(
		.INIT('h69)
	) name13291 (
		_w13293_,
		_w13322_,
		_w13286_,
		_w13325_
	);
	LUT3 #(
		.INIT('h82)
	) name13292 (
		_w6335_,
		_w13292_,
		_w13325_,
		_w13326_
	);
	LUT3 #(
		.INIT('h82)
	) name13293 (
		_w6657_,
		_w13293_,
		_w13322_,
		_w13327_
	);
	LUT2 #(
		.INIT('h8)
	) name13294 (
		_w6334_,
		_w13247_,
		_w13328_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13295 (
		_w6650_,
		_w13243_,
		_w13245_,
		_w13285_,
		_w13329_
	);
	LUT2 #(
		.INIT('h1)
	) name13296 (
		_w13328_,
		_w13329_,
		_w13330_
	);
	LUT2 #(
		.INIT('h4)
	) name13297 (
		_w13327_,
		_w13330_,
		_w13331_
	);
	LUT3 #(
		.INIT('h9a)
	) name13298 (
		\a[2] ,
		_w13326_,
		_w13331_,
		_w13332_
	);
	LUT4 #(
		.INIT('h4844)
	) name13299 (
		\a[2] ,
		_w13201_,
		_w13326_,
		_w13331_,
		_w13333_
	);
	LUT4 #(
		.INIT('h9699)
	) name13300 (
		\a[2] ,
		_w13201_,
		_w13326_,
		_w13331_,
		_w13334_
	);
	LUT4 #(
		.INIT('h54ab)
	) name13301 (
		_w12805_,
		_w13056_,
		_w13057_,
		_w13059_,
		_w13335_
	);
	LUT2 #(
		.INIT('h9)
	) name13302 (
		_w13056_,
		_w13058_,
		_w13336_
	);
	LUT3 #(
		.INIT('h82)
	) name13303 (
		_w6335_,
		_w13061_,
		_w13102_,
		_w13337_
	);
	LUT3 #(
		.INIT('h82)
	) name13304 (
		_w6657_,
		_w13062_,
		_w13099_,
		_w13338_
	);
	LUT2 #(
		.INIT('h8)
	) name13305 (
		_w6334_,
		_w11377_,
		_w13339_
	);
	LUT4 #(
		.INIT('h2228)
	) name13306 (
		_w6650_,
		_w11549_,
		_w11373_,
		_w11375_,
		_w13340_
	);
	LUT2 #(
		.INIT('h1)
	) name13307 (
		_w13339_,
		_w13340_,
		_w13341_
	);
	LUT2 #(
		.INIT('h4)
	) name13308 (
		_w13338_,
		_w13341_,
		_w13342_
	);
	LUT3 #(
		.INIT('h1e)
	) name13309 (
		_w12820_,
		_w13054_,
		_w13055_,
		_w13343_
	);
	LUT4 #(
		.INIT('h009a)
	) name13310 (
		\a[2] ,
		_w13337_,
		_w13342_,
		_w13343_,
		_w13344_
	);
	LUT4 #(
		.INIT('h6500)
	) name13311 (
		\a[2] ,
		_w13337_,
		_w13342_,
		_w13343_,
		_w13345_
	);
	LUT4 #(
		.INIT('h54ab)
	) name13312 (
		_w12826_,
		_w13050_,
		_w13051_,
		_w13053_,
		_w13346_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13313 (
		_w6335_,
		_w11378_,
		_w11494_,
		_w11552_,
		_w13347_
	);
	LUT4 #(
		.INIT('h2228)
	) name13314 (
		_w6657_,
		_w11549_,
		_w11373_,
		_w11375_,
		_w13348_
	);
	LUT3 #(
		.INIT('h82)
	) name13315 (
		_w6334_,
		_w11286_,
		_w11335_,
		_w13349_
	);
	LUT3 #(
		.INIT('h07)
	) name13316 (
		_w6650_,
		_w11377_,
		_w13349_,
		_w13350_
	);
	LUT2 #(
		.INIT('h4)
	) name13317 (
		_w13348_,
		_w13350_,
		_w13351_
	);
	LUT4 #(
		.INIT('h2122)
	) name13318 (
		\a[2] ,
		_w13346_,
		_w13347_,
		_w13351_,
		_w13352_
	);
	LUT4 #(
		.INIT('h4844)
	) name13319 (
		\a[2] ,
		_w13346_,
		_w13347_,
		_w13351_,
		_w13353_
	);
	LUT2 #(
		.INIT('h9)
	) name13320 (
		_w13050_,
		_w13052_,
		_w13354_
	);
	LUT4 #(
		.INIT('h2228)
	) name13321 (
		_w6334_,
		_w7695_,
		_w7750_,
		_w11285_,
		_w13355_
	);
	LUT4 #(
		.INIT('h007d)
	) name13322 (
		_w6650_,
		_w11286_,
		_w11335_,
		_w13355_,
		_w13356_
	);
	LUT3 #(
		.INIT('h70)
	) name13323 (
		_w6657_,
		_w11377_,
		_w13356_,
		_w13357_
	);
	LUT4 #(
		.INIT('h6a55)
	) name13324 (
		\a[2] ,
		_w6335_,
		_w12799_,
		_w13357_,
		_w13358_
	);
	LUT3 #(
		.INIT('h82)
	) name13325 (
		_w6335_,
		_w11490_,
		_w11492_,
		_w13359_
	);
	LUT3 #(
		.INIT('h82)
	) name13326 (
		_w6657_,
		_w11286_,
		_w11335_,
		_w13360_
	);
	LUT2 #(
		.INIT('h8)
	) name13327 (
		_w6334_,
		_w11382_,
		_w13361_
	);
	LUT4 #(
		.INIT('h2228)
	) name13328 (
		_w6650_,
		_w7695_,
		_w7750_,
		_w11285_,
		_w13362_
	);
	LUT2 #(
		.INIT('h1)
	) name13329 (
		_w13361_,
		_w13362_,
		_w13363_
	);
	LUT2 #(
		.INIT('h4)
	) name13330 (
		_w13360_,
		_w13363_,
		_w13364_
	);
	LUT3 #(
		.INIT('h1e)
	) name13331 (
		_w12841_,
		_w13048_,
		_w13049_,
		_w13365_
	);
	LUT4 #(
		.INIT('h009a)
	) name13332 (
		\a[2] ,
		_w13359_,
		_w13364_,
		_w13365_,
		_w13366_
	);
	LUT4 #(
		.INIT('h6500)
	) name13333 (
		\a[2] ,
		_w13359_,
		_w13364_,
		_w13365_,
		_w13367_
	);
	LUT4 #(
		.INIT('h54ab)
	) name13334 (
		_w12847_,
		_w13044_,
		_w13045_,
		_w13047_,
		_w13368_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13335 (
		_w6335_,
		_w11384_,
		_w11488_,
		_w11489_,
		_w13369_
	);
	LUT4 #(
		.INIT('h2228)
	) name13336 (
		_w6657_,
		_w7695_,
		_w7750_,
		_w11285_,
		_w13370_
	);
	LUT3 #(
		.INIT('h82)
	) name13337 (
		_w6334_,
		_w11280_,
		_w11282_,
		_w13371_
	);
	LUT3 #(
		.INIT('h07)
	) name13338 (
		_w6650_,
		_w11382_,
		_w13371_,
		_w13372_
	);
	LUT2 #(
		.INIT('h4)
	) name13339 (
		_w13370_,
		_w13372_,
		_w13373_
	);
	LUT4 #(
		.INIT('h2122)
	) name13340 (
		\a[2] ,
		_w13368_,
		_w13369_,
		_w13373_,
		_w13374_
	);
	LUT4 #(
		.INIT('h4844)
	) name13341 (
		\a[2] ,
		_w13368_,
		_w13369_,
		_w13373_,
		_w13375_
	);
	LUT4 #(
		.INIT('h2228)
	) name13342 (
		_w6334_,
		_w7935_,
		_w8077_,
		_w11279_,
		_w13376_
	);
	LUT4 #(
		.INIT('h007d)
	) name13343 (
		_w6650_,
		_w11280_,
		_w11282_,
		_w13376_,
		_w13377_
	);
	LUT3 #(
		.INIT('h70)
	) name13344 (
		_w6657_,
		_w11382_,
		_w13377_,
		_w13378_
	);
	LUT4 #(
		.INIT('h95aa)
	) name13345 (
		\a[2] ,
		_w6335_,
		_w12476_,
		_w13378_,
		_w13379_
	);
	LUT2 #(
		.INIT('h9)
	) name13346 (
		_w13044_,
		_w13046_,
		_w13380_
	);
	LUT3 #(
		.INIT('h1e)
	) name13347 (
		_w12862_,
		_w13042_,
		_w13043_,
		_w13381_
	);
	LUT3 #(
		.INIT('h82)
	) name13348 (
		_w6335_,
		_w11484_,
		_w11486_,
		_w13382_
	);
	LUT3 #(
		.INIT('h82)
	) name13349 (
		_w6657_,
		_w11280_,
		_w11282_,
		_w13383_
	);
	LUT2 #(
		.INIT('h8)
	) name13350 (
		_w6334_,
		_w11388_,
		_w13384_
	);
	LUT4 #(
		.INIT('h2228)
	) name13351 (
		_w6650_,
		_w7935_,
		_w8077_,
		_w11279_,
		_w13385_
	);
	LUT2 #(
		.INIT('h1)
	) name13352 (
		_w13384_,
		_w13385_,
		_w13386_
	);
	LUT2 #(
		.INIT('h4)
	) name13353 (
		_w13383_,
		_w13386_,
		_w13387_
	);
	LUT4 #(
		.INIT('h2122)
	) name13354 (
		\a[2] ,
		_w13381_,
		_w13382_,
		_w13387_,
		_w13388_
	);
	LUT4 #(
		.INIT('h4844)
	) name13355 (
		\a[2] ,
		_w13381_,
		_w13382_,
		_w13387_,
		_w13389_
	);
	LUT4 #(
		.INIT('h54ab)
	) name13356 (
		_w12868_,
		_w13038_,
		_w13039_,
		_w13041_,
		_w13390_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13357 (
		_w6335_,
		_w11390_,
		_w11482_,
		_w11483_,
		_w13391_
	);
	LUT4 #(
		.INIT('h2228)
	) name13358 (
		_w6657_,
		_w7935_,
		_w8077_,
		_w11279_,
		_w13392_
	);
	LUT3 #(
		.INIT('h82)
	) name13359 (
		_w6334_,
		_w11274_,
		_w11276_,
		_w13393_
	);
	LUT3 #(
		.INIT('h07)
	) name13360 (
		_w6650_,
		_w11388_,
		_w13393_,
		_w13394_
	);
	LUT2 #(
		.INIT('h4)
	) name13361 (
		_w13392_,
		_w13394_,
		_w13395_
	);
	LUT4 #(
		.INIT('h2122)
	) name13362 (
		\a[2] ,
		_w13390_,
		_w13391_,
		_w13395_,
		_w13396_
	);
	LUT4 #(
		.INIT('h4844)
	) name13363 (
		\a[2] ,
		_w13390_,
		_w13391_,
		_w13395_,
		_w13397_
	);
	LUT2 #(
		.INIT('h9)
	) name13364 (
		_w13038_,
		_w13040_,
		_w13398_
	);
	LUT4 #(
		.INIT('h2228)
	) name13365 (
		_w6334_,
		_w8466_,
		_w8541_,
		_w11273_,
		_w13399_
	);
	LUT4 #(
		.INIT('h007d)
	) name13366 (
		_w6650_,
		_w11274_,
		_w11276_,
		_w13399_,
		_w13400_
	);
	LUT3 #(
		.INIT('h70)
	) name13367 (
		_w6657_,
		_w11388_,
		_w13400_,
		_w13401_
	);
	LUT4 #(
		.INIT('h95aa)
	) name13368 (
		\a[2] ,
		_w6335_,
		_w12391_,
		_w13401_,
		_w13402_
	);
	LUT3 #(
		.INIT('h82)
	) name13369 (
		_w6335_,
		_w11478_,
		_w11480_,
		_w13403_
	);
	LUT3 #(
		.INIT('h82)
	) name13370 (
		_w6657_,
		_w11274_,
		_w11276_,
		_w13404_
	);
	LUT2 #(
		.INIT('h8)
	) name13371 (
		_w6334_,
		_w11394_,
		_w13405_
	);
	LUT4 #(
		.INIT('h2228)
	) name13372 (
		_w6650_,
		_w8466_,
		_w8541_,
		_w11273_,
		_w13406_
	);
	LUT2 #(
		.INIT('h1)
	) name13373 (
		_w13405_,
		_w13406_,
		_w13407_
	);
	LUT2 #(
		.INIT('h4)
	) name13374 (
		_w13404_,
		_w13407_,
		_w13408_
	);
	LUT3 #(
		.INIT('h1e)
	) name13375 (
		_w12883_,
		_w13036_,
		_w13037_,
		_w13409_
	);
	LUT4 #(
		.INIT('h009a)
	) name13376 (
		\a[2] ,
		_w13403_,
		_w13408_,
		_w13409_,
		_w13410_
	);
	LUT4 #(
		.INIT('h6500)
	) name13377 (
		\a[2] ,
		_w13403_,
		_w13408_,
		_w13409_,
		_w13411_
	);
	LUT4 #(
		.INIT('h54ab)
	) name13378 (
		_w12889_,
		_w13032_,
		_w13033_,
		_w13035_,
		_w13412_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13379 (
		_w6335_,
		_w11396_,
		_w11476_,
		_w11477_,
		_w13413_
	);
	LUT4 #(
		.INIT('h2228)
	) name13380 (
		_w6657_,
		_w8466_,
		_w8541_,
		_w11273_,
		_w13414_
	);
	LUT3 #(
		.INIT('h82)
	) name13381 (
		_w6334_,
		_w11268_,
		_w11270_,
		_w13415_
	);
	LUT3 #(
		.INIT('h07)
	) name13382 (
		_w6650_,
		_w11394_,
		_w13415_,
		_w13416_
	);
	LUT2 #(
		.INIT('h4)
	) name13383 (
		_w13414_,
		_w13416_,
		_w13417_
	);
	LUT4 #(
		.INIT('h2122)
	) name13384 (
		\a[2] ,
		_w13412_,
		_w13413_,
		_w13417_,
		_w13418_
	);
	LUT4 #(
		.INIT('h4844)
	) name13385 (
		\a[2] ,
		_w13412_,
		_w13413_,
		_w13417_,
		_w13419_
	);
	LUT4 #(
		.INIT('h2228)
	) name13386 (
		_w6334_,
		_w8794_,
		_w8994_,
		_w11267_,
		_w13420_
	);
	LUT4 #(
		.INIT('h007d)
	) name13387 (
		_w6650_,
		_w11268_,
		_w11270_,
		_w13420_,
		_w13421_
	);
	LUT3 #(
		.INIT('h70)
	) name13388 (
		_w6657_,
		_w11394_,
		_w13421_,
		_w13422_
	);
	LUT4 #(
		.INIT('h95aa)
	) name13389 (
		\a[2] ,
		_w6335_,
		_w12209_,
		_w13422_,
		_w13423_
	);
	LUT2 #(
		.INIT('h9)
	) name13390 (
		_w13032_,
		_w13034_,
		_w13424_
	);
	LUT3 #(
		.INIT('h1e)
	) name13391 (
		_w12904_,
		_w13030_,
		_w13031_,
		_w13425_
	);
	LUT3 #(
		.INIT('h82)
	) name13392 (
		_w6335_,
		_w11472_,
		_w11474_,
		_w13426_
	);
	LUT3 #(
		.INIT('h82)
	) name13393 (
		_w6657_,
		_w11268_,
		_w11270_,
		_w13427_
	);
	LUT2 #(
		.INIT('h8)
	) name13394 (
		_w6334_,
		_w11400_,
		_w13428_
	);
	LUT4 #(
		.INIT('h2228)
	) name13395 (
		_w6650_,
		_w8794_,
		_w8994_,
		_w11267_,
		_w13429_
	);
	LUT2 #(
		.INIT('h1)
	) name13396 (
		_w13428_,
		_w13429_,
		_w13430_
	);
	LUT2 #(
		.INIT('h4)
	) name13397 (
		_w13427_,
		_w13430_,
		_w13431_
	);
	LUT4 #(
		.INIT('h2122)
	) name13398 (
		\a[2] ,
		_w13425_,
		_w13426_,
		_w13431_,
		_w13432_
	);
	LUT4 #(
		.INIT('h4844)
	) name13399 (
		\a[2] ,
		_w13425_,
		_w13426_,
		_w13431_,
		_w13433_
	);
	LUT4 #(
		.INIT('h54ab)
	) name13400 (
		_w12910_,
		_w13026_,
		_w13027_,
		_w13029_,
		_w13434_
	);
	LUT3 #(
		.INIT('h82)
	) name13401 (
		_w6335_,
		_w11469_,
		_w11471_,
		_w13435_
	);
	LUT4 #(
		.INIT('h2228)
	) name13402 (
		_w6657_,
		_w8794_,
		_w8994_,
		_w11267_,
		_w13436_
	);
	LUT3 #(
		.INIT('h82)
	) name13403 (
		_w6334_,
		_w11262_,
		_w11264_,
		_w13437_
	);
	LUT3 #(
		.INIT('h07)
	) name13404 (
		_w6650_,
		_w11400_,
		_w13437_,
		_w13438_
	);
	LUT2 #(
		.INIT('h4)
	) name13405 (
		_w13436_,
		_w13438_,
		_w13439_
	);
	LUT4 #(
		.INIT('h2122)
	) name13406 (
		\a[2] ,
		_w13434_,
		_w13435_,
		_w13439_,
		_w13440_
	);
	LUT4 #(
		.INIT('h4844)
	) name13407 (
		\a[2] ,
		_w13434_,
		_w13435_,
		_w13439_,
		_w13441_
	);
	LUT2 #(
		.INIT('h9)
	) name13408 (
		_w13026_,
		_w13028_,
		_w13442_
	);
	LUT4 #(
		.INIT('h2228)
	) name13409 (
		_w6334_,
		_w9446_,
		_w9702_,
		_w11261_,
		_w13443_
	);
	LUT4 #(
		.INIT('h007d)
	) name13410 (
		_w6650_,
		_w11262_,
		_w11264_,
		_w13443_,
		_w13444_
	);
	LUT3 #(
		.INIT('h70)
	) name13411 (
		_w6657_,
		_w11400_,
		_w13444_,
		_w13445_
	);
	LUT4 #(
		.INIT('h6a55)
	) name13412 (
		\a[2] ,
		_w6335_,
		_w11967_,
		_w13445_,
		_w13446_
	);
	LUT3 #(
		.INIT('h82)
	) name13413 (
		_w6335_,
		_w11465_,
		_w11467_,
		_w13447_
	);
	LUT3 #(
		.INIT('h82)
	) name13414 (
		_w6657_,
		_w11262_,
		_w11264_,
		_w13448_
	);
	LUT2 #(
		.INIT('h8)
	) name13415 (
		_w6334_,
		_w11406_,
		_w13449_
	);
	LUT4 #(
		.INIT('h2228)
	) name13416 (
		_w6650_,
		_w9446_,
		_w9702_,
		_w11261_,
		_w13450_
	);
	LUT2 #(
		.INIT('h1)
	) name13417 (
		_w13449_,
		_w13450_,
		_w13451_
	);
	LUT2 #(
		.INIT('h4)
	) name13418 (
		_w13448_,
		_w13451_,
		_w13452_
	);
	LUT2 #(
		.INIT('h9)
	) name13419 (
		_w13023_,
		_w13025_,
		_w13453_
	);
	LUT4 #(
		.INIT('h009a)
	) name13420 (
		\a[2] ,
		_w13447_,
		_w13452_,
		_w13453_,
		_w13454_
	);
	LUT4 #(
		.INIT('h6500)
	) name13421 (
		\a[2] ,
		_w13447_,
		_w13452_,
		_w13453_,
		_w13455_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13422 (
		_w6335_,
		_w11408_,
		_w11463_,
		_w11464_,
		_w13456_
	);
	LUT4 #(
		.INIT('h2228)
	) name13423 (
		_w6657_,
		_w9446_,
		_w9702_,
		_w11261_,
		_w13457_
	);
	LUT3 #(
		.INIT('h82)
	) name13424 (
		_w6334_,
		_w11256_,
		_w11258_,
		_w13458_
	);
	LUT3 #(
		.INIT('h07)
	) name13425 (
		_w6650_,
		_w11406_,
		_w13458_,
		_w13459_
	);
	LUT2 #(
		.INIT('h4)
	) name13426 (
		_w13457_,
		_w13459_,
		_w13460_
	);
	LUT2 #(
		.INIT('h9)
	) name13427 (
		_w13020_,
		_w13022_,
		_w13461_
	);
	LUT4 #(
		.INIT('h009a)
	) name13428 (
		\a[2] ,
		_w13456_,
		_w13460_,
		_w13461_,
		_w13462_
	);
	LUT4 #(
		.INIT('h6500)
	) name13429 (
		\a[2] ,
		_w13456_,
		_w13460_,
		_w13461_,
		_w13463_
	);
	LUT3 #(
		.INIT('h82)
	) name13430 (
		_w6334_,
		_w10268_,
		_w11255_,
		_w13464_
	);
	LUT4 #(
		.INIT('h007d)
	) name13431 (
		_w6650_,
		_w11256_,
		_w11258_,
		_w13464_,
		_w13465_
	);
	LUT3 #(
		.INIT('h70)
	) name13432 (
		_w6657_,
		_w11406_,
		_w13465_,
		_w13466_
	);
	LUT4 #(
		.INIT('h95aa)
	) name13433 (
		\a[2] ,
		_w6335_,
		_w11796_,
		_w13466_,
		_w13467_
	);
	LUT2 #(
		.INIT('h9)
	) name13434 (
		_w13017_,
		_w13019_,
		_w13468_
	);
	LUT2 #(
		.INIT('h9)
	) name13435 (
		_w13014_,
		_w13016_,
		_w13469_
	);
	LUT3 #(
		.INIT('h82)
	) name13436 (
		_w6334_,
		_w10580_,
		_w11254_,
		_w13470_
	);
	LUT4 #(
		.INIT('h007d)
	) name13437 (
		_w6650_,
		_w10268_,
		_w11255_,
		_w13470_,
		_w13471_
	);
	LUT4 #(
		.INIT('h7d00)
	) name13438 (
		_w6657_,
		_w11256_,
		_w11258_,
		_w13471_,
		_w13472_
	);
	LUT4 #(
		.INIT('h7d00)
	) name13439 (
		_w6335_,
		_w11459_,
		_w11461_,
		_w13472_,
		_w13473_
	);
	LUT2 #(
		.INIT('h9)
	) name13440 (
		\a[2] ,
		_w13473_,
		_w13474_
	);
	LUT2 #(
		.INIT('h9)
	) name13441 (
		_w13011_,
		_w13013_,
		_w13475_
	);
	LUT3 #(
		.INIT('h82)
	) name13442 (
		_w6334_,
		_w10599_,
		_w11253_,
		_w13476_
	);
	LUT4 #(
		.INIT('h007d)
	) name13443 (
		_w6650_,
		_w10580_,
		_w11254_,
		_w13476_,
		_w13477_
	);
	LUT4 #(
		.INIT('h7d00)
	) name13444 (
		_w6657_,
		_w10268_,
		_w11255_,
		_w13477_,
		_w13478_
	);
	LUT4 #(
		.INIT('h7d00)
	) name13445 (
		_w6335_,
		_w11456_,
		_w11458_,
		_w13478_,
		_w13479_
	);
	LUT3 #(
		.INIT('h84)
	) name13446 (
		\a[2] ,
		_w13475_,
		_w13479_,
		_w13480_
	);
	LUT3 #(
		.INIT('h12)
	) name13447 (
		\a[2] ,
		_w13475_,
		_w13479_,
		_w13481_
	);
	LUT3 #(
		.INIT('h1e)
	) name13448 (
		_w12955_,
		_w13009_,
		_w13010_,
		_w13482_
	);
	LUT2 #(
		.INIT('h8)
	) name13449 (
		_w6334_,
		_w11415_,
		_w13483_
	);
	LUT4 #(
		.INIT('h007d)
	) name13450 (
		_w6650_,
		_w10599_,
		_w11253_,
		_w13483_,
		_w13484_
	);
	LUT4 #(
		.INIT('h7d00)
	) name13451 (
		_w6657_,
		_w10580_,
		_w11254_,
		_w13484_,
		_w13485_
	);
	LUT4 #(
		.INIT('h7d00)
	) name13452 (
		_w6335_,
		_w11453_,
		_w11455_,
		_w13485_,
		_w13486_
	);
	LUT3 #(
		.INIT('h84)
	) name13453 (
		\a[2] ,
		_w13482_,
		_w13486_,
		_w13487_
	);
	LUT3 #(
		.INIT('h12)
	) name13454 (
		\a[2] ,
		_w13482_,
		_w13486_,
		_w13488_
	);
	LUT4 #(
		.INIT('h54ab)
	) name13455 (
		_w12961_,
		_w13005_,
		_w13006_,
		_w13008_,
		_w13489_
	);
	LUT3 #(
		.INIT('h82)
	) name13456 (
		_w6334_,
		_w11249_,
		_w11251_,
		_w13490_
	);
	LUT3 #(
		.INIT('h07)
	) name13457 (
		_w6650_,
		_w11415_,
		_w13490_,
		_w13491_
	);
	LUT4 #(
		.INIT('h7d00)
	) name13458 (
		_w6657_,
		_w10599_,
		_w11253_,
		_w13491_,
		_w13492_
	);
	LUT4 #(
		.INIT('h7d00)
	) name13459 (
		_w6335_,
		_w11450_,
		_w11452_,
		_w13492_,
		_w13493_
	);
	LUT3 #(
		.INIT('h84)
	) name13460 (
		\a[2] ,
		_w13489_,
		_w13493_,
		_w13494_
	);
	LUT3 #(
		.INIT('h12)
	) name13461 (
		\a[2] ,
		_w13489_,
		_w13493_,
		_w13495_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13462 (
		_w6334_,
		_w10945_,
		_w11246_,
		_w11248_,
		_w13496_
	);
	LUT4 #(
		.INIT('h007d)
	) name13463 (
		_w6650_,
		_w11249_,
		_w11251_,
		_w13496_,
		_w13497_
	);
	LUT3 #(
		.INIT('h70)
	) name13464 (
		_w6657_,
		_w11415_,
		_w13497_,
		_w13498_
	);
	LUT4 #(
		.INIT('h95aa)
	) name13465 (
		\a[2] ,
		_w6335_,
		_w11675_,
		_w13498_,
		_w13499_
	);
	LUT2 #(
		.INIT('h9)
	) name13466 (
		_w13005_,
		_w13007_,
		_w13500_
	);
	LUT2 #(
		.INIT('h4)
	) name13467 (
		_w13499_,
		_w13500_,
		_w13501_
	);
	LUT2 #(
		.INIT('h2)
	) name13468 (
		_w13499_,
		_w13500_,
		_w13502_
	);
	LUT3 #(
		.INIT('h82)
	) name13469 (
		_w6335_,
		_w11445_,
		_w11447_,
		_w13503_
	);
	LUT3 #(
		.INIT('h82)
	) name13470 (
		_w6657_,
		_w11249_,
		_w11251_,
		_w13504_
	);
	LUT2 #(
		.INIT('h8)
	) name13471 (
		_w6334_,
		_w11421_,
		_w13505_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13472 (
		_w6650_,
		_w10945_,
		_w11246_,
		_w11248_,
		_w13506_
	);
	LUT2 #(
		.INIT('h1)
	) name13473 (
		_w13505_,
		_w13506_,
		_w13507_
	);
	LUT2 #(
		.INIT('h4)
	) name13474 (
		_w13504_,
		_w13507_,
		_w13508_
	);
	LUT2 #(
		.INIT('h9)
	) name13475 (
		_w13002_,
		_w13004_,
		_w13509_
	);
	LUT4 #(
		.INIT('h6500)
	) name13476 (
		\a[2] ,
		_w13503_,
		_w13508_,
		_w13509_,
		_w13510_
	);
	LUT4 #(
		.INIT('h009a)
	) name13477 (
		\a[2] ,
		_w13503_,
		_w13508_,
		_w13509_,
		_w13511_
	);
	LUT2 #(
		.INIT('h9)
	) name13478 (
		_w12999_,
		_w13001_,
		_w13512_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13479 (
		_w6335_,
		_w11423_,
		_w11443_,
		_w11444_,
		_w13513_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13480 (
		_w6657_,
		_w10945_,
		_w11246_,
		_w11248_,
		_w13514_
	);
	LUT3 #(
		.INIT('h82)
	) name13481 (
		_w6334_,
		_w11241_,
		_w11243_,
		_w13515_
	);
	LUT3 #(
		.INIT('h07)
	) name13482 (
		_w6650_,
		_w11421_,
		_w13515_,
		_w13516_
	);
	LUT2 #(
		.INIT('h4)
	) name13483 (
		_w13514_,
		_w13516_,
		_w13517_
	);
	LUT4 #(
		.INIT('h4844)
	) name13484 (
		\a[2] ,
		_w13512_,
		_w13513_,
		_w13517_,
		_w13518_
	);
	LUT4 #(
		.INIT('h2122)
	) name13485 (
		\a[2] ,
		_w13512_,
		_w13513_,
		_w13517_,
		_w13519_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13486 (
		_w6334_,
		_w10968_,
		_w11238_,
		_w11240_,
		_w13520_
	);
	LUT4 #(
		.INIT('h007d)
	) name13487 (
		_w6650_,
		_w11241_,
		_w11243_,
		_w13520_,
		_w13521_
	);
	LUT3 #(
		.INIT('h70)
	) name13488 (
		_w6657_,
		_w11421_,
		_w13521_,
		_w13522_
	);
	LUT4 #(
		.INIT('h95aa)
	) name13489 (
		\a[2] ,
		_w6335_,
		_w11569_,
		_w13522_,
		_w13523_
	);
	LUT3 #(
		.INIT('h8a)
	) name13490 (
		\a[5] ,
		_w12982_,
		_w12981_,
		_w13524_
	);
	LUT2 #(
		.INIT('h9)
	) name13491 (
		_w12990_,
		_w13524_,
		_w13525_
	);
	LUT3 #(
		.INIT('h82)
	) name13492 (
		_w6335_,
		_w11439_,
		_w11441_,
		_w13526_
	);
	LUT3 #(
		.INIT('h82)
	) name13493 (
		_w6657_,
		_w11241_,
		_w11243_,
		_w13527_
	);
	LUT2 #(
		.INIT('h8)
	) name13494 (
		_w6334_,
		_w11427_,
		_w13528_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13495 (
		_w6650_,
		_w10968_,
		_w11238_,
		_w11240_,
		_w13529_
	);
	LUT2 #(
		.INIT('h1)
	) name13496 (
		_w13528_,
		_w13529_,
		_w13530_
	);
	LUT2 #(
		.INIT('h4)
	) name13497 (
		_w13527_,
		_w13530_,
		_w13531_
	);
	LUT3 #(
		.INIT('h65)
	) name13498 (
		\a[2] ,
		_w13526_,
		_w13531_,
		_w13532_
	);
	LUT3 #(
		.INIT('h28)
	) name13499 (
		_w6335_,
		_w11431_,
		_w11435_,
		_w13533_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13500 (
		_w6334_,
		_w10991_,
		_w11230_,
		_w11232_,
		_w13534_
	);
	LUT4 #(
		.INIT('h007d)
	) name13501 (
		_w6650_,
		_w11233_,
		_w11235_,
		_w13534_,
		_w13535_
	);
	LUT3 #(
		.INIT('h70)
	) name13502 (
		_w6657_,
		_w11427_,
		_w13535_,
		_w13536_
	);
	LUT2 #(
		.INIT('h4)
	) name13503 (
		\a[2] ,
		_w11434_,
		_w13537_
	);
	LUT3 #(
		.INIT('h0b)
	) name13504 (
		_w13533_,
		_w13536_,
		_w13537_,
		_w13538_
	);
	LUT4 #(
		.INIT('h3c28)
	) name13505 (
		_w6333_,
		_w11233_,
		_w11235_,
		_w11581_,
		_w13539_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13506 (
		_w10590_,
		_w10991_,
		_w11230_,
		_w11232_,
		_w13540_
	);
	LUT2 #(
		.INIT('h1)
	) name13507 (
		_w11434_,
		_w13540_,
		_w13541_
	);
	LUT4 #(
		.INIT('h0233)
	) name13508 (
		\a[0] ,
		_w12982_,
		_w13539_,
		_w13541_,
		_w13542_
	);
	LUT4 #(
		.INIT('h00ef)
	) name13509 (
		\a[2] ,
		_w13533_,
		_w13536_,
		_w13542_,
		_w13543_
	);
	LUT2 #(
		.INIT('h4)
	) name13510 (
		_w13538_,
		_w13543_,
		_w13544_
	);
	LUT3 #(
		.INIT('h20)
	) name13511 (
		\a[5] ,
		_w34_,
		_w11434_,
		_w13545_
	);
	LUT2 #(
		.INIT('h9)
	) name13512 (
		_w12981_,
		_w13545_,
		_w13546_
	);
	LUT3 #(
		.INIT('h82)
	) name13513 (
		_w6335_,
		_w11436_,
		_w11438_,
		_w13547_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13514 (
		_w6657_,
		_w10968_,
		_w11238_,
		_w11240_,
		_w13548_
	);
	LUT3 #(
		.INIT('h82)
	) name13515 (
		_w6334_,
		_w11233_,
		_w11235_,
		_w13549_
	);
	LUT3 #(
		.INIT('h07)
	) name13516 (
		_w6650_,
		_w11427_,
		_w13549_,
		_w13550_
	);
	LUT2 #(
		.INIT('h4)
	) name13517 (
		_w13548_,
		_w13550_,
		_w13551_
	);
	LUT3 #(
		.INIT('h9a)
	) name13518 (
		\a[2] ,
		_w13547_,
		_w13551_,
		_w13552_
	);
	LUT3 #(
		.INIT('h8e)
	) name13519 (
		_w13544_,
		_w13546_,
		_w13552_,
		_w13553_
	);
	LUT4 #(
		.INIT('h022a)
	) name13520 (
		_w13523_,
		_w13525_,
		_w13532_,
		_w13553_,
		_w13554_
	);
	LUT2 #(
		.INIT('h9)
	) name13521 (
		_w12996_,
		_w12998_,
		_w13555_
	);
	LUT4 #(
		.INIT('h5440)
	) name13522 (
		_w13523_,
		_w13525_,
		_w13532_,
		_w13553_,
		_w13556_
	);
	LUT4 #(
		.INIT('h5510)
	) name13523 (
		_w13519_,
		_w13554_,
		_w13555_,
		_w13556_,
		_w13557_
	);
	LUT4 #(
		.INIT('h4445)
	) name13524 (
		_w13510_,
		_w13511_,
		_w13518_,
		_w13557_,
		_w13558_
	);
	LUT3 #(
		.INIT('h54)
	) name13525 (
		_w13501_,
		_w13502_,
		_w13558_,
		_w13559_
	);
	LUT3 #(
		.INIT('h54)
	) name13526 (
		_w13494_,
		_w13495_,
		_w13559_,
		_w13560_
	);
	LUT3 #(
		.INIT('h54)
	) name13527 (
		_w13487_,
		_w13488_,
		_w13560_,
		_w13561_
	);
	LUT3 #(
		.INIT('h54)
	) name13528 (
		_w13480_,
		_w13481_,
		_w13561_,
		_w13562_
	);
	LUT3 #(
		.INIT('h8e)
	) name13529 (
		_w13469_,
		_w13474_,
		_w13562_,
		_w13563_
	);
	LUT4 #(
		.INIT('h0445)
	) name13530 (
		_w13463_,
		_w13467_,
		_w13468_,
		_w13563_,
		_w13564_
	);
	LUT4 #(
		.INIT('h4445)
	) name13531 (
		_w13454_,
		_w13455_,
		_w13462_,
		_w13564_,
		_w13565_
	);
	LUT4 #(
		.INIT('h0115)
	) name13532 (
		_w13441_,
		_w13442_,
		_w13446_,
		_w13565_,
		_w13566_
	);
	LUT4 #(
		.INIT('h4445)
	) name13533 (
		_w13432_,
		_w13433_,
		_w13440_,
		_w13566_,
		_w13567_
	);
	LUT4 #(
		.INIT('h0445)
	) name13534 (
		_w13419_,
		_w13423_,
		_w13424_,
		_w13567_,
		_w13568_
	);
	LUT4 #(
		.INIT('h4445)
	) name13535 (
		_w13410_,
		_w13411_,
		_w13418_,
		_w13568_,
		_w13569_
	);
	LUT4 #(
		.INIT('h1051)
	) name13536 (
		_w13397_,
		_w13398_,
		_w13402_,
		_w13569_,
		_w13570_
	);
	LUT4 #(
		.INIT('h4445)
	) name13537 (
		_w13388_,
		_w13389_,
		_w13396_,
		_w13570_,
		_w13571_
	);
	LUT4 #(
		.INIT('h0445)
	) name13538 (
		_w13375_,
		_w13379_,
		_w13380_,
		_w13571_,
		_w13572_
	);
	LUT4 #(
		.INIT('h4445)
	) name13539 (
		_w13366_,
		_w13367_,
		_w13374_,
		_w13572_,
		_w13573_
	);
	LUT4 #(
		.INIT('h0115)
	) name13540 (
		_w13353_,
		_w13354_,
		_w13358_,
		_w13573_,
		_w13574_
	);
	LUT4 #(
		.INIT('h4445)
	) name13541 (
		_w13344_,
		_w13345_,
		_w13352_,
		_w13574_,
		_w13575_
	);
	LUT4 #(
		.INIT('h32cd)
	) name13542 (
		_w13061_,
		_w13100_,
		_w13101_,
		_w13289_,
		_w13576_
	);
	LUT4 #(
		.INIT('h2228)
	) name13543 (
		_w6334_,
		_w11549_,
		_w11373_,
		_w11375_,
		_w13577_
	);
	LUT4 #(
		.INIT('h007d)
	) name13544 (
		_w6650_,
		_w13062_,
		_w13099_,
		_w13577_,
		_w13578_
	);
	LUT3 #(
		.INIT('h70)
	) name13545 (
		_w6657_,
		_w13247_,
		_w13578_,
		_w13579_
	);
	LUT4 #(
		.INIT('h95aa)
	) name13546 (
		\a[2] ,
		_w6335_,
		_w13576_,
		_w13579_,
		_w13580_
	);
	LUT3 #(
		.INIT('h8e)
	) name13547 (
		_w13336_,
		_w13575_,
		_w13580_,
		_w13581_
	);
	LUT4 #(
		.INIT('h1501)
	) name13548 (
		_w13335_,
		_w13336_,
		_w13575_,
		_w13580_,
		_w13582_
	);
	LUT4 #(
		.INIT('h80a8)
	) name13549 (
		_w13335_,
		_w13336_,
		_w13575_,
		_w13580_,
		_w13583_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13550 (
		_w6335_,
		_w13288_,
		_w13290_,
		_w13291_,
		_w13584_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13551 (
		_w6657_,
		_w13243_,
		_w13245_,
		_w13285_,
		_w13585_
	);
	LUT3 #(
		.INIT('h82)
	) name13552 (
		_w6334_,
		_w13062_,
		_w13099_,
		_w13586_
	);
	LUT3 #(
		.INIT('h07)
	) name13553 (
		_w6650_,
		_w13247_,
		_w13586_,
		_w13587_
	);
	LUT2 #(
		.INIT('h4)
	) name13554 (
		_w13585_,
		_w13587_,
		_w13588_
	);
	LUT3 #(
		.INIT('h9a)
	) name13555 (
		\a[2] ,
		_w13584_,
		_w13588_,
		_w13589_
	);
	LUT3 #(
		.INIT('h45)
	) name13556 (
		_w13582_,
		_w13583_,
		_w13589_,
		_w13590_
	);
	LUT4 #(
		.INIT('h80a8)
	) name13557 (
		_w13334_,
		_w13335_,
		_w13581_,
		_w13589_,
		_w13591_
	);
	LUT4 #(
		.INIT('h010f)
	) name13558 (
		_w12798_,
		_w13060_,
		_w13199_,
		_w13200_,
		_w13592_
	);
	LUT4 #(
		.INIT('h2228)
	) name13559 (
		_w5524_,
		_w11549_,
		_w11373_,
		_w11375_,
		_w13593_
	);
	LUT4 #(
		.INIT('h007d)
	) name13560 (
		_w6031_,
		_w13062_,
		_w13099_,
		_w13593_,
		_w13594_
	);
	LUT3 #(
		.INIT('h70)
	) name13561 (
		_w6324_,
		_w13247_,
		_w13594_,
		_w13595_
	);
	LUT4 #(
		.INIT('h95aa)
	) name13562 (
		\a[5] ,
		_w35_,
		_w13576_,
		_w13595_,
		_w13596_
	);
	LUT4 #(
		.INIT('h010f)
	) name13563 (
		_w12794_,
		_w12796_,
		_w13196_,
		_w13197_,
		_w13597_
	);
	LUT4 #(
		.INIT('h010f)
	) name13564 (
		_w12785_,
		_w12787_,
		_w13187_,
		_w13188_,
		_w13598_
	);
	LUT4 #(
		.INIT('h2228)
	) name13565 (
		_w4458_,
		_w7935_,
		_w8077_,
		_w11279_,
		_w13599_
	);
	LUT4 #(
		.INIT('h007d)
	) name13566 (
		_w4684_,
		_w11280_,
		_w11282_,
		_w13599_,
		_w13600_
	);
	LUT3 #(
		.INIT('h70)
	) name13567 (
		_w4700_,
		_w11382_,
		_w13600_,
		_w13601_
	);
	LUT4 #(
		.INIT('h95aa)
	) name13568 (
		\a[11] ,
		_w4459_,
		_w12476_,
		_w13601_,
		_w13602_
	);
	LUT4 #(
		.INIT('h010f)
	) name13569 (
		_w12781_,
		_w12783_,
		_w13184_,
		_w13185_,
		_w13603_
	);
	LUT4 #(
		.INIT('h010f)
	) name13570 (
		_w12772_,
		_w12774_,
		_w13175_,
		_w13176_,
		_w13604_
	);
	LUT4 #(
		.INIT('h2228)
	) name13571 (
		_w3709_,
		_w8794_,
		_w8994_,
		_w11267_,
		_w13605_
	);
	LUT4 #(
		.INIT('h007d)
	) name13572 (
		_w3877_,
		_w11268_,
		_w11270_,
		_w13605_,
		_w13606_
	);
	LUT3 #(
		.INIT('h70)
	) name13573 (
		_w3886_,
		_w11394_,
		_w13606_,
		_w13607_
	);
	LUT4 #(
		.INIT('h95aa)
	) name13574 (
		\a[17] ,
		_w3710_,
		_w12209_,
		_w13607_,
		_w13608_
	);
	LUT4 #(
		.INIT('h010f)
	) name13575 (
		_w12768_,
		_w12770_,
		_w13172_,
		_w13173_,
		_w13609_
	);
	LUT3 #(
		.INIT('h32)
	) name13576 (
		_w13121_,
		_w13162_,
		_w13163_,
		_w13610_
	);
	LUT3 #(
		.INIT('h82)
	) name13577 (
		_w3214_,
		_w10268_,
		_w11255_,
		_w13611_
	);
	LUT4 #(
		.INIT('h007d)
	) name13578 (
		_w3249_,
		_w11256_,
		_w11258_,
		_w13611_,
		_w13612_
	);
	LUT3 #(
		.INIT('h70)
	) name13579 (
		_w3262_,
		_w11406_,
		_w13612_,
		_w13613_
	);
	LUT4 #(
		.INIT('h95aa)
	) name13580 (
		\a[23] ,
		_w37_,
		_w11796_,
		_w13613_,
		_w13614_
	);
	LUT3 #(
		.INIT('h32)
	) name13581 (
		_w13126_,
		_w13158_,
		_w13159_,
		_w13615_
	);
	LUT3 #(
		.INIT('h82)
	) name13582 (
		_w2550_,
		_w11445_,
		_w11447_,
		_w13616_
	);
	LUT3 #(
		.INIT('h82)
	) name13583 (
		_w2854_,
		_w11249_,
		_w11251_,
		_w13617_
	);
	LUT2 #(
		.INIT('h8)
	) name13584 (
		_w2549_,
		_w11421_,
		_w13618_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13585 (
		_w2617_,
		_w10945_,
		_w11246_,
		_w11248_,
		_w13619_
	);
	LUT2 #(
		.INIT('h1)
	) name13586 (
		_w13618_,
		_w13619_,
		_w13620_
	);
	LUT2 #(
		.INIT('h4)
	) name13587 (
		_w13617_,
		_w13620_,
		_w13621_
	);
	LUT3 #(
		.INIT('h32)
	) name13588 (
		_w13132_,
		_w13146_,
		_w13147_,
		_w13622_
	);
	LUT3 #(
		.INIT('h80)
	) name13589 (
		_w1669_,
		_w2370_,
		_w7212_,
		_w13623_
	);
	LUT3 #(
		.INIT('h80)
	) name13590 (
		_w3345_,
		_w7219_,
		_w13623_,
		_w13624_
	);
	LUT4 #(
		.INIT('h4000)
	) name13591 (
		_w437_,
		_w713_,
		_w924_,
		_w1472_,
		_w13625_
	);
	LUT4 #(
		.INIT('h4000)
	) name13592 (
		_w482_,
		_w1668_,
		_w1776_,
		_w1777_,
		_w13626_
	);
	LUT4 #(
		.INIT('h8000)
	) name13593 (
		_w2821_,
		_w2824_,
		_w13625_,
		_w13626_,
		_w13627_
	);
	LUT4 #(
		.INIT('h8000)
	) name13594 (
		_w3112_,
		_w3117_,
		_w13624_,
		_w13627_,
		_w13628_
	);
	LUT2 #(
		.INIT('h8)
	) name13595 (
		_w7308_,
		_w13628_,
		_w13629_
	);
	LUT3 #(
		.INIT('h82)
	) name13596 (
		_w377_,
		_w11439_,
		_w11441_,
		_w13630_
	);
	LUT3 #(
		.INIT('h82)
	) name13597 (
		_w2527_,
		_w11241_,
		_w11243_,
		_w13631_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13598 (
		_w2407_,
		_w10968_,
		_w11238_,
		_w11240_,
		_w13632_
	);
	LUT2 #(
		.INIT('h8)
	) name13599 (
		_w376_,
		_w11427_,
		_w13633_
	);
	LUT2 #(
		.INIT('h1)
	) name13600 (
		_w13632_,
		_w13633_,
		_w13634_
	);
	LUT2 #(
		.INIT('h4)
	) name13601 (
		_w13631_,
		_w13634_,
		_w13635_
	);
	LUT2 #(
		.INIT('h4)
	) name13602 (
		_w13630_,
		_w13635_,
		_w13636_
	);
	LUT3 #(
		.INIT('h45)
	) name13603 (
		_w13629_,
		_w13630_,
		_w13635_,
		_w13637_
	);
	LUT3 #(
		.INIT('h20)
	) name13604 (
		_w13629_,
		_w13630_,
		_w13635_,
		_w13638_
	);
	LUT3 #(
		.INIT('h9a)
	) name13605 (
		_w13629_,
		_w13630_,
		_w13635_,
		_w13639_
	);
	LUT2 #(
		.INIT('h9)
	) name13606 (
		_w13622_,
		_w13639_,
		_w13640_
	);
	LUT4 #(
		.INIT('h6500)
	) name13607 (
		\a[29] ,
		_w13616_,
		_w13621_,
		_w13640_,
		_w13641_
	);
	LUT4 #(
		.INIT('h9a65)
	) name13608 (
		\a[29] ,
		_w13616_,
		_w13621_,
		_w13640_,
		_w13642_
	);
	LUT3 #(
		.INIT('h1e)
	) name13609 (
		_w13150_,
		_w13152_,
		_w13642_,
		_w13643_
	);
	LUT2 #(
		.INIT('h8)
	) name13610 (
		_w2874_,
		_w11415_,
		_w13644_
	);
	LUT4 #(
		.INIT('h007d)
	) name13611 (
		_w2975_,
		_w10599_,
		_w11253_,
		_w13644_,
		_w13645_
	);
	LUT4 #(
		.INIT('h7d00)
	) name13612 (
		_w2986_,
		_w10580_,
		_w11254_,
		_w13645_,
		_w13646_
	);
	LUT4 #(
		.INIT('h7d00)
	) name13613 (
		_w2875_,
		_w11453_,
		_w11455_,
		_w13646_,
		_w13647_
	);
	LUT3 #(
		.INIT('h84)
	) name13614 (
		\a[26] ,
		_w13643_,
		_w13647_,
		_w13648_
	);
	LUT3 #(
		.INIT('h12)
	) name13615 (
		\a[26] ,
		_w13643_,
		_w13647_,
		_w13649_
	);
	LUT3 #(
		.INIT('h69)
	) name13616 (
		\a[26] ,
		_w13643_,
		_w13647_,
		_w13650_
	);
	LUT2 #(
		.INIT('h9)
	) name13617 (
		_w13615_,
		_w13650_,
		_w13651_
	);
	LUT2 #(
		.INIT('h4)
	) name13618 (
		_w13614_,
		_w13651_,
		_w13652_
	);
	LUT2 #(
		.INIT('h2)
	) name13619 (
		_w13614_,
		_w13651_,
		_w13653_
	);
	LUT2 #(
		.INIT('h9)
	) name13620 (
		_w13614_,
		_w13651_,
		_w13654_
	);
	LUT2 #(
		.INIT('h9)
	) name13621 (
		_w13610_,
		_w13654_,
		_w13655_
	);
	LUT4 #(
		.INIT('h2228)
	) name13622 (
		_w3311_,
		_w9446_,
		_w9702_,
		_w11261_,
		_w13656_
	);
	LUT4 #(
		.INIT('h007d)
	) name13623 (
		_w3645_,
		_w11262_,
		_w11264_,
		_w13656_,
		_w13657_
	);
	LUT3 #(
		.INIT('h70)
	) name13624 (
		_w3654_,
		_w11400_,
		_w13657_,
		_w13658_
	);
	LUT4 #(
		.INIT('h95aa)
	) name13625 (
		\a[20] ,
		_w3312_,
		_w11967_,
		_w13658_,
		_w13659_
	);
	LUT2 #(
		.INIT('h2)
	) name13626 (
		_w13655_,
		_w13659_,
		_w13660_
	);
	LUT2 #(
		.INIT('h4)
	) name13627 (
		_w13655_,
		_w13659_,
		_w13661_
	);
	LUT2 #(
		.INIT('h9)
	) name13628 (
		_w13655_,
		_w13659_,
		_w13662_
	);
	LUT2 #(
		.INIT('h9)
	) name13629 (
		_w13609_,
		_w13662_,
		_w13663_
	);
	LUT2 #(
		.INIT('h4)
	) name13630 (
		_w13608_,
		_w13663_,
		_w13664_
	);
	LUT2 #(
		.INIT('h2)
	) name13631 (
		_w13608_,
		_w13663_,
		_w13665_
	);
	LUT2 #(
		.INIT('h9)
	) name13632 (
		_w13608_,
		_w13663_,
		_w13666_
	);
	LUT2 #(
		.INIT('h9)
	) name13633 (
		_w13604_,
		_w13666_,
		_w13667_
	);
	LUT4 #(
		.INIT('h2228)
	) name13634 (
		_w4033_,
		_w8466_,
		_w8541_,
		_w11273_,
		_w13668_
	);
	LUT4 #(
		.INIT('h007d)
	) name13635 (
		_w4367_,
		_w11274_,
		_w11276_,
		_w13668_,
		_w13669_
	);
	LUT3 #(
		.INIT('h70)
	) name13636 (
		_w4382_,
		_w11388_,
		_w13669_,
		_w13670_
	);
	LUT4 #(
		.INIT('h95aa)
	) name13637 (
		\a[14] ,
		_w4034_,
		_w12391_,
		_w13670_,
		_w13671_
	);
	LUT2 #(
		.INIT('h2)
	) name13638 (
		_w13667_,
		_w13671_,
		_w13672_
	);
	LUT2 #(
		.INIT('h4)
	) name13639 (
		_w13667_,
		_w13671_,
		_w13673_
	);
	LUT2 #(
		.INIT('h9)
	) name13640 (
		_w13667_,
		_w13671_,
		_w13674_
	);
	LUT2 #(
		.INIT('h9)
	) name13641 (
		_w13603_,
		_w13674_,
		_w13675_
	);
	LUT2 #(
		.INIT('h4)
	) name13642 (
		_w13602_,
		_w13675_,
		_w13676_
	);
	LUT2 #(
		.INIT('h2)
	) name13643 (
		_w13602_,
		_w13675_,
		_w13677_
	);
	LUT2 #(
		.INIT('h9)
	) name13644 (
		_w13602_,
		_w13675_,
		_w13678_
	);
	LUT2 #(
		.INIT('h9)
	) name13645 (
		_w13598_,
		_w13678_,
		_w13679_
	);
	LUT4 #(
		.INIT('h2228)
	) name13646 (
		_w4875_,
		_w7695_,
		_w7750_,
		_w11285_,
		_w13680_
	);
	LUT4 #(
		.INIT('h007d)
	) name13647 (
		_w5271_,
		_w11286_,
		_w11335_,
		_w13680_,
		_w13681_
	);
	LUT3 #(
		.INIT('h70)
	) name13648 (
		_w5286_,
		_w11377_,
		_w13681_,
		_w13682_
	);
	LUT4 #(
		.INIT('h95aa)
	) name13649 (
		\a[8] ,
		_w4876_,
		_w12799_,
		_w13682_,
		_w13683_
	);
	LUT2 #(
		.INIT('h2)
	) name13650 (
		_w13679_,
		_w13683_,
		_w13684_
	);
	LUT2 #(
		.INIT('h4)
	) name13651 (
		_w13679_,
		_w13683_,
		_w13685_
	);
	LUT2 #(
		.INIT('h9)
	) name13652 (
		_w13679_,
		_w13683_,
		_w13686_
	);
	LUT2 #(
		.INIT('h9)
	) name13653 (
		_w13597_,
		_w13686_,
		_w13687_
	);
	LUT2 #(
		.INIT('h4)
	) name13654 (
		_w13596_,
		_w13687_,
		_w13688_
	);
	LUT2 #(
		.INIT('h2)
	) name13655 (
		_w13596_,
		_w13687_,
		_w13689_
	);
	LUT2 #(
		.INIT('h9)
	) name13656 (
		_w13596_,
		_w13687_,
		_w13690_
	);
	LUT2 #(
		.INIT('h9)
	) name13657 (
		_w13592_,
		_w13690_,
		_w13691_
	);
	LUT4 #(
		.INIT('h0f01)
	) name13658 (
		_w13264_,
		_w13266_,
		_w13315_,
		_w13316_,
		_w13692_
	);
	LUT3 #(
		.INIT('h0d)
	) name13659 (
		_w13301_,
		_w13307_,
		_w13308_,
		_w13693_
	);
	LUT3 #(
		.INIT('h08)
	) name13660 (
		_w279_,
		_w350_,
		_w420_,
		_w13694_
	);
	LUT3 #(
		.INIT('h80)
	) name13661 (
		_w486_,
		_w13302_,
		_w13694_,
		_w13695_
	);
	LUT4 #(
		.INIT('h0df2)
	) name13662 (
		_w13301_,
		_w13307_,
		_w13308_,
		_w13695_,
		_w13696_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13663 (
		_w377_,
		_w6998_,
		_w7133_,
		_w7134_,
		_w13697_
	);
	LUT4 #(
		.INIT('h04c8)
	) name13664 (
		_w2411_,
		_w2527_,
		_w6983_,
		_w6993_,
		_w13698_
	);
	LUT3 #(
		.INIT('h82)
	) name13665 (
		_w376_,
		_w2546_,
		_w6981_,
		_w13699_
	);
	LUT3 #(
		.INIT('h07)
	) name13666 (
		_w2407_,
		_w6996_,
		_w13699_,
		_w13700_
	);
	LUT2 #(
		.INIT('h4)
	) name13667 (
		_w13698_,
		_w13700_,
		_w13701_
	);
	LUT2 #(
		.INIT('h4)
	) name13668 (
		_w13697_,
		_w13701_,
		_w13702_
	);
	LUT4 #(
		.INIT('h147d)
	) name13669 (
		_w13299_,
		_w13301_,
		_w13309_,
		_w13313_,
		_w13703_
	);
	LUT3 #(
		.INIT('h90)
	) name13670 (
		_w13696_,
		_w13702_,
		_w13703_,
		_w13704_
	);
	LUT3 #(
		.INIT('h69)
	) name13671 (
		_w13696_,
		_w13702_,
		_w13703_,
		_w13705_
	);
	LUT4 #(
		.INIT('h0a02)
	) name13672 (
		_w2550_,
		_w7169_,
		_w7419_,
		_w7686_,
		_w13706_
	);
	LUT4 #(
		.INIT('h3111)
	) name13673 (
		_w2617_,
		_w2854_,
		_w7136_,
		_w7167_,
		_w13707_
	);
	LUT3 #(
		.INIT('h28)
	) name13674 (
		_w2549_,
		_w7136_,
		_w7168_,
		_w13708_
	);
	LUT3 #(
		.INIT('h0e)
	) name13675 (
		_w7244_,
		_w13707_,
		_w13708_,
		_w13709_
	);
	LUT4 #(
		.INIT('h4844)
	) name13676 (
		\a[29] ,
		_w13705_,
		_w13706_,
		_w13709_,
		_w13710_
	);
	LUT4 #(
		.INIT('h9699)
	) name13677 (
		\a[29] ,
		_w13705_,
		_w13706_,
		_w13709_,
		_w13711_
	);
	LUT2 #(
		.INIT('h4)
	) name13678 (
		_w13692_,
		_w13711_,
		_w13712_
	);
	LUT2 #(
		.INIT('h9)
	) name13679 (
		_w13692_,
		_w13711_,
		_w13713_
	);
	LUT4 #(
		.INIT('h4d00)
	) name13680 (
		_w13293_,
		_w13318_,
		_w13319_,
		_w13713_,
		_w13714_
	);
	LUT4 #(
		.INIT('h00b2)
	) name13681 (
		_w13293_,
		_w13318_,
		_w13319_,
		_w13713_,
		_w13715_
	);
	LUT4 #(
		.INIT('h32cd)
	) name13682 (
		_w13293_,
		_w13320_,
		_w13321_,
		_w13713_,
		_w13716_
	);
	LUT4 #(
		.INIT('h1244)
	) name13683 (
		_w13293_,
		_w13320_,
		_w13321_,
		_w13713_,
		_w13717_
	);
	LUT4 #(
		.INIT('h8679)
	) name13684 (
		_w13293_,
		_w13320_,
		_w13322_,
		_w13713_,
		_w13718_
	);
	LUT4 #(
		.INIT('hdc00)
	) name13685 (
		_w13292_,
		_w13323_,
		_w13325_,
		_w13718_,
		_w13719_
	);
	LUT4 #(
		.INIT('h32cd)
	) name13686 (
		_w13292_,
		_w13323_,
		_w13324_,
		_w13718_,
		_w13720_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13687 (
		_w6334_,
		_w13243_,
		_w13245_,
		_w13285_,
		_w13721_
	);
	LUT4 #(
		.INIT('h007d)
	) name13688 (
		_w6650_,
		_w13293_,
		_w13322_,
		_w13721_,
		_w13722_
	);
	LUT3 #(
		.INIT('h70)
	) name13689 (
		_w6657_,
		_w13716_,
		_w13722_,
		_w13723_
	);
	LUT4 #(
		.INIT('h95aa)
	) name13690 (
		\a[2] ,
		_w6335_,
		_w13720_,
		_w13723_,
		_w13724_
	);
	LUT2 #(
		.INIT('h2)
	) name13691 (
		_w13691_,
		_w13724_,
		_w13725_
	);
	LUT2 #(
		.INIT('h4)
	) name13692 (
		_w13691_,
		_w13724_,
		_w13726_
	);
	LUT2 #(
		.INIT('h9)
	) name13693 (
		_w13691_,
		_w13724_,
		_w13727_
	);
	LUT4 #(
		.INIT('h1501)
	) name13694 (
		_w13334_,
		_w13335_,
		_w13581_,
		_w13589_,
		_w13728_
	);
	LUT4 #(
		.INIT('h4920)
	) name13695 (
		_w13201_,
		_w13332_,
		_w13590_,
		_w13727_,
		_w13729_
	);
	LUT4 #(
		.INIT('h1e2d)
	) name13696 (
		_w13333_,
		_w13591_,
		_w13727_,
		_w13728_,
		_w13730_
	);
	LUT4 #(
		.INIT('h0f01)
	) name13697 (
		_w13333_,
		_w13591_,
		_w13725_,
		_w13726_,
		_w13731_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13698 (
		_w35_,
		_w13288_,
		_w13290_,
		_w13291_,
		_w13732_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13699 (
		_w6324_,
		_w13243_,
		_w13245_,
		_w13285_,
		_w13733_
	);
	LUT3 #(
		.INIT('h82)
	) name13700 (
		_w5524_,
		_w13062_,
		_w13099_,
		_w13734_
	);
	LUT3 #(
		.INIT('h07)
	) name13701 (
		_w6031_,
		_w13247_,
		_w13734_,
		_w13735_
	);
	LUT2 #(
		.INIT('h4)
	) name13702 (
		_w13733_,
		_w13735_,
		_w13736_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13703 (
		_w4459_,
		_w11384_,
		_w11488_,
		_w11489_,
		_w13737_
	);
	LUT4 #(
		.INIT('h2228)
	) name13704 (
		_w4700_,
		_w7695_,
		_w7750_,
		_w11285_,
		_w13738_
	);
	LUT3 #(
		.INIT('h82)
	) name13705 (
		_w4458_,
		_w11280_,
		_w11282_,
		_w13739_
	);
	LUT3 #(
		.INIT('h07)
	) name13706 (
		_w4684_,
		_w11382_,
		_w13739_,
		_w13740_
	);
	LUT2 #(
		.INIT('h4)
	) name13707 (
		_w13738_,
		_w13740_,
		_w13741_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13708 (
		_w3710_,
		_w11396_,
		_w11476_,
		_w11477_,
		_w13742_
	);
	LUT4 #(
		.INIT('h2228)
	) name13709 (
		_w3886_,
		_w8466_,
		_w8541_,
		_w11273_,
		_w13743_
	);
	LUT3 #(
		.INIT('h82)
	) name13710 (
		_w3709_,
		_w11268_,
		_w11270_,
		_w13744_
	);
	LUT3 #(
		.INIT('h07)
	) name13711 (
		_w3877_,
		_w11394_,
		_w13744_,
		_w13745_
	);
	LUT2 #(
		.INIT('h4)
	) name13712 (
		_w13743_,
		_w13745_,
		_w13746_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13713 (
		_w37_,
		_w11408_,
		_w11463_,
		_w11464_,
		_w13747_
	);
	LUT4 #(
		.INIT('h2228)
	) name13714 (
		_w3262_,
		_w9446_,
		_w9702_,
		_w11261_,
		_w13748_
	);
	LUT3 #(
		.INIT('h82)
	) name13715 (
		_w3214_,
		_w11256_,
		_w11258_,
		_w13749_
	);
	LUT3 #(
		.INIT('h07)
	) name13716 (
		_w3249_,
		_w11406_,
		_w13749_,
		_w13750_
	);
	LUT2 #(
		.INIT('h4)
	) name13717 (
		_w13748_,
		_w13750_,
		_w13751_
	);
	LUT3 #(
		.INIT('h32)
	) name13718 (
		_w13615_,
		_w13648_,
		_w13649_,
		_w13752_
	);
	LUT4 #(
		.INIT('h010f)
	) name13719 (
		_w13150_,
		_w13152_,
		_w13641_,
		_w13642_,
		_w13753_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13720 (
		_w2549_,
		_w10945_,
		_w11246_,
		_w11248_,
		_w13754_
	);
	LUT4 #(
		.INIT('h007d)
	) name13721 (
		_w2617_,
		_w11249_,
		_w11251_,
		_w13754_,
		_w13755_
	);
	LUT3 #(
		.INIT('h70)
	) name13722 (
		_w2854_,
		_w11415_,
		_w13755_,
		_w13756_
	);
	LUT4 #(
		.INIT('h95aa)
	) name13723 (
		\a[29] ,
		_w2550_,
		_w11675_,
		_w13756_,
		_w13757_
	);
	LUT4 #(
		.INIT('h135f)
	) name13724 (
		_w106_,
		_w90_,
		_w65_,
		_w236_,
		_w13758_
	);
	LUT4 #(
		.INIT('h8000)
	) name13725 (
		_w292_,
		_w1575_,
		_w1624_,
		_w13758_,
		_w13759_
	);
	LUT4 #(
		.INIT('h135f)
	) name13726 (
		_w55_,
		_w65_,
		_w236_,
		_w176_,
		_w13760_
	);
	LUT4 #(
		.INIT('h2000)
	) name13727 (
		_w132_,
		_w334_,
		_w797_,
		_w13760_,
		_w13761_
	);
	LUT3 #(
		.INIT('h80)
	) name13728 (
		_w4183_,
		_w13759_,
		_w13761_,
		_w13762_
	);
	LUT2 #(
		.INIT('h8)
	) name13729 (
		_w738_,
		_w3561_,
		_w13763_
	);
	LUT4 #(
		.INIT('h4000)
	) name13730 (
		_w141_,
		_w1472_,
		_w1865_,
		_w1866_,
		_w13764_
	);
	LUT4 #(
		.INIT('h8000)
	) name13731 (
		_w4245_,
		_w4246_,
		_w13763_,
		_w13764_,
		_w13765_
	);
	LUT4 #(
		.INIT('h8000)
	) name13732 (
		_w2085_,
		_w7612_,
		_w13762_,
		_w13765_,
		_w13766_
	);
	LUT2 #(
		.INIT('h8)
	) name13733 (
		_w871_,
		_w13766_,
		_w13767_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13734 (
		_w376_,
		_w10968_,
		_w11238_,
		_w11240_,
		_w13768_
	);
	LUT4 #(
		.INIT('h007d)
	) name13735 (
		_w2407_,
		_w11241_,
		_w11243_,
		_w13768_,
		_w13769_
	);
	LUT3 #(
		.INIT('h70)
	) name13736 (
		_w2527_,
		_w11421_,
		_w13769_,
		_w13770_
	);
	LUT4 #(
		.INIT('h080f)
	) name13737 (
		_w377_,
		_w11569_,
		_w13767_,
		_w13770_,
		_w13771_
	);
	LUT4 #(
		.INIT('h87f0)
	) name13738 (
		_w377_,
		_w11569_,
		_w13767_,
		_w13770_,
		_w13772_
	);
	LUT4 #(
		.INIT('h1700)
	) name13739 (
		_w13622_,
		_w13629_,
		_w13636_,
		_w13772_,
		_w13773_
	);
	LUT4 #(
		.INIT('h32cd)
	) name13740 (
		_w13622_,
		_w13637_,
		_w13638_,
		_w13772_,
		_w13774_
	);
	LUT2 #(
		.INIT('h4)
	) name13741 (
		_w13757_,
		_w13774_,
		_w13775_
	);
	LUT2 #(
		.INIT('h2)
	) name13742 (
		_w13757_,
		_w13774_,
		_w13776_
	);
	LUT2 #(
		.INIT('h9)
	) name13743 (
		_w13757_,
		_w13774_,
		_w13777_
	);
	LUT2 #(
		.INIT('h9)
	) name13744 (
		_w13753_,
		_w13777_,
		_w13778_
	);
	LUT3 #(
		.INIT('h82)
	) name13745 (
		_w2874_,
		_w10599_,
		_w11253_,
		_w13779_
	);
	LUT4 #(
		.INIT('h007d)
	) name13746 (
		_w2975_,
		_w10580_,
		_w11254_,
		_w13779_,
		_w13780_
	);
	LUT4 #(
		.INIT('h7d00)
	) name13747 (
		_w2986_,
		_w10268_,
		_w11255_,
		_w13780_,
		_w13781_
	);
	LUT4 #(
		.INIT('h7d00)
	) name13748 (
		_w2875_,
		_w11456_,
		_w11458_,
		_w13781_,
		_w13782_
	);
	LUT3 #(
		.INIT('h84)
	) name13749 (
		\a[26] ,
		_w13778_,
		_w13782_,
		_w13783_
	);
	LUT3 #(
		.INIT('h12)
	) name13750 (
		\a[26] ,
		_w13778_,
		_w13782_,
		_w13784_
	);
	LUT3 #(
		.INIT('h69)
	) name13751 (
		\a[26] ,
		_w13778_,
		_w13782_,
		_w13785_
	);
	LUT2 #(
		.INIT('h9)
	) name13752 (
		_w13752_,
		_w13785_,
		_w13786_
	);
	LUT4 #(
		.INIT('h6500)
	) name13753 (
		\a[23] ,
		_w13747_,
		_w13751_,
		_w13786_,
		_w13787_
	);
	LUT4 #(
		.INIT('h9a65)
	) name13754 (
		\a[23] ,
		_w13747_,
		_w13751_,
		_w13786_,
		_w13788_
	);
	LUT4 #(
		.INIT('h7100)
	) name13755 (
		_w13610_,
		_w13614_,
		_w13651_,
		_w13788_,
		_w13789_
	);
	LUT4 #(
		.INIT('h32cd)
	) name13756 (
		_w13610_,
		_w13652_,
		_w13653_,
		_w13788_,
		_w13790_
	);
	LUT3 #(
		.INIT('h82)
	) name13757 (
		_w3312_,
		_w11469_,
		_w11471_,
		_w13791_
	);
	LUT4 #(
		.INIT('h2228)
	) name13758 (
		_w3654_,
		_w8794_,
		_w8994_,
		_w11267_,
		_w13792_
	);
	LUT3 #(
		.INIT('h82)
	) name13759 (
		_w3311_,
		_w11262_,
		_w11264_,
		_w13793_
	);
	LUT3 #(
		.INIT('h07)
	) name13760 (
		_w3645_,
		_w11400_,
		_w13793_,
		_w13794_
	);
	LUT2 #(
		.INIT('h4)
	) name13761 (
		_w13792_,
		_w13794_,
		_w13795_
	);
	LUT4 #(
		.INIT('h4844)
	) name13762 (
		\a[20] ,
		_w13790_,
		_w13791_,
		_w13795_,
		_w13796_
	);
	LUT4 #(
		.INIT('h9699)
	) name13763 (
		\a[20] ,
		_w13790_,
		_w13791_,
		_w13795_,
		_w13797_
	);
	LUT4 #(
		.INIT('h4d00)
	) name13764 (
		_w13609_,
		_w13655_,
		_w13659_,
		_w13797_,
		_w13798_
	);
	LUT4 #(
		.INIT('h32cd)
	) name13765 (
		_w13609_,
		_w13660_,
		_w13661_,
		_w13797_,
		_w13799_
	);
	LUT4 #(
		.INIT('h6500)
	) name13766 (
		\a[17] ,
		_w13742_,
		_w13746_,
		_w13799_,
		_w13800_
	);
	LUT4 #(
		.INIT('h9a65)
	) name13767 (
		\a[17] ,
		_w13742_,
		_w13746_,
		_w13799_,
		_w13801_
	);
	LUT4 #(
		.INIT('h7100)
	) name13768 (
		_w13604_,
		_w13608_,
		_w13663_,
		_w13801_,
		_w13802_
	);
	LUT4 #(
		.INIT('h32cd)
	) name13769 (
		_w13604_,
		_w13664_,
		_w13665_,
		_w13801_,
		_w13803_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13770 (
		_w4034_,
		_w11390_,
		_w11482_,
		_w11483_,
		_w13804_
	);
	LUT4 #(
		.INIT('h2228)
	) name13771 (
		_w4382_,
		_w7935_,
		_w8077_,
		_w11279_,
		_w13805_
	);
	LUT3 #(
		.INIT('h82)
	) name13772 (
		_w4033_,
		_w11274_,
		_w11276_,
		_w13806_
	);
	LUT3 #(
		.INIT('h07)
	) name13773 (
		_w4367_,
		_w11388_,
		_w13806_,
		_w13807_
	);
	LUT2 #(
		.INIT('h4)
	) name13774 (
		_w13805_,
		_w13807_,
		_w13808_
	);
	LUT4 #(
		.INIT('h4844)
	) name13775 (
		\a[14] ,
		_w13803_,
		_w13804_,
		_w13808_,
		_w13809_
	);
	LUT4 #(
		.INIT('h9699)
	) name13776 (
		\a[14] ,
		_w13803_,
		_w13804_,
		_w13808_,
		_w13810_
	);
	LUT4 #(
		.INIT('h4d00)
	) name13777 (
		_w13603_,
		_w13667_,
		_w13671_,
		_w13810_,
		_w13811_
	);
	LUT4 #(
		.INIT('h32cd)
	) name13778 (
		_w13603_,
		_w13672_,
		_w13673_,
		_w13810_,
		_w13812_
	);
	LUT4 #(
		.INIT('h6500)
	) name13779 (
		\a[11] ,
		_w13737_,
		_w13741_,
		_w13812_,
		_w13813_
	);
	LUT4 #(
		.INIT('h9a65)
	) name13780 (
		\a[11] ,
		_w13737_,
		_w13741_,
		_w13812_,
		_w13814_
	);
	LUT4 #(
		.INIT('h7100)
	) name13781 (
		_w13598_,
		_w13602_,
		_w13675_,
		_w13814_,
		_w13815_
	);
	LUT4 #(
		.INIT('h32cd)
	) name13782 (
		_w13598_,
		_w13676_,
		_w13677_,
		_w13814_,
		_w13816_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13783 (
		_w4876_,
		_w11378_,
		_w11494_,
		_w11552_,
		_w13817_
	);
	LUT4 #(
		.INIT('h2228)
	) name13784 (
		_w5286_,
		_w11549_,
		_w11373_,
		_w11375_,
		_w13818_
	);
	LUT3 #(
		.INIT('h82)
	) name13785 (
		_w4875_,
		_w11286_,
		_w11335_,
		_w13819_
	);
	LUT3 #(
		.INIT('h07)
	) name13786 (
		_w5271_,
		_w11377_,
		_w13819_,
		_w13820_
	);
	LUT2 #(
		.INIT('h4)
	) name13787 (
		_w13818_,
		_w13820_,
		_w13821_
	);
	LUT4 #(
		.INIT('h4844)
	) name13788 (
		\a[8] ,
		_w13816_,
		_w13817_,
		_w13821_,
		_w13822_
	);
	LUT4 #(
		.INIT('h9699)
	) name13789 (
		\a[8] ,
		_w13816_,
		_w13817_,
		_w13821_,
		_w13823_
	);
	LUT4 #(
		.INIT('h4d00)
	) name13790 (
		_w13597_,
		_w13679_,
		_w13683_,
		_w13823_,
		_w13824_
	);
	LUT4 #(
		.INIT('h32cd)
	) name13791 (
		_w13597_,
		_w13684_,
		_w13685_,
		_w13823_,
		_w13825_
	);
	LUT4 #(
		.INIT('h6500)
	) name13792 (
		\a[5] ,
		_w13732_,
		_w13736_,
		_w13825_,
		_w13826_
	);
	LUT4 #(
		.INIT('h9a65)
	) name13793 (
		\a[5] ,
		_w13732_,
		_w13736_,
		_w13825_,
		_w13827_
	);
	LUT4 #(
		.INIT('h7100)
	) name13794 (
		_w13592_,
		_w13596_,
		_w13687_,
		_w13827_,
		_w13828_
	);
	LUT4 #(
		.INIT('h32cd)
	) name13795 (
		_w13592_,
		_w13688_,
		_w13689_,
		_w13827_,
		_w13829_
	);
	LUT2 #(
		.INIT('h8)
	) name13796 (
		_w121_,
		_w352_,
		_w13830_
	);
	LUT4 #(
		.INIT('h817e)
	) name13797 (
		_w13693_,
		_w13695_,
		_w13702_,
		_w13830_,
		_w13831_
	);
	LUT4 #(
		.INIT('h028a)
	) name13798 (
		_w2549_,
		_w7136_,
		_w7166_,
		_w7167_,
		_w13832_
	);
	LUT4 #(
		.INIT('h781e)
	) name13799 (
		\a[26] ,
		\a[27] ,
		\a[28] ,
		\a[29] ,
		_w13833_
	);
	LUT3 #(
		.INIT('hb0)
	) name13800 (
		_w7136_,
		_w7166_,
		_w13833_,
		_w13834_
	);
	LUT2 #(
		.INIT('h1)
	) name13801 (
		_w13832_,
		_w13834_,
		_w13835_
	);
	LUT4 #(
		.INIT('h5700)
	) name13802 (
		_w2550_,
		_w7418_,
		_w7419_,
		_w13835_,
		_w13836_
	);
	LUT3 #(
		.INIT('h82)
	) name13803 (
		_w377_,
		_w7135_,
		_w7172_,
		_w13837_
	);
	LUT3 #(
		.INIT('h28)
	) name13804 (
		_w2527_,
		_w7136_,
		_w7168_,
		_w13838_
	);
	LUT2 #(
		.INIT('h8)
	) name13805 (
		_w376_,
		_w6996_,
		_w13839_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13806 (
		_w2407_,
		_w2411_,
		_w6983_,
		_w6993_,
		_w13840_
	);
	LUT2 #(
		.INIT('h1)
	) name13807 (
		_w13839_,
		_w13840_,
		_w13841_
	);
	LUT2 #(
		.INIT('h4)
	) name13808 (
		_w13838_,
		_w13841_,
		_w13842_
	);
	LUT2 #(
		.INIT('h4)
	) name13809 (
		_w13837_,
		_w13842_,
		_w13843_
	);
	LUT4 #(
		.INIT('h6996)
	) name13810 (
		\a[29] ,
		_w13831_,
		_w13836_,
		_w13843_,
		_w13844_
	);
	LUT3 #(
		.INIT('he0)
	) name13811 (
		_w13704_,
		_w13710_,
		_w13844_,
		_w13845_
	);
	LUT3 #(
		.INIT('h01)
	) name13812 (
		_w13704_,
		_w13710_,
		_w13844_,
		_w13846_
	);
	LUT3 #(
		.INIT('h1e)
	) name13813 (
		_w13704_,
		_w13710_,
		_w13844_,
		_w13847_
	);
	LUT3 #(
		.INIT('h1e)
	) name13814 (
		_w13712_,
		_w13714_,
		_w13847_,
		_w13848_
	);
	LUT4 #(
		.INIT('h10e0)
	) name13815 (
		_w13712_,
		_w13714_,
		_w13716_,
		_w13847_,
		_w13849_
	);
	LUT4 #(
		.INIT('h12ed)
	) name13816 (
		_w13712_,
		_w13714_,
		_w13715_,
		_w13847_,
		_w13850_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13817 (
		_w6335_,
		_w13717_,
		_w13719_,
		_w13850_,
		_w13851_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13818 (
		_w6657_,
		_w13712_,
		_w13714_,
		_w13847_,
		_w13852_
	);
	LUT3 #(
		.INIT('h82)
	) name13819 (
		_w6334_,
		_w13293_,
		_w13322_,
		_w13853_
	);
	LUT3 #(
		.INIT('h07)
	) name13820 (
		_w6650_,
		_w13716_,
		_w13853_,
		_w13854_
	);
	LUT2 #(
		.INIT('h4)
	) name13821 (
		_w13852_,
		_w13854_,
		_w13855_
	);
	LUT3 #(
		.INIT('h9a)
	) name13822 (
		\a[2] ,
		_w13851_,
		_w13855_,
		_w13856_
	);
	LUT4 #(
		.INIT('h4844)
	) name13823 (
		\a[2] ,
		_w13829_,
		_w13851_,
		_w13855_,
		_w13857_
	);
	LUT4 #(
		.INIT('h2122)
	) name13824 (
		\a[2] ,
		_w13829_,
		_w13851_,
		_w13855_,
		_w13858_
	);
	LUT4 #(
		.INIT('h9699)
	) name13825 (
		\a[2] ,
		_w13829_,
		_w13851_,
		_w13855_,
		_w13859_
	);
	LUT3 #(
		.INIT('h82)
	) name13826 (
		_w13729_,
		_w13731_,
		_w13859_,
		_w13860_
	);
	LUT3 #(
		.INIT('h69)
	) name13827 (
		_w13729_,
		_w13731_,
		_w13859_,
		_w13861_
	);
	LUT3 #(
		.INIT('h82)
	) name13828 (
		_w35_,
		_w13292_,
		_w13325_,
		_w13862_
	);
	LUT3 #(
		.INIT('h82)
	) name13829 (
		_w6324_,
		_w13293_,
		_w13322_,
		_w13863_
	);
	LUT2 #(
		.INIT('h8)
	) name13830 (
		_w5524_,
		_w13247_,
		_w13864_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13831 (
		_w6031_,
		_w13243_,
		_w13245_,
		_w13285_,
		_w13865_
	);
	LUT2 #(
		.INIT('h1)
	) name13832 (
		_w13864_,
		_w13865_,
		_w13866_
	);
	LUT2 #(
		.INIT('h4)
	) name13833 (
		_w13863_,
		_w13866_,
		_w13867_
	);
	LUT3 #(
		.INIT('h82)
	) name13834 (
		_w4459_,
		_w11490_,
		_w11492_,
		_w13868_
	);
	LUT3 #(
		.INIT('h82)
	) name13835 (
		_w4700_,
		_w11286_,
		_w11335_,
		_w13869_
	);
	LUT2 #(
		.INIT('h8)
	) name13836 (
		_w4458_,
		_w11382_,
		_w13870_
	);
	LUT4 #(
		.INIT('h2228)
	) name13837 (
		_w4684_,
		_w7695_,
		_w7750_,
		_w11285_,
		_w13871_
	);
	LUT2 #(
		.INIT('h1)
	) name13838 (
		_w13870_,
		_w13871_,
		_w13872_
	);
	LUT2 #(
		.INIT('h4)
	) name13839 (
		_w13869_,
		_w13872_,
		_w13873_
	);
	LUT3 #(
		.INIT('h82)
	) name13840 (
		_w3710_,
		_w11478_,
		_w11480_,
		_w13874_
	);
	LUT3 #(
		.INIT('h82)
	) name13841 (
		_w3886_,
		_w11274_,
		_w11276_,
		_w13875_
	);
	LUT2 #(
		.INIT('h8)
	) name13842 (
		_w3709_,
		_w11394_,
		_w13876_
	);
	LUT4 #(
		.INIT('h2228)
	) name13843 (
		_w3877_,
		_w8466_,
		_w8541_,
		_w11273_,
		_w13877_
	);
	LUT2 #(
		.INIT('h1)
	) name13844 (
		_w13876_,
		_w13877_,
		_w13878_
	);
	LUT2 #(
		.INIT('h4)
	) name13845 (
		_w13875_,
		_w13878_,
		_w13879_
	);
	LUT3 #(
		.INIT('h82)
	) name13846 (
		_w37_,
		_w11465_,
		_w11467_,
		_w13880_
	);
	LUT3 #(
		.INIT('h82)
	) name13847 (
		_w3262_,
		_w11262_,
		_w11264_,
		_w13881_
	);
	LUT2 #(
		.INIT('h8)
	) name13848 (
		_w3214_,
		_w11406_,
		_w13882_
	);
	LUT4 #(
		.INIT('h2228)
	) name13849 (
		_w3249_,
		_w9446_,
		_w9702_,
		_w11261_,
		_w13883_
	);
	LUT2 #(
		.INIT('h1)
	) name13850 (
		_w13882_,
		_w13883_,
		_w13884_
	);
	LUT2 #(
		.INIT('h4)
	) name13851 (
		_w13881_,
		_w13884_,
		_w13885_
	);
	LUT3 #(
		.INIT('h32)
	) name13852 (
		_w13752_,
		_w13783_,
		_w13784_,
		_w13886_
	);
	LUT3 #(
		.INIT('h32)
	) name13853 (
		_w13753_,
		_w13775_,
		_w13776_,
		_w13887_
	);
	LUT3 #(
		.INIT('h82)
	) name13854 (
		_w2549_,
		_w11249_,
		_w11251_,
		_w13888_
	);
	LUT3 #(
		.INIT('h07)
	) name13855 (
		_w2617_,
		_w11415_,
		_w13888_,
		_w13889_
	);
	LUT4 #(
		.INIT('h7d00)
	) name13856 (
		_w2854_,
		_w10599_,
		_w11253_,
		_w13889_,
		_w13890_
	);
	LUT4 #(
		.INIT('h7d00)
	) name13857 (
		_w2550_,
		_w11450_,
		_w11452_,
		_w13890_,
		_w13891_
	);
	LUT4 #(
		.INIT('h8000)
	) name13858 (
		_w514_,
		_w777_,
		_w2060_,
		_w7997_,
		_w13892_
	);
	LUT4 #(
		.INIT('h135f)
	) name13859 (
		_w55_,
		_w56_,
		_w43_,
		_w158_,
		_w13893_
	);
	LUT4 #(
		.INIT('h2000)
	) name13860 (
		_w168_,
		_w353_,
		_w538_,
		_w13893_,
		_w13894_
	);
	LUT4 #(
		.INIT('h8000)
	) name13861 (
		_w1737_,
		_w4286_,
		_w13892_,
		_w13894_,
		_w13895_
	);
	LUT4 #(
		.INIT('h4000)
	) name13862 (
		_w295_,
		_w650_,
		_w951_,
		_w1184_,
		_w13896_
	);
	LUT4 #(
		.INIT('h8000)
	) name13863 (
		_w2795_,
		_w2798_,
		_w7623_,
		_w13896_,
		_w13897_
	);
	LUT4 #(
		.INIT('h8000)
	) name13864 (
		_w1612_,
		_w1619_,
		_w13895_,
		_w13897_,
		_w13898_
	);
	LUT2 #(
		.INIT('h8)
	) name13865 (
		_w2814_,
		_w13898_,
		_w13899_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13866 (
		_w377_,
		_w11423_,
		_w11443_,
		_w11444_,
		_w13900_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13867 (
		_w2527_,
		_w10945_,
		_w11246_,
		_w11248_,
		_w13901_
	);
	LUT3 #(
		.INIT('h82)
	) name13868 (
		_w376_,
		_w11241_,
		_w11243_,
		_w13902_
	);
	LUT3 #(
		.INIT('h07)
	) name13869 (
		_w2407_,
		_w11421_,
		_w13902_,
		_w13903_
	);
	LUT2 #(
		.INIT('h4)
	) name13870 (
		_w13901_,
		_w13903_,
		_w13904_
	);
	LUT3 #(
		.INIT('h45)
	) name13871 (
		_w13899_,
		_w13900_,
		_w13904_,
		_w13905_
	);
	LUT3 #(
		.INIT('h9a)
	) name13872 (
		_w13899_,
		_w13900_,
		_w13904_,
		_w13906_
	);
	LUT3 #(
		.INIT('h1e)
	) name13873 (
		_w13771_,
		_w13773_,
		_w13906_,
		_w13907_
	);
	LUT3 #(
		.INIT('h90)
	) name13874 (
		\a[29] ,
		_w13891_,
		_w13907_,
		_w13908_
	);
	LUT3 #(
		.INIT('h06)
	) name13875 (
		\a[29] ,
		_w13891_,
		_w13907_,
		_w13909_
	);
	LUT3 #(
		.INIT('h69)
	) name13876 (
		\a[29] ,
		_w13891_,
		_w13907_,
		_w13910_
	);
	LUT2 #(
		.INIT('h9)
	) name13877 (
		_w13887_,
		_w13910_,
		_w13911_
	);
	LUT3 #(
		.INIT('h82)
	) name13878 (
		_w2874_,
		_w10580_,
		_w11254_,
		_w13912_
	);
	LUT4 #(
		.INIT('h007d)
	) name13879 (
		_w2975_,
		_w10268_,
		_w11255_,
		_w13912_,
		_w13913_
	);
	LUT4 #(
		.INIT('h7d00)
	) name13880 (
		_w2986_,
		_w11256_,
		_w11258_,
		_w13913_,
		_w13914_
	);
	LUT4 #(
		.INIT('h7d00)
	) name13881 (
		_w2875_,
		_w11459_,
		_w11461_,
		_w13914_,
		_w13915_
	);
	LUT3 #(
		.INIT('h84)
	) name13882 (
		\a[26] ,
		_w13911_,
		_w13915_,
		_w13916_
	);
	LUT3 #(
		.INIT('h12)
	) name13883 (
		\a[26] ,
		_w13911_,
		_w13915_,
		_w13917_
	);
	LUT3 #(
		.INIT('h69)
	) name13884 (
		\a[26] ,
		_w13911_,
		_w13915_,
		_w13918_
	);
	LUT2 #(
		.INIT('h9)
	) name13885 (
		_w13886_,
		_w13918_,
		_w13919_
	);
	LUT4 #(
		.INIT('h6500)
	) name13886 (
		\a[23] ,
		_w13880_,
		_w13885_,
		_w13919_,
		_w13920_
	);
	LUT4 #(
		.INIT('h9a65)
	) name13887 (
		\a[23] ,
		_w13880_,
		_w13885_,
		_w13919_,
		_w13921_
	);
	LUT3 #(
		.INIT('h1e)
	) name13888 (
		_w13787_,
		_w13789_,
		_w13921_,
		_w13922_
	);
	LUT3 #(
		.INIT('h82)
	) name13889 (
		_w3312_,
		_w11472_,
		_w11474_,
		_w13923_
	);
	LUT3 #(
		.INIT('h82)
	) name13890 (
		_w3654_,
		_w11268_,
		_w11270_,
		_w13924_
	);
	LUT2 #(
		.INIT('h8)
	) name13891 (
		_w3311_,
		_w11400_,
		_w13925_
	);
	LUT4 #(
		.INIT('h2228)
	) name13892 (
		_w3645_,
		_w8794_,
		_w8994_,
		_w11267_,
		_w13926_
	);
	LUT2 #(
		.INIT('h1)
	) name13893 (
		_w13925_,
		_w13926_,
		_w13927_
	);
	LUT2 #(
		.INIT('h4)
	) name13894 (
		_w13924_,
		_w13927_,
		_w13928_
	);
	LUT4 #(
		.INIT('h4844)
	) name13895 (
		\a[20] ,
		_w13922_,
		_w13923_,
		_w13928_,
		_w13929_
	);
	LUT4 #(
		.INIT('h9699)
	) name13896 (
		\a[20] ,
		_w13922_,
		_w13923_,
		_w13928_,
		_w13930_
	);
	LUT3 #(
		.INIT('h1e)
	) name13897 (
		_w13796_,
		_w13798_,
		_w13930_,
		_w13931_
	);
	LUT4 #(
		.INIT('h6500)
	) name13898 (
		\a[17] ,
		_w13874_,
		_w13879_,
		_w13931_,
		_w13932_
	);
	LUT4 #(
		.INIT('h9a65)
	) name13899 (
		\a[17] ,
		_w13874_,
		_w13879_,
		_w13931_,
		_w13933_
	);
	LUT3 #(
		.INIT('h1e)
	) name13900 (
		_w13800_,
		_w13802_,
		_w13933_,
		_w13934_
	);
	LUT3 #(
		.INIT('h82)
	) name13901 (
		_w4034_,
		_w11484_,
		_w11486_,
		_w13935_
	);
	LUT3 #(
		.INIT('h82)
	) name13902 (
		_w4382_,
		_w11280_,
		_w11282_,
		_w13936_
	);
	LUT2 #(
		.INIT('h8)
	) name13903 (
		_w4033_,
		_w11388_,
		_w13937_
	);
	LUT4 #(
		.INIT('h2228)
	) name13904 (
		_w4367_,
		_w7935_,
		_w8077_,
		_w11279_,
		_w13938_
	);
	LUT2 #(
		.INIT('h1)
	) name13905 (
		_w13937_,
		_w13938_,
		_w13939_
	);
	LUT2 #(
		.INIT('h4)
	) name13906 (
		_w13936_,
		_w13939_,
		_w13940_
	);
	LUT4 #(
		.INIT('h4844)
	) name13907 (
		\a[14] ,
		_w13934_,
		_w13935_,
		_w13940_,
		_w13941_
	);
	LUT4 #(
		.INIT('h9699)
	) name13908 (
		\a[14] ,
		_w13934_,
		_w13935_,
		_w13940_,
		_w13942_
	);
	LUT3 #(
		.INIT('h1e)
	) name13909 (
		_w13809_,
		_w13811_,
		_w13942_,
		_w13943_
	);
	LUT4 #(
		.INIT('h6500)
	) name13910 (
		\a[11] ,
		_w13868_,
		_w13873_,
		_w13943_,
		_w13944_
	);
	LUT4 #(
		.INIT('h9a65)
	) name13911 (
		\a[11] ,
		_w13868_,
		_w13873_,
		_w13943_,
		_w13945_
	);
	LUT3 #(
		.INIT('h1e)
	) name13912 (
		_w13813_,
		_w13815_,
		_w13945_,
		_w13946_
	);
	LUT3 #(
		.INIT('h82)
	) name13913 (
		_w4876_,
		_w13061_,
		_w13102_,
		_w13947_
	);
	LUT3 #(
		.INIT('h82)
	) name13914 (
		_w5286_,
		_w13062_,
		_w13099_,
		_w13948_
	);
	LUT2 #(
		.INIT('h8)
	) name13915 (
		_w4875_,
		_w11377_,
		_w13949_
	);
	LUT4 #(
		.INIT('h2228)
	) name13916 (
		_w5271_,
		_w11549_,
		_w11373_,
		_w11375_,
		_w13950_
	);
	LUT2 #(
		.INIT('h1)
	) name13917 (
		_w13949_,
		_w13950_,
		_w13951_
	);
	LUT2 #(
		.INIT('h4)
	) name13918 (
		_w13948_,
		_w13951_,
		_w13952_
	);
	LUT4 #(
		.INIT('h4844)
	) name13919 (
		\a[8] ,
		_w13946_,
		_w13947_,
		_w13952_,
		_w13953_
	);
	LUT4 #(
		.INIT('h9699)
	) name13920 (
		\a[8] ,
		_w13946_,
		_w13947_,
		_w13952_,
		_w13954_
	);
	LUT3 #(
		.INIT('h1e)
	) name13921 (
		_w13822_,
		_w13824_,
		_w13954_,
		_w13955_
	);
	LUT4 #(
		.INIT('h6500)
	) name13922 (
		\a[5] ,
		_w13862_,
		_w13867_,
		_w13955_,
		_w13956_
	);
	LUT4 #(
		.INIT('h9a65)
	) name13923 (
		\a[5] ,
		_w13862_,
		_w13867_,
		_w13955_,
		_w13957_
	);
	LUT3 #(
		.INIT('h1e)
	) name13924 (
		_w13826_,
		_w13828_,
		_w13957_,
		_w13958_
	);
	LUT4 #(
		.INIT('h010f)
	) name13925 (
		_w13717_,
		_w13719_,
		_w13849_,
		_w13850_,
		_w13959_
	);
	LUT4 #(
		.INIT('h0f01)
	) name13926 (
		_w13712_,
		_w13714_,
		_w13845_,
		_w13846_,
		_w13960_
	);
	LUT4 #(
		.INIT('h7b12)
	) name13927 (
		\a[29] ,
		_w13831_,
		_w13836_,
		_w13843_,
		_w13961_
	);
	LUT4 #(
		.INIT('h80fe)
	) name13928 (
		_w13693_,
		_w13695_,
		_w13702_,
		_w13830_,
		_w13962_
	);
	LUT4 #(
		.INIT('h8001)
	) name13929 (
		\a[26] ,
		\a[27] ,
		\a[28] ,
		\a[29] ,
		_w13963_
	);
	LUT4 #(
		.INIT('h559a)
	) name13930 (
		\a[29] ,
		_w7136_,
		_w7166_,
		_w13963_,
		_w13964_
	);
	LUT3 #(
		.INIT('h80)
	) name13931 (
		_w7148_,
		_w7162_,
		_w13830_,
		_w13965_
	);
	LUT3 #(
		.INIT('h07)
	) name13932 (
		_w7148_,
		_w7162_,
		_w13830_,
		_w13966_
	);
	LUT3 #(
		.INIT('h78)
	) name13933 (
		_w7148_,
		_w7162_,
		_w13830_,
		_w13967_
	);
	LUT2 #(
		.INIT('h6)
	) name13934 (
		_w13964_,
		_w13967_,
		_w13968_
	);
	LUT3 #(
		.INIT('h28)
	) name13935 (
		_w2407_,
		_w7136_,
		_w7168_,
		_w13969_
	);
	LUT4 #(
		.INIT('h028a)
	) name13936 (
		_w2527_,
		_w7136_,
		_w7166_,
		_w7167_,
		_w13970_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13937 (
		_w376_,
		_w2411_,
		_w6983_,
		_w6993_,
		_w13971_
	);
	LUT3 #(
		.INIT('h01)
	) name13938 (
		_w13970_,
		_w13971_,
		_w13969_,
		_w13972_
	);
	LUT4 #(
		.INIT('h80f0)
	) name13939 (
		_w377_,
		_w7696_,
		_w13968_,
		_w13972_,
		_w13973_
	);
	LUT4 #(
		.INIT('h0700)
	) name13940 (
		_w377_,
		_w7696_,
		_w13968_,
		_w13972_,
		_w13974_
	);
	LUT4 #(
		.INIT('h780f)
	) name13941 (
		_w377_,
		_w7696_,
		_w13968_,
		_w13972_,
		_w13975_
	);
	LUT2 #(
		.INIT('h9)
	) name13942 (
		_w13962_,
		_w13975_,
		_w13976_
	);
	LUT2 #(
		.INIT('h4)
	) name13943 (
		_w13961_,
		_w13976_,
		_w13977_
	);
	LUT2 #(
		.INIT('h2)
	) name13944 (
		_w13961_,
		_w13976_,
		_w13978_
	);
	LUT2 #(
		.INIT('h9)
	) name13945 (
		_w13961_,
		_w13976_,
		_w13979_
	);
	LUT3 #(
		.INIT('h14)
	) name13946 (
		_w13848_,
		_w13960_,
		_w13979_,
		_w13980_
	);
	LUT3 #(
		.INIT('h82)
	) name13947 (
		_w13848_,
		_w13960_,
		_w13979_,
		_w13981_
	);
	LUT3 #(
		.INIT('h69)
	) name13948 (
		_w13848_,
		_w13960_,
		_w13979_,
		_w13982_
	);
	LUT3 #(
		.INIT('h82)
	) name13949 (
		_w6335_,
		_w13959_,
		_w13982_,
		_w13983_
	);
	LUT3 #(
		.INIT('h82)
	) name13950 (
		_w6657_,
		_w13960_,
		_w13979_,
		_w13984_
	);
	LUT2 #(
		.INIT('h8)
	) name13951 (
		_w6334_,
		_w13716_,
		_w13985_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13952 (
		_w6650_,
		_w13712_,
		_w13714_,
		_w13847_,
		_w13986_
	);
	LUT2 #(
		.INIT('h1)
	) name13953 (
		_w13985_,
		_w13986_,
		_w13987_
	);
	LUT2 #(
		.INIT('h4)
	) name13954 (
		_w13984_,
		_w13987_,
		_w13988_
	);
	LUT4 #(
		.INIT('h4844)
	) name13955 (
		\a[2] ,
		_w13958_,
		_w13983_,
		_w13988_,
		_w13989_
	);
	LUT4 #(
		.INIT('h9699)
	) name13956 (
		\a[2] ,
		_w13958_,
		_w13983_,
		_w13988_,
		_w13990_
	);
	LUT4 #(
		.INIT('h4d00)
	) name13957 (
		_w13731_,
		_w13829_,
		_w13856_,
		_w13990_,
		_w13991_
	);
	LUT4 #(
		.INIT('h32cd)
	) name13958 (
		_w13731_,
		_w13857_,
		_w13858_,
		_w13990_,
		_w13992_
	);
	LUT2 #(
		.INIT('h8)
	) name13959 (
		_w13860_,
		_w13992_,
		_w13993_
	);
	LUT2 #(
		.INIT('h6)
	) name13960 (
		_w13860_,
		_w13992_,
		_w13994_
	);
	LUT4 #(
		.INIT('h010f)
	) name13961 (
		_w13826_,
		_w13828_,
		_w13956_,
		_w13957_,
		_w13995_
	);
	LUT4 #(
		.INIT('h02a8)
	) name13962 (
		_w5524_,
		_w13243_,
		_w13245_,
		_w13285_,
		_w13996_
	);
	LUT4 #(
		.INIT('h007d)
	) name13963 (
		_w6031_,
		_w13293_,
		_w13322_,
		_w13996_,
		_w13997_
	);
	LUT3 #(
		.INIT('h70)
	) name13964 (
		_w6324_,
		_w13716_,
		_w13997_,
		_w13998_
	);
	LUT4 #(
		.INIT('h95aa)
	) name13965 (
		\a[5] ,
		_w35_,
		_w13720_,
		_w13998_,
		_w13999_
	);
	LUT4 #(
		.INIT('h010f)
	) name13966 (
		_w13822_,
		_w13824_,
		_w13953_,
		_w13954_,
		_w14000_
	);
	LUT4 #(
		.INIT('h010f)
	) name13967 (
		_w13813_,
		_w13815_,
		_w13944_,
		_w13945_,
		_w14001_
	);
	LUT4 #(
		.INIT('h2228)
	) name13968 (
		_w4458_,
		_w7695_,
		_w7750_,
		_w11285_,
		_w14002_
	);
	LUT4 #(
		.INIT('h007d)
	) name13969 (
		_w4684_,
		_w11286_,
		_w11335_,
		_w14002_,
		_w14003_
	);
	LUT3 #(
		.INIT('h70)
	) name13970 (
		_w4700_,
		_w11377_,
		_w14003_,
		_w14004_
	);
	LUT4 #(
		.INIT('h95aa)
	) name13971 (
		\a[11] ,
		_w4459_,
		_w12799_,
		_w14004_,
		_w14005_
	);
	LUT4 #(
		.INIT('h010f)
	) name13972 (
		_w13809_,
		_w13811_,
		_w13941_,
		_w13942_,
		_w14006_
	);
	LUT4 #(
		.INIT('h010f)
	) name13973 (
		_w13800_,
		_w13802_,
		_w13932_,
		_w13933_,
		_w14007_
	);
	LUT4 #(
		.INIT('h2228)
	) name13974 (
		_w3709_,
		_w8466_,
		_w8541_,
		_w11273_,
		_w14008_
	);
	LUT4 #(
		.INIT('h007d)
	) name13975 (
		_w3877_,
		_w11274_,
		_w11276_,
		_w14008_,
		_w14009_
	);
	LUT3 #(
		.INIT('h70)
	) name13976 (
		_w3886_,
		_w11388_,
		_w14009_,
		_w14010_
	);
	LUT4 #(
		.INIT('h95aa)
	) name13977 (
		\a[17] ,
		_w3710_,
		_w12391_,
		_w14010_,
		_w14011_
	);
	LUT4 #(
		.INIT('h010f)
	) name13978 (
		_w13796_,
		_w13798_,
		_w13929_,
		_w13930_,
		_w14012_
	);
	LUT4 #(
		.INIT('h010f)
	) name13979 (
		_w13787_,
		_w13789_,
		_w13920_,
		_w13921_,
		_w14013_
	);
	LUT4 #(
		.INIT('h2228)
	) name13980 (
		_w3214_,
		_w9446_,
		_w9702_,
		_w11261_,
		_w14014_
	);
	LUT4 #(
		.INIT('h007d)
	) name13981 (
		_w3249_,
		_w11262_,
		_w11264_,
		_w14014_,
		_w14015_
	);
	LUT3 #(
		.INIT('h70)
	) name13982 (
		_w3262_,
		_w11400_,
		_w14015_,
		_w14016_
	);
	LUT4 #(
		.INIT('h95aa)
	) name13983 (
		\a[23] ,
		_w37_,
		_w11967_,
		_w14016_,
		_w14017_
	);
	LUT3 #(
		.INIT('h32)
	) name13984 (
		_w13886_,
		_w13916_,
		_w13917_,
		_w14018_
	);
	LUT3 #(
		.INIT('h32)
	) name13985 (
		_w13887_,
		_w13908_,
		_w13909_,
		_w14019_
	);
	LUT2 #(
		.INIT('h8)
	) name13986 (
		_w2549_,
		_w11415_,
		_w14020_
	);
	LUT4 #(
		.INIT('h007d)
	) name13987 (
		_w2617_,
		_w10599_,
		_w11253_,
		_w14020_,
		_w14021_
	);
	LUT4 #(
		.INIT('h7d00)
	) name13988 (
		_w2854_,
		_w10580_,
		_w11254_,
		_w14021_,
		_w14022_
	);
	LUT4 #(
		.INIT('h7d00)
	) name13989 (
		_w2550_,
		_w11453_,
		_w11455_,
		_w14022_,
		_w14023_
	);
	LUT4 #(
		.INIT('h010f)
	) name13990 (
		_w13771_,
		_w13773_,
		_w13905_,
		_w13906_,
		_w14024_
	);
	LUT4 #(
		.INIT('h153f)
	) name13991 (
		_w122_,
		_w67_,
		_w39_,
		_w46_,
		_w14025_
	);
	LUT4 #(
		.INIT('h8000)
	) name13992 (
		_w649_,
		_w1624_,
		_w1697_,
		_w14025_,
		_w14026_
	);
	LUT4 #(
		.INIT('h4000)
	) name13993 (
		_w369_,
		_w776_,
		_w1707_,
		_w3341_,
		_w14027_
	);
	LUT3 #(
		.INIT('h80)
	) name13994 (
		_w245_,
		_w760_,
		_w856_,
		_w14028_
	);
	LUT3 #(
		.INIT('h80)
	) name13995 (
		_w697_,
		_w1014_,
		_w2060_,
		_w14029_
	);
	LUT4 #(
		.INIT('h8000)
	) name13996 (
		_w14028_,
		_w14029_,
		_w14026_,
		_w14027_,
		_w14030_
	);
	LUT3 #(
		.INIT('h80)
	) name13997 (
		_w1955_,
		_w8190_,
		_w14030_,
		_w14031_
	);
	LUT4 #(
		.INIT('h8000)
	) name13998 (
		_w2674_,
		_w2677_,
		_w4279_,
		_w4288_,
		_w14032_
	);
	LUT2 #(
		.INIT('h8)
	) name13999 (
		_w14031_,
		_w14032_,
		_w14033_
	);
	LUT3 #(
		.INIT('h82)
	) name14000 (
		_w377_,
		_w11445_,
		_w11447_,
		_w14034_
	);
	LUT3 #(
		.INIT('h82)
	) name14001 (
		_w2527_,
		_w11249_,
		_w11251_,
		_w14035_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14002 (
		_w2407_,
		_w10945_,
		_w11246_,
		_w11248_,
		_w14036_
	);
	LUT2 #(
		.INIT('h8)
	) name14003 (
		_w376_,
		_w11421_,
		_w14037_
	);
	LUT2 #(
		.INIT('h1)
	) name14004 (
		_w14036_,
		_w14037_,
		_w14038_
	);
	LUT2 #(
		.INIT('h4)
	) name14005 (
		_w14035_,
		_w14038_,
		_w14039_
	);
	LUT2 #(
		.INIT('h4)
	) name14006 (
		_w14034_,
		_w14039_,
		_w14040_
	);
	LUT3 #(
		.INIT('h45)
	) name14007 (
		_w14033_,
		_w14034_,
		_w14039_,
		_w14041_
	);
	LUT3 #(
		.INIT('h20)
	) name14008 (
		_w14033_,
		_w14034_,
		_w14039_,
		_w14042_
	);
	LUT3 #(
		.INIT('h9a)
	) name14009 (
		_w14033_,
		_w14034_,
		_w14039_,
		_w14043_
	);
	LUT2 #(
		.INIT('h9)
	) name14010 (
		_w14024_,
		_w14043_,
		_w14044_
	);
	LUT3 #(
		.INIT('h90)
	) name14011 (
		\a[29] ,
		_w14023_,
		_w14044_,
		_w14045_
	);
	LUT3 #(
		.INIT('h06)
	) name14012 (
		\a[29] ,
		_w14023_,
		_w14044_,
		_w14046_
	);
	LUT3 #(
		.INIT('h69)
	) name14013 (
		\a[29] ,
		_w14023_,
		_w14044_,
		_w14047_
	);
	LUT2 #(
		.INIT('h9)
	) name14014 (
		_w14019_,
		_w14047_,
		_w14048_
	);
	LUT3 #(
		.INIT('h82)
	) name14015 (
		_w2874_,
		_w10268_,
		_w11255_,
		_w14049_
	);
	LUT4 #(
		.INIT('h007d)
	) name14016 (
		_w2975_,
		_w11256_,
		_w11258_,
		_w14049_,
		_w14050_
	);
	LUT3 #(
		.INIT('h70)
	) name14017 (
		_w2986_,
		_w11406_,
		_w14050_,
		_w14051_
	);
	LUT4 #(
		.INIT('h95aa)
	) name14018 (
		\a[26] ,
		_w2875_,
		_w11796_,
		_w14051_,
		_w14052_
	);
	LUT2 #(
		.INIT('h2)
	) name14019 (
		_w14048_,
		_w14052_,
		_w14053_
	);
	LUT2 #(
		.INIT('h4)
	) name14020 (
		_w14048_,
		_w14052_,
		_w14054_
	);
	LUT2 #(
		.INIT('h9)
	) name14021 (
		_w14048_,
		_w14052_,
		_w14055_
	);
	LUT2 #(
		.INIT('h9)
	) name14022 (
		_w14018_,
		_w14055_,
		_w14056_
	);
	LUT2 #(
		.INIT('h4)
	) name14023 (
		_w14017_,
		_w14056_,
		_w14057_
	);
	LUT2 #(
		.INIT('h2)
	) name14024 (
		_w14017_,
		_w14056_,
		_w14058_
	);
	LUT2 #(
		.INIT('h9)
	) name14025 (
		_w14017_,
		_w14056_,
		_w14059_
	);
	LUT2 #(
		.INIT('h9)
	) name14026 (
		_w14013_,
		_w14059_,
		_w14060_
	);
	LUT4 #(
		.INIT('h2228)
	) name14027 (
		_w3311_,
		_w8794_,
		_w8994_,
		_w11267_,
		_w14061_
	);
	LUT4 #(
		.INIT('h007d)
	) name14028 (
		_w3645_,
		_w11268_,
		_w11270_,
		_w14061_,
		_w14062_
	);
	LUT3 #(
		.INIT('h70)
	) name14029 (
		_w3654_,
		_w11394_,
		_w14062_,
		_w14063_
	);
	LUT4 #(
		.INIT('h95aa)
	) name14030 (
		\a[20] ,
		_w3312_,
		_w12209_,
		_w14063_,
		_w14064_
	);
	LUT2 #(
		.INIT('h2)
	) name14031 (
		_w14060_,
		_w14064_,
		_w14065_
	);
	LUT2 #(
		.INIT('h4)
	) name14032 (
		_w14060_,
		_w14064_,
		_w14066_
	);
	LUT2 #(
		.INIT('h9)
	) name14033 (
		_w14060_,
		_w14064_,
		_w14067_
	);
	LUT2 #(
		.INIT('h9)
	) name14034 (
		_w14012_,
		_w14067_,
		_w14068_
	);
	LUT2 #(
		.INIT('h4)
	) name14035 (
		_w14011_,
		_w14068_,
		_w14069_
	);
	LUT2 #(
		.INIT('h2)
	) name14036 (
		_w14011_,
		_w14068_,
		_w14070_
	);
	LUT2 #(
		.INIT('h9)
	) name14037 (
		_w14011_,
		_w14068_,
		_w14071_
	);
	LUT2 #(
		.INIT('h9)
	) name14038 (
		_w14007_,
		_w14071_,
		_w14072_
	);
	LUT4 #(
		.INIT('h2228)
	) name14039 (
		_w4033_,
		_w7935_,
		_w8077_,
		_w11279_,
		_w14073_
	);
	LUT4 #(
		.INIT('h007d)
	) name14040 (
		_w4367_,
		_w11280_,
		_w11282_,
		_w14073_,
		_w14074_
	);
	LUT3 #(
		.INIT('h70)
	) name14041 (
		_w4382_,
		_w11382_,
		_w14074_,
		_w14075_
	);
	LUT4 #(
		.INIT('h95aa)
	) name14042 (
		\a[14] ,
		_w4034_,
		_w12476_,
		_w14075_,
		_w14076_
	);
	LUT2 #(
		.INIT('h2)
	) name14043 (
		_w14072_,
		_w14076_,
		_w14077_
	);
	LUT2 #(
		.INIT('h4)
	) name14044 (
		_w14072_,
		_w14076_,
		_w14078_
	);
	LUT2 #(
		.INIT('h9)
	) name14045 (
		_w14072_,
		_w14076_,
		_w14079_
	);
	LUT2 #(
		.INIT('h9)
	) name14046 (
		_w14006_,
		_w14079_,
		_w14080_
	);
	LUT2 #(
		.INIT('h4)
	) name14047 (
		_w14005_,
		_w14080_,
		_w14081_
	);
	LUT2 #(
		.INIT('h2)
	) name14048 (
		_w14005_,
		_w14080_,
		_w14082_
	);
	LUT2 #(
		.INIT('h9)
	) name14049 (
		_w14005_,
		_w14080_,
		_w14083_
	);
	LUT2 #(
		.INIT('h9)
	) name14050 (
		_w14001_,
		_w14083_,
		_w14084_
	);
	LUT4 #(
		.INIT('h2228)
	) name14051 (
		_w4875_,
		_w11549_,
		_w11373_,
		_w11375_,
		_w14085_
	);
	LUT4 #(
		.INIT('h007d)
	) name14052 (
		_w5271_,
		_w13062_,
		_w13099_,
		_w14085_,
		_w14086_
	);
	LUT3 #(
		.INIT('h70)
	) name14053 (
		_w5286_,
		_w13247_,
		_w14086_,
		_w14087_
	);
	LUT4 #(
		.INIT('h95aa)
	) name14054 (
		\a[8] ,
		_w4876_,
		_w13576_,
		_w14087_,
		_w14088_
	);
	LUT2 #(
		.INIT('h2)
	) name14055 (
		_w14084_,
		_w14088_,
		_w14089_
	);
	LUT2 #(
		.INIT('h4)
	) name14056 (
		_w14084_,
		_w14088_,
		_w14090_
	);
	LUT2 #(
		.INIT('h9)
	) name14057 (
		_w14084_,
		_w14088_,
		_w14091_
	);
	LUT2 #(
		.INIT('h9)
	) name14058 (
		_w14000_,
		_w14091_,
		_w14092_
	);
	LUT2 #(
		.INIT('h4)
	) name14059 (
		_w13999_,
		_w14092_,
		_w14093_
	);
	LUT2 #(
		.INIT('h2)
	) name14060 (
		_w13999_,
		_w14092_,
		_w14094_
	);
	LUT2 #(
		.INIT('h9)
	) name14061 (
		_w13999_,
		_w14092_,
		_w14095_
	);
	LUT2 #(
		.INIT('h9)
	) name14062 (
		_w13995_,
		_w14095_,
		_w14096_
	);
	LUT3 #(
		.INIT('h32)
	) name14063 (
		_w13962_,
		_w13973_,
		_w13974_,
		_w14097_
	);
	LUT4 #(
		.INIT('h2a02)
	) name14064 (
		_w373_,
		_w7163_,
		_w13830_,
		_w13964_,
		_w14098_
	);
	LUT4 #(
		.INIT('h4054)
	) name14065 (
		_w373_,
		_w7163_,
		_w13830_,
		_w13964_,
		_w14099_
	);
	LUT4 #(
		.INIT('h55a6)
	) name14066 (
		_w373_,
		_w13964_,
		_w13965_,
		_w13966_,
		_w14100_
	);
	LUT4 #(
		.INIT('h0a02)
	) name14067 (
		_w377_,
		_w7169_,
		_w7419_,
		_w7686_,
		_w14101_
	);
	LUT3 #(
		.INIT('h28)
	) name14068 (
		_w376_,
		_w7136_,
		_w7168_,
		_w14102_
	);
	LUT3 #(
		.INIT('h40)
	) name14069 (
		_w2527_,
		_w7136_,
		_w7167_,
		_w14103_
	);
	LUT3 #(
		.INIT('he1)
	) name14070 (
		\a[29] ,
		\a[30] ,
		\a[31] ,
		_w14104_
	);
	LUT3 #(
		.INIT('h0b)
	) name14071 (
		_w7136_,
		_w7166_,
		_w14104_,
		_w14105_
	);
	LUT3 #(
		.INIT('h45)
	) name14072 (
		_w14102_,
		_w14103_,
		_w14105_,
		_w14106_
	);
	LUT3 #(
		.INIT('h65)
	) name14073 (
		_w14100_,
		_w14101_,
		_w14106_,
		_w14107_
	);
	LUT2 #(
		.INIT('h4)
	) name14074 (
		_w14097_,
		_w14107_,
		_w14108_
	);
	LUT2 #(
		.INIT('h9)
	) name14075 (
		_w14097_,
		_w14107_,
		_w14109_
	);
	LUT4 #(
		.INIT('h008e)
	) name14076 (
		_w13960_,
		_w13961_,
		_w13976_,
		_w14109_,
		_w14110_
	);
	LUT4 #(
		.INIT('h7100)
	) name14077 (
		_w13960_,
		_w13961_,
		_w13976_,
		_w14109_,
		_w14111_
	);
	LUT4 #(
		.INIT('h32cd)
	) name14078 (
		_w13960_,
		_w13977_,
		_w13978_,
		_w14109_,
		_w14112_
	);
	LUT4 #(
		.INIT('h1244)
	) name14079 (
		_w13960_,
		_w13977_,
		_w13978_,
		_w14109_,
		_w14113_
	);
	LUT4 #(
		.INIT('h8679)
	) name14080 (
		_w13960_,
		_w13977_,
		_w13979_,
		_w14109_,
		_w14114_
	);
	LUT4 #(
		.INIT('hdc00)
	) name14081 (
		_w13959_,
		_w13981_,
		_w13982_,
		_w14114_,
		_w14115_
	);
	LUT4 #(
		.INIT('h0ef1)
	) name14082 (
		_w13959_,
		_w13980_,
		_w13981_,
		_w14114_,
		_w14116_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14083 (
		_w6334_,
		_w13712_,
		_w13714_,
		_w13847_,
		_w14117_
	);
	LUT4 #(
		.INIT('h007d)
	) name14084 (
		_w6650_,
		_w13960_,
		_w13979_,
		_w14117_,
		_w14118_
	);
	LUT3 #(
		.INIT('h70)
	) name14085 (
		_w6657_,
		_w14112_,
		_w14118_,
		_w14119_
	);
	LUT4 #(
		.INIT('h95aa)
	) name14086 (
		\a[2] ,
		_w6335_,
		_w14116_,
		_w14119_,
		_w14120_
	);
	LUT2 #(
		.INIT('h2)
	) name14087 (
		_w14096_,
		_w14120_,
		_w14121_
	);
	LUT2 #(
		.INIT('h4)
	) name14088 (
		_w14096_,
		_w14120_,
		_w14122_
	);
	LUT2 #(
		.INIT('h9)
	) name14089 (
		_w14096_,
		_w14120_,
		_w14123_
	);
	LUT3 #(
		.INIT('h1e)
	) name14090 (
		_w13989_,
		_w13991_,
		_w14123_,
		_w14124_
	);
	LUT2 #(
		.INIT('h6)
	) name14091 (
		_w13993_,
		_w14124_,
		_w14125_
	);
	LUT4 #(
		.INIT('h0f01)
	) name14092 (
		_w13989_,
		_w13991_,
		_w14121_,
		_w14122_,
		_w14126_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14093 (
		_w35_,
		_w13717_,
		_w13719_,
		_w13850_,
		_w14127_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14094 (
		_w6324_,
		_w13712_,
		_w13714_,
		_w13847_,
		_w14128_
	);
	LUT3 #(
		.INIT('h82)
	) name14095 (
		_w5524_,
		_w13293_,
		_w13322_,
		_w14129_
	);
	LUT3 #(
		.INIT('h07)
	) name14096 (
		_w6031_,
		_w13716_,
		_w14129_,
		_w14130_
	);
	LUT2 #(
		.INIT('h4)
	) name14097 (
		_w14128_,
		_w14130_,
		_w14131_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14098 (
		_w4459_,
		_w11378_,
		_w11494_,
		_w11552_,
		_w14132_
	);
	LUT4 #(
		.INIT('h2228)
	) name14099 (
		_w4700_,
		_w11549_,
		_w11373_,
		_w11375_,
		_w14133_
	);
	LUT3 #(
		.INIT('h82)
	) name14100 (
		_w4458_,
		_w11286_,
		_w11335_,
		_w14134_
	);
	LUT3 #(
		.INIT('h07)
	) name14101 (
		_w4684_,
		_w11377_,
		_w14134_,
		_w14135_
	);
	LUT2 #(
		.INIT('h4)
	) name14102 (
		_w14133_,
		_w14135_,
		_w14136_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14103 (
		_w3710_,
		_w11390_,
		_w11482_,
		_w11483_,
		_w14137_
	);
	LUT4 #(
		.INIT('h2228)
	) name14104 (
		_w3886_,
		_w7935_,
		_w8077_,
		_w11279_,
		_w14138_
	);
	LUT3 #(
		.INIT('h82)
	) name14105 (
		_w3709_,
		_w11274_,
		_w11276_,
		_w14139_
	);
	LUT3 #(
		.INIT('h07)
	) name14106 (
		_w3877_,
		_w11388_,
		_w14139_,
		_w14140_
	);
	LUT2 #(
		.INIT('h4)
	) name14107 (
		_w14138_,
		_w14140_,
		_w14141_
	);
	LUT3 #(
		.INIT('h82)
	) name14108 (
		_w37_,
		_w11469_,
		_w11471_,
		_w14142_
	);
	LUT4 #(
		.INIT('h2228)
	) name14109 (
		_w3262_,
		_w8794_,
		_w8994_,
		_w11267_,
		_w14143_
	);
	LUT3 #(
		.INIT('h82)
	) name14110 (
		_w3214_,
		_w11262_,
		_w11264_,
		_w14144_
	);
	LUT3 #(
		.INIT('h07)
	) name14111 (
		_w3249_,
		_w11400_,
		_w14144_,
		_w14145_
	);
	LUT2 #(
		.INIT('h4)
	) name14112 (
		_w14143_,
		_w14145_,
		_w14146_
	);
	LUT3 #(
		.INIT('h32)
	) name14113 (
		_w14019_,
		_w14045_,
		_w14046_,
		_w14147_
	);
	LUT3 #(
		.INIT('h82)
	) name14114 (
		_w2549_,
		_w10599_,
		_w11253_,
		_w14148_
	);
	LUT4 #(
		.INIT('h007d)
	) name14115 (
		_w2617_,
		_w10580_,
		_w11254_,
		_w14148_,
		_w14149_
	);
	LUT4 #(
		.INIT('h7d00)
	) name14116 (
		_w2854_,
		_w10268_,
		_w11255_,
		_w14149_,
		_w14150_
	);
	LUT4 #(
		.INIT('h7d00)
	) name14117 (
		_w2550_,
		_w11456_,
		_w11458_,
		_w14150_,
		_w14151_
	);
	LUT3 #(
		.INIT('h80)
	) name14118 (
		_w3932_,
		_w7149_,
		_w7537_,
		_w14152_
	);
	LUT4 #(
		.INIT('h135f)
	) name14119 (
		_w55_,
		_w46_,
		_w184_,
		_w201_,
		_w14153_
	);
	LUT4 #(
		.INIT('h1000)
	) name14120 (
		_w146_,
		_w482_,
		_w868_,
		_w14153_,
		_w14154_
	);
	LUT3 #(
		.INIT('h80)
	) name14121 (
		_w13763_,
		_w14152_,
		_w14154_,
		_w14155_
	);
	LUT4 #(
		.INIT('h1000)
	) name14122 (
		_w114_,
		_w413_,
		_w714_,
		_w1362_,
		_w14156_
	);
	LUT4 #(
		.INIT('h8000)
	) name14123 (
		_w305_,
		_w609_,
		_w1463_,
		_w1464_,
		_w14157_
	);
	LUT2 #(
		.INIT('h8)
	) name14124 (
		_w14156_,
		_w14157_,
		_w14158_
	);
	LUT4 #(
		.INIT('h8000)
	) name14125 (
		_w780_,
		_w937_,
		_w1687_,
		_w1878_,
		_w14159_
	);
	LUT4 #(
		.INIT('h135f)
	) name14126 (
		_w122_,
		_w55_,
		_w93_,
		_w236_,
		_w14160_
	);
	LUT4 #(
		.INIT('h2000)
	) name14127 (
		_w48_,
		_w409_,
		_w806_,
		_w14160_,
		_w14161_
	);
	LUT3 #(
		.INIT('h80)
	) name14128 (
		_w1860_,
		_w14159_,
		_w14161_,
		_w14162_
	);
	LUT3 #(
		.INIT('h80)
	) name14129 (
		_w14155_,
		_w14158_,
		_w14162_,
		_w14163_
	);
	LUT3 #(
		.INIT('h80)
	) name14130 (
		_w2785_,
		_w3151_,
		_w14163_,
		_w14164_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14131 (
		_w376_,
		_w10945_,
		_w11246_,
		_w11248_,
		_w14165_
	);
	LUT4 #(
		.INIT('h007d)
	) name14132 (
		_w2407_,
		_w11249_,
		_w11251_,
		_w14165_,
		_w14166_
	);
	LUT3 #(
		.INIT('h70)
	) name14133 (
		_w2527_,
		_w11415_,
		_w14166_,
		_w14167_
	);
	LUT4 #(
		.INIT('h080f)
	) name14134 (
		_w377_,
		_w11675_,
		_w14164_,
		_w14167_,
		_w14168_
	);
	LUT4 #(
		.INIT('h87f0)
	) name14135 (
		_w377_,
		_w11675_,
		_w14164_,
		_w14167_,
		_w14169_
	);
	LUT4 #(
		.INIT('h1700)
	) name14136 (
		_w14024_,
		_w14033_,
		_w14040_,
		_w14169_,
		_w14170_
	);
	LUT4 #(
		.INIT('h32cd)
	) name14137 (
		_w14024_,
		_w14041_,
		_w14042_,
		_w14169_,
		_w14171_
	);
	LUT3 #(
		.INIT('h90)
	) name14138 (
		\a[29] ,
		_w14151_,
		_w14171_,
		_w14172_
	);
	LUT3 #(
		.INIT('h06)
	) name14139 (
		\a[29] ,
		_w14151_,
		_w14171_,
		_w14173_
	);
	LUT3 #(
		.INIT('h69)
	) name14140 (
		\a[29] ,
		_w14151_,
		_w14171_,
		_w14174_
	);
	LUT2 #(
		.INIT('h9)
	) name14141 (
		_w14147_,
		_w14174_,
		_w14175_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14142 (
		_w2875_,
		_w11408_,
		_w11463_,
		_w11464_,
		_w14176_
	);
	LUT4 #(
		.INIT('h2228)
	) name14143 (
		_w2986_,
		_w9446_,
		_w9702_,
		_w11261_,
		_w14177_
	);
	LUT3 #(
		.INIT('h82)
	) name14144 (
		_w2874_,
		_w11256_,
		_w11258_,
		_w14178_
	);
	LUT3 #(
		.INIT('h07)
	) name14145 (
		_w2975_,
		_w11406_,
		_w14178_,
		_w14179_
	);
	LUT2 #(
		.INIT('h4)
	) name14146 (
		_w14177_,
		_w14179_,
		_w14180_
	);
	LUT4 #(
		.INIT('h4844)
	) name14147 (
		\a[26] ,
		_w14175_,
		_w14176_,
		_w14180_,
		_w14181_
	);
	LUT4 #(
		.INIT('h9699)
	) name14148 (
		\a[26] ,
		_w14175_,
		_w14176_,
		_w14180_,
		_w14182_
	);
	LUT4 #(
		.INIT('h4d00)
	) name14149 (
		_w14018_,
		_w14048_,
		_w14052_,
		_w14182_,
		_w14183_
	);
	LUT4 #(
		.INIT('h32cd)
	) name14150 (
		_w14018_,
		_w14053_,
		_w14054_,
		_w14182_,
		_w14184_
	);
	LUT4 #(
		.INIT('h6500)
	) name14151 (
		\a[23] ,
		_w14142_,
		_w14146_,
		_w14184_,
		_w14185_
	);
	LUT4 #(
		.INIT('h9a65)
	) name14152 (
		\a[23] ,
		_w14142_,
		_w14146_,
		_w14184_,
		_w14186_
	);
	LUT4 #(
		.INIT('h7100)
	) name14153 (
		_w14013_,
		_w14017_,
		_w14056_,
		_w14186_,
		_w14187_
	);
	LUT4 #(
		.INIT('h32cd)
	) name14154 (
		_w14013_,
		_w14057_,
		_w14058_,
		_w14186_,
		_w14188_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14155 (
		_w3312_,
		_w11396_,
		_w11476_,
		_w11477_,
		_w14189_
	);
	LUT4 #(
		.INIT('h2228)
	) name14156 (
		_w3654_,
		_w8466_,
		_w8541_,
		_w11273_,
		_w14190_
	);
	LUT3 #(
		.INIT('h82)
	) name14157 (
		_w3311_,
		_w11268_,
		_w11270_,
		_w14191_
	);
	LUT3 #(
		.INIT('h07)
	) name14158 (
		_w3645_,
		_w11394_,
		_w14191_,
		_w14192_
	);
	LUT2 #(
		.INIT('h4)
	) name14159 (
		_w14190_,
		_w14192_,
		_w14193_
	);
	LUT4 #(
		.INIT('h4844)
	) name14160 (
		\a[20] ,
		_w14188_,
		_w14189_,
		_w14193_,
		_w14194_
	);
	LUT4 #(
		.INIT('h9699)
	) name14161 (
		\a[20] ,
		_w14188_,
		_w14189_,
		_w14193_,
		_w14195_
	);
	LUT4 #(
		.INIT('h4d00)
	) name14162 (
		_w14012_,
		_w14060_,
		_w14064_,
		_w14195_,
		_w14196_
	);
	LUT4 #(
		.INIT('h32cd)
	) name14163 (
		_w14012_,
		_w14065_,
		_w14066_,
		_w14195_,
		_w14197_
	);
	LUT4 #(
		.INIT('h6500)
	) name14164 (
		\a[17] ,
		_w14137_,
		_w14141_,
		_w14197_,
		_w14198_
	);
	LUT4 #(
		.INIT('h9a65)
	) name14165 (
		\a[17] ,
		_w14137_,
		_w14141_,
		_w14197_,
		_w14199_
	);
	LUT4 #(
		.INIT('h7100)
	) name14166 (
		_w14007_,
		_w14011_,
		_w14068_,
		_w14199_,
		_w14200_
	);
	LUT4 #(
		.INIT('h32cd)
	) name14167 (
		_w14007_,
		_w14069_,
		_w14070_,
		_w14199_,
		_w14201_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14168 (
		_w4034_,
		_w11384_,
		_w11488_,
		_w11489_,
		_w14202_
	);
	LUT4 #(
		.INIT('h2228)
	) name14169 (
		_w4382_,
		_w7695_,
		_w7750_,
		_w11285_,
		_w14203_
	);
	LUT3 #(
		.INIT('h82)
	) name14170 (
		_w4033_,
		_w11280_,
		_w11282_,
		_w14204_
	);
	LUT3 #(
		.INIT('h07)
	) name14171 (
		_w4367_,
		_w11382_,
		_w14204_,
		_w14205_
	);
	LUT2 #(
		.INIT('h4)
	) name14172 (
		_w14203_,
		_w14205_,
		_w14206_
	);
	LUT4 #(
		.INIT('h4844)
	) name14173 (
		\a[14] ,
		_w14201_,
		_w14202_,
		_w14206_,
		_w14207_
	);
	LUT4 #(
		.INIT('h9699)
	) name14174 (
		\a[14] ,
		_w14201_,
		_w14202_,
		_w14206_,
		_w14208_
	);
	LUT4 #(
		.INIT('h4d00)
	) name14175 (
		_w14006_,
		_w14072_,
		_w14076_,
		_w14208_,
		_w14209_
	);
	LUT4 #(
		.INIT('h32cd)
	) name14176 (
		_w14006_,
		_w14077_,
		_w14078_,
		_w14208_,
		_w14210_
	);
	LUT4 #(
		.INIT('h6500)
	) name14177 (
		\a[11] ,
		_w14132_,
		_w14136_,
		_w14210_,
		_w14211_
	);
	LUT4 #(
		.INIT('h9a65)
	) name14178 (
		\a[11] ,
		_w14132_,
		_w14136_,
		_w14210_,
		_w14212_
	);
	LUT4 #(
		.INIT('h7100)
	) name14179 (
		_w14001_,
		_w14005_,
		_w14080_,
		_w14212_,
		_w14213_
	);
	LUT4 #(
		.INIT('h32cd)
	) name14180 (
		_w14001_,
		_w14081_,
		_w14082_,
		_w14212_,
		_w14214_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14181 (
		_w4876_,
		_w13288_,
		_w13290_,
		_w13291_,
		_w14215_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14182 (
		_w5286_,
		_w13243_,
		_w13245_,
		_w13285_,
		_w14216_
	);
	LUT3 #(
		.INIT('h82)
	) name14183 (
		_w4875_,
		_w13062_,
		_w13099_,
		_w14217_
	);
	LUT3 #(
		.INIT('h07)
	) name14184 (
		_w5271_,
		_w13247_,
		_w14217_,
		_w14218_
	);
	LUT2 #(
		.INIT('h4)
	) name14185 (
		_w14216_,
		_w14218_,
		_w14219_
	);
	LUT4 #(
		.INIT('h4844)
	) name14186 (
		\a[8] ,
		_w14214_,
		_w14215_,
		_w14219_,
		_w14220_
	);
	LUT4 #(
		.INIT('h9699)
	) name14187 (
		\a[8] ,
		_w14214_,
		_w14215_,
		_w14219_,
		_w14221_
	);
	LUT4 #(
		.INIT('h4d00)
	) name14188 (
		_w14000_,
		_w14084_,
		_w14088_,
		_w14221_,
		_w14222_
	);
	LUT4 #(
		.INIT('h32cd)
	) name14189 (
		_w14000_,
		_w14089_,
		_w14090_,
		_w14221_,
		_w14223_
	);
	LUT4 #(
		.INIT('h6500)
	) name14190 (
		\a[5] ,
		_w14127_,
		_w14131_,
		_w14223_,
		_w14224_
	);
	LUT4 #(
		.INIT('h9a65)
	) name14191 (
		\a[5] ,
		_w14127_,
		_w14131_,
		_w14223_,
		_w14225_
	);
	LUT4 #(
		.INIT('h7100)
	) name14192 (
		_w13995_,
		_w13999_,
		_w14092_,
		_w14225_,
		_w14226_
	);
	LUT4 #(
		.INIT('h32cd)
	) name14193 (
		_w13995_,
		_w14093_,
		_w14094_,
		_w14225_,
		_w14227_
	);
	LUT4 #(
		.INIT('h028a)
	) name14194 (
		_w376_,
		_w7136_,
		_w7166_,
		_w7167_,
		_w14228_
	);
	LUT2 #(
		.INIT('h1)
	) name14195 (
		_w14105_,
		_w14228_,
		_w14229_
	);
	LUT4 #(
		.INIT('h5700)
	) name14196 (
		_w377_,
		_w7418_,
		_w7419_,
		_w14229_,
		_w14230_
	);
	LUT2 #(
		.INIT('h6)
	) name14197 (
		_w373_,
		_w14230_,
		_w14231_
	);
	LUT4 #(
		.INIT('h3233)
	) name14198 (
		_w14098_,
		_w14099_,
		_w14101_,
		_w14106_,
		_w14232_
	);
	LUT2 #(
		.INIT('h2)
	) name14199 (
		_w14231_,
		_w14232_,
		_w14233_
	);
	LUT2 #(
		.INIT('h4)
	) name14200 (
		_w14231_,
		_w14232_,
		_w14234_
	);
	LUT2 #(
		.INIT('h9)
	) name14201 (
		_w14231_,
		_w14232_,
		_w14235_
	);
	LUT3 #(
		.INIT('h1e)
	) name14202 (
		_w14108_,
		_w14111_,
		_w14235_,
		_w14236_
	);
	LUT4 #(
		.INIT('h10e0)
	) name14203 (
		_w14108_,
		_w14111_,
		_w14112_,
		_w14235_,
		_w14237_
	);
	LUT4 #(
		.INIT('h06f9)
	) name14204 (
		_w14108_,
		_w14110_,
		_w14111_,
		_w14235_,
		_w14238_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14205 (
		_w6335_,
		_w14113_,
		_w14115_,
		_w14238_,
		_w14239_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14206 (
		_w6657_,
		_w14108_,
		_w14111_,
		_w14235_,
		_w14240_
	);
	LUT3 #(
		.INIT('h82)
	) name14207 (
		_w6334_,
		_w13960_,
		_w13979_,
		_w14241_
	);
	LUT3 #(
		.INIT('h07)
	) name14208 (
		_w6650_,
		_w14112_,
		_w14241_,
		_w14242_
	);
	LUT2 #(
		.INIT('h4)
	) name14209 (
		_w14240_,
		_w14242_,
		_w14243_
	);
	LUT3 #(
		.INIT('h9a)
	) name14210 (
		\a[2] ,
		_w14239_,
		_w14243_,
		_w14244_
	);
	LUT4 #(
		.INIT('h4844)
	) name14211 (
		\a[2] ,
		_w14227_,
		_w14239_,
		_w14243_,
		_w14245_
	);
	LUT4 #(
		.INIT('h2122)
	) name14212 (
		\a[2] ,
		_w14227_,
		_w14239_,
		_w14243_,
		_w14246_
	);
	LUT4 #(
		.INIT('h9699)
	) name14213 (
		\a[2] ,
		_w14227_,
		_w14239_,
		_w14243_,
		_w14247_
	);
	LUT4 #(
		.INIT('h8008)
	) name14214 (
		_w13993_,
		_w14124_,
		_w14126_,
		_w14247_,
		_w14248_
	);
	LUT4 #(
		.INIT('h7887)
	) name14215 (
		_w13993_,
		_w14124_,
		_w14126_,
		_w14247_,
		_w14249_
	);
	LUT3 #(
		.INIT('h82)
	) name14216 (
		_w35_,
		_w13959_,
		_w13982_,
		_w14250_
	);
	LUT3 #(
		.INIT('h82)
	) name14217 (
		_w6324_,
		_w13960_,
		_w13979_,
		_w14251_
	);
	LUT2 #(
		.INIT('h8)
	) name14218 (
		_w5524_,
		_w13716_,
		_w14252_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14219 (
		_w6031_,
		_w13712_,
		_w13714_,
		_w13847_,
		_w14253_
	);
	LUT2 #(
		.INIT('h1)
	) name14220 (
		_w14252_,
		_w14253_,
		_w14254_
	);
	LUT2 #(
		.INIT('h4)
	) name14221 (
		_w14251_,
		_w14254_,
		_w14255_
	);
	LUT3 #(
		.INIT('h82)
	) name14222 (
		_w4459_,
		_w13061_,
		_w13102_,
		_w14256_
	);
	LUT3 #(
		.INIT('h82)
	) name14223 (
		_w4700_,
		_w13062_,
		_w13099_,
		_w14257_
	);
	LUT2 #(
		.INIT('h8)
	) name14224 (
		_w4458_,
		_w11377_,
		_w14258_
	);
	LUT4 #(
		.INIT('h2228)
	) name14225 (
		_w4684_,
		_w11549_,
		_w11373_,
		_w11375_,
		_w14259_
	);
	LUT2 #(
		.INIT('h1)
	) name14226 (
		_w14258_,
		_w14259_,
		_w14260_
	);
	LUT2 #(
		.INIT('h4)
	) name14227 (
		_w14257_,
		_w14260_,
		_w14261_
	);
	LUT3 #(
		.INIT('h82)
	) name14228 (
		_w3710_,
		_w11484_,
		_w11486_,
		_w14262_
	);
	LUT3 #(
		.INIT('h82)
	) name14229 (
		_w3886_,
		_w11280_,
		_w11282_,
		_w14263_
	);
	LUT2 #(
		.INIT('h8)
	) name14230 (
		_w3709_,
		_w11388_,
		_w14264_
	);
	LUT4 #(
		.INIT('h2228)
	) name14231 (
		_w3877_,
		_w7935_,
		_w8077_,
		_w11279_,
		_w14265_
	);
	LUT2 #(
		.INIT('h1)
	) name14232 (
		_w14264_,
		_w14265_,
		_w14266_
	);
	LUT2 #(
		.INIT('h4)
	) name14233 (
		_w14263_,
		_w14266_,
		_w14267_
	);
	LUT3 #(
		.INIT('h82)
	) name14234 (
		_w37_,
		_w11472_,
		_w11474_,
		_w14268_
	);
	LUT3 #(
		.INIT('h82)
	) name14235 (
		_w3262_,
		_w11268_,
		_w11270_,
		_w14269_
	);
	LUT2 #(
		.INIT('h8)
	) name14236 (
		_w3214_,
		_w11400_,
		_w14270_
	);
	LUT4 #(
		.INIT('h2228)
	) name14237 (
		_w3249_,
		_w8794_,
		_w8994_,
		_w11267_,
		_w14271_
	);
	LUT2 #(
		.INIT('h1)
	) name14238 (
		_w14270_,
		_w14271_,
		_w14272_
	);
	LUT2 #(
		.INIT('h4)
	) name14239 (
		_w14269_,
		_w14272_,
		_w14273_
	);
	LUT3 #(
		.INIT('h32)
	) name14240 (
		_w14147_,
		_w14172_,
		_w14173_,
		_w14274_
	);
	LUT3 #(
		.INIT('h82)
	) name14241 (
		_w2549_,
		_w10580_,
		_w11254_,
		_w14275_
	);
	LUT4 #(
		.INIT('h007d)
	) name14242 (
		_w2617_,
		_w10268_,
		_w11255_,
		_w14275_,
		_w14276_
	);
	LUT4 #(
		.INIT('h7d00)
	) name14243 (
		_w2854_,
		_w11256_,
		_w11258_,
		_w14276_,
		_w14277_
	);
	LUT4 #(
		.INIT('h7d00)
	) name14244 (
		_w2550_,
		_w11459_,
		_w11461_,
		_w14277_,
		_w14278_
	);
	LUT4 #(
		.INIT('h8000)
	) name14245 (
		_w750_,
		_w1631_,
		_w2451_,
		_w7337_,
		_w14279_
	);
	LUT3 #(
		.INIT('h80)
	) name14246 (
		_w699_,
		_w2680_,
		_w14279_,
		_w14280_
	);
	LUT4 #(
		.INIT('h135f)
	) name14247 (
		_w55_,
		_w52_,
		_w39_,
		_w176_,
		_w14281_
	);
	LUT4 #(
		.INIT('h0400)
	) name14248 (
		_w80_,
		_w348_,
		_w451_,
		_w14281_,
		_w14282_
	);
	LUT4 #(
		.INIT('h8000)
	) name14249 (
		_w2639_,
		_w2641_,
		_w3934_,
		_w14282_,
		_w14283_
	);
	LUT4 #(
		.INIT('h8000)
	) name14250 (
		_w3563_,
		_w3575_,
		_w14280_,
		_w14283_,
		_w14284_
	);
	LUT2 #(
		.INIT('h8)
	) name14251 (
		_w8314_,
		_w14284_,
		_w14285_
	);
	LUT3 #(
		.INIT('h82)
	) name14252 (
		_w376_,
		_w11249_,
		_w11251_,
		_w14286_
	);
	LUT3 #(
		.INIT('h07)
	) name14253 (
		_w2407_,
		_w11415_,
		_w14286_,
		_w14287_
	);
	LUT4 #(
		.INIT('h7d00)
	) name14254 (
		_w2527_,
		_w10599_,
		_w11253_,
		_w14287_,
		_w14288_
	);
	LUT4 #(
		.INIT('h7d00)
	) name14255 (
		_w377_,
		_w11450_,
		_w11452_,
		_w14288_,
		_w14289_
	);
	LUT4 #(
		.INIT('he11e)
	) name14256 (
		_w14168_,
		_w14170_,
		_w14285_,
		_w14289_,
		_w14290_
	);
	LUT3 #(
		.INIT('h90)
	) name14257 (
		\a[29] ,
		_w14278_,
		_w14290_,
		_w14291_
	);
	LUT3 #(
		.INIT('h06)
	) name14258 (
		\a[29] ,
		_w14278_,
		_w14290_,
		_w14292_
	);
	LUT3 #(
		.INIT('h69)
	) name14259 (
		\a[29] ,
		_w14278_,
		_w14290_,
		_w14293_
	);
	LUT2 #(
		.INIT('h9)
	) name14260 (
		_w14274_,
		_w14293_,
		_w14294_
	);
	LUT3 #(
		.INIT('h82)
	) name14261 (
		_w2875_,
		_w11465_,
		_w11467_,
		_w14295_
	);
	LUT3 #(
		.INIT('h82)
	) name14262 (
		_w2986_,
		_w11262_,
		_w11264_,
		_w14296_
	);
	LUT2 #(
		.INIT('h8)
	) name14263 (
		_w2874_,
		_w11406_,
		_w14297_
	);
	LUT4 #(
		.INIT('h2228)
	) name14264 (
		_w2975_,
		_w9446_,
		_w9702_,
		_w11261_,
		_w14298_
	);
	LUT2 #(
		.INIT('h1)
	) name14265 (
		_w14297_,
		_w14298_,
		_w14299_
	);
	LUT2 #(
		.INIT('h4)
	) name14266 (
		_w14296_,
		_w14299_,
		_w14300_
	);
	LUT4 #(
		.INIT('h4844)
	) name14267 (
		\a[26] ,
		_w14294_,
		_w14295_,
		_w14300_,
		_w14301_
	);
	LUT4 #(
		.INIT('h9699)
	) name14268 (
		\a[26] ,
		_w14294_,
		_w14295_,
		_w14300_,
		_w14302_
	);
	LUT3 #(
		.INIT('h1e)
	) name14269 (
		_w14181_,
		_w14183_,
		_w14302_,
		_w14303_
	);
	LUT4 #(
		.INIT('h6500)
	) name14270 (
		\a[23] ,
		_w14268_,
		_w14273_,
		_w14303_,
		_w14304_
	);
	LUT4 #(
		.INIT('h9a65)
	) name14271 (
		\a[23] ,
		_w14268_,
		_w14273_,
		_w14303_,
		_w14305_
	);
	LUT3 #(
		.INIT('h1e)
	) name14272 (
		_w14185_,
		_w14187_,
		_w14305_,
		_w14306_
	);
	LUT3 #(
		.INIT('h82)
	) name14273 (
		_w3312_,
		_w11478_,
		_w11480_,
		_w14307_
	);
	LUT3 #(
		.INIT('h82)
	) name14274 (
		_w3654_,
		_w11274_,
		_w11276_,
		_w14308_
	);
	LUT2 #(
		.INIT('h8)
	) name14275 (
		_w3311_,
		_w11394_,
		_w14309_
	);
	LUT4 #(
		.INIT('h2228)
	) name14276 (
		_w3645_,
		_w8466_,
		_w8541_,
		_w11273_,
		_w14310_
	);
	LUT2 #(
		.INIT('h1)
	) name14277 (
		_w14309_,
		_w14310_,
		_w14311_
	);
	LUT2 #(
		.INIT('h4)
	) name14278 (
		_w14308_,
		_w14311_,
		_w14312_
	);
	LUT4 #(
		.INIT('h4844)
	) name14279 (
		\a[20] ,
		_w14306_,
		_w14307_,
		_w14312_,
		_w14313_
	);
	LUT4 #(
		.INIT('h9699)
	) name14280 (
		\a[20] ,
		_w14306_,
		_w14307_,
		_w14312_,
		_w14314_
	);
	LUT3 #(
		.INIT('h1e)
	) name14281 (
		_w14194_,
		_w14196_,
		_w14314_,
		_w14315_
	);
	LUT4 #(
		.INIT('h6500)
	) name14282 (
		\a[17] ,
		_w14262_,
		_w14267_,
		_w14315_,
		_w14316_
	);
	LUT4 #(
		.INIT('h9a65)
	) name14283 (
		\a[17] ,
		_w14262_,
		_w14267_,
		_w14315_,
		_w14317_
	);
	LUT3 #(
		.INIT('h1e)
	) name14284 (
		_w14198_,
		_w14200_,
		_w14317_,
		_w14318_
	);
	LUT3 #(
		.INIT('h82)
	) name14285 (
		_w4034_,
		_w11490_,
		_w11492_,
		_w14319_
	);
	LUT3 #(
		.INIT('h82)
	) name14286 (
		_w4382_,
		_w11286_,
		_w11335_,
		_w14320_
	);
	LUT2 #(
		.INIT('h8)
	) name14287 (
		_w4033_,
		_w11382_,
		_w14321_
	);
	LUT4 #(
		.INIT('h2228)
	) name14288 (
		_w4367_,
		_w7695_,
		_w7750_,
		_w11285_,
		_w14322_
	);
	LUT2 #(
		.INIT('h1)
	) name14289 (
		_w14321_,
		_w14322_,
		_w14323_
	);
	LUT2 #(
		.INIT('h4)
	) name14290 (
		_w14320_,
		_w14323_,
		_w14324_
	);
	LUT4 #(
		.INIT('h4844)
	) name14291 (
		\a[14] ,
		_w14318_,
		_w14319_,
		_w14324_,
		_w14325_
	);
	LUT4 #(
		.INIT('h9699)
	) name14292 (
		\a[14] ,
		_w14318_,
		_w14319_,
		_w14324_,
		_w14326_
	);
	LUT3 #(
		.INIT('h1e)
	) name14293 (
		_w14207_,
		_w14209_,
		_w14326_,
		_w14327_
	);
	LUT4 #(
		.INIT('h6500)
	) name14294 (
		\a[11] ,
		_w14256_,
		_w14261_,
		_w14327_,
		_w14328_
	);
	LUT4 #(
		.INIT('h9a65)
	) name14295 (
		\a[11] ,
		_w14256_,
		_w14261_,
		_w14327_,
		_w14329_
	);
	LUT3 #(
		.INIT('h1e)
	) name14296 (
		_w14211_,
		_w14213_,
		_w14329_,
		_w14330_
	);
	LUT3 #(
		.INIT('h82)
	) name14297 (
		_w4876_,
		_w13292_,
		_w13325_,
		_w14331_
	);
	LUT3 #(
		.INIT('h82)
	) name14298 (
		_w5286_,
		_w13293_,
		_w13322_,
		_w14332_
	);
	LUT2 #(
		.INIT('h8)
	) name14299 (
		_w4875_,
		_w13247_,
		_w14333_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14300 (
		_w5271_,
		_w13243_,
		_w13245_,
		_w13285_,
		_w14334_
	);
	LUT2 #(
		.INIT('h1)
	) name14301 (
		_w14333_,
		_w14334_,
		_w14335_
	);
	LUT2 #(
		.INIT('h4)
	) name14302 (
		_w14332_,
		_w14335_,
		_w14336_
	);
	LUT4 #(
		.INIT('h4844)
	) name14303 (
		\a[8] ,
		_w14330_,
		_w14331_,
		_w14336_,
		_w14337_
	);
	LUT4 #(
		.INIT('h9699)
	) name14304 (
		\a[8] ,
		_w14330_,
		_w14331_,
		_w14336_,
		_w14338_
	);
	LUT3 #(
		.INIT('h1e)
	) name14305 (
		_w14220_,
		_w14222_,
		_w14338_,
		_w14339_
	);
	LUT4 #(
		.INIT('h6500)
	) name14306 (
		\a[5] ,
		_w14250_,
		_w14255_,
		_w14339_,
		_w14340_
	);
	LUT4 #(
		.INIT('h9a65)
	) name14307 (
		\a[5] ,
		_w14250_,
		_w14255_,
		_w14339_,
		_w14341_
	);
	LUT3 #(
		.INIT('h1e)
	) name14308 (
		_w14224_,
		_w14226_,
		_w14341_,
		_w14342_
	);
	LUT4 #(
		.INIT('h010f)
	) name14309 (
		_w14113_,
		_w14115_,
		_w14237_,
		_w14238_,
		_w14343_
	);
	LUT4 #(
		.INIT('h00f1)
	) name14310 (
		_w14108_,
		_w14111_,
		_w14233_,
		_w14234_,
		_w14344_
	);
	LUT3 #(
		.INIT('h01)
	) name14311 (
		\a[29] ,
		\a[30] ,
		\a[31] ,
		_w14345_
	);
	LUT3 #(
		.INIT('h0b)
	) name14312 (
		_w7136_,
		_w7166_,
		_w14345_,
		_w14346_
	);
	LUT3 #(
		.INIT('h87)
	) name14313 (
		_w373_,
		_w14230_,
		_w14346_,
		_w14347_
	);
	LUT3 #(
		.INIT('h28)
	) name14314 (
		_w14236_,
		_w14344_,
		_w14347_,
		_w14348_
	);
	LUT3 #(
		.INIT('h96)
	) name14315 (
		_w14236_,
		_w14344_,
		_w14347_,
		_w14349_
	);
	LUT3 #(
		.INIT('h82)
	) name14316 (
		_w6335_,
		_w14343_,
		_w14349_,
		_w14350_
	);
	LUT3 #(
		.INIT('h28)
	) name14317 (
		_w6657_,
		_w14344_,
		_w14347_,
		_w14351_
	);
	LUT2 #(
		.INIT('h8)
	) name14318 (
		_w6334_,
		_w14112_,
		_w14352_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14319 (
		_w6650_,
		_w14108_,
		_w14111_,
		_w14235_,
		_w14353_
	);
	LUT2 #(
		.INIT('h1)
	) name14320 (
		_w14352_,
		_w14353_,
		_w14354_
	);
	LUT2 #(
		.INIT('h4)
	) name14321 (
		_w14351_,
		_w14354_,
		_w14355_
	);
	LUT4 #(
		.INIT('h4844)
	) name14322 (
		\a[2] ,
		_w14342_,
		_w14350_,
		_w14355_,
		_w14356_
	);
	LUT4 #(
		.INIT('h9699)
	) name14323 (
		\a[2] ,
		_w14342_,
		_w14350_,
		_w14355_,
		_w14357_
	);
	LUT4 #(
		.INIT('h4d00)
	) name14324 (
		_w14126_,
		_w14227_,
		_w14244_,
		_w14357_,
		_w14358_
	);
	LUT4 #(
		.INIT('h32cd)
	) name14325 (
		_w14126_,
		_w14245_,
		_w14246_,
		_w14357_,
		_w14359_
	);
	LUT2 #(
		.INIT('h8)
	) name14326 (
		_w14248_,
		_w14359_,
		_w14360_
	);
	LUT2 #(
		.INIT('h6)
	) name14327 (
		_w14248_,
		_w14359_,
		_w14361_
	);
	LUT4 #(
		.INIT('h010f)
	) name14328 (
		_w14224_,
		_w14226_,
		_w14340_,
		_w14341_,
		_w14362_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name14329 (
		_w6335_,
		_w14343_,
		_w14348_,
		_w14349_,
		_w14363_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14330 (
		_w6334_,
		_w14108_,
		_w14111_,
		_w14235_,
		_w14364_
	);
	LUT4 #(
		.INIT('h00d7)
	) name14331 (
		_w10590_,
		_w14344_,
		_w14347_,
		_w14364_,
		_w14365_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14332 (
		_w5524_,
		_w13712_,
		_w13714_,
		_w13847_,
		_w14366_
	);
	LUT4 #(
		.INIT('h007d)
	) name14333 (
		_w6031_,
		_w13960_,
		_w13979_,
		_w14366_,
		_w14367_
	);
	LUT3 #(
		.INIT('h70)
	) name14334 (
		_w6324_,
		_w14112_,
		_w14367_,
		_w14368_
	);
	LUT4 #(
		.INIT('h95aa)
	) name14335 (
		\a[5] ,
		_w35_,
		_w14116_,
		_w14368_,
		_w14369_
	);
	LUT4 #(
		.INIT('h010f)
	) name14336 (
		_w14220_,
		_w14222_,
		_w14337_,
		_w14338_,
		_w14370_
	);
	LUT4 #(
		.INIT('h010f)
	) name14337 (
		_w14211_,
		_w14213_,
		_w14328_,
		_w14329_,
		_w14371_
	);
	LUT4 #(
		.INIT('h2228)
	) name14338 (
		_w4458_,
		_w11549_,
		_w11373_,
		_w11375_,
		_w14372_
	);
	LUT4 #(
		.INIT('h007d)
	) name14339 (
		_w4684_,
		_w13062_,
		_w13099_,
		_w14372_,
		_w14373_
	);
	LUT3 #(
		.INIT('h70)
	) name14340 (
		_w4700_,
		_w13247_,
		_w14373_,
		_w14374_
	);
	LUT4 #(
		.INIT('h95aa)
	) name14341 (
		\a[11] ,
		_w4459_,
		_w13576_,
		_w14374_,
		_w14375_
	);
	LUT4 #(
		.INIT('h010f)
	) name14342 (
		_w14207_,
		_w14209_,
		_w14325_,
		_w14326_,
		_w14376_
	);
	LUT4 #(
		.INIT('h010f)
	) name14343 (
		_w14198_,
		_w14200_,
		_w14316_,
		_w14317_,
		_w14377_
	);
	LUT4 #(
		.INIT('h2228)
	) name14344 (
		_w3709_,
		_w7935_,
		_w8077_,
		_w11279_,
		_w14378_
	);
	LUT4 #(
		.INIT('h007d)
	) name14345 (
		_w3877_,
		_w11280_,
		_w11282_,
		_w14378_,
		_w14379_
	);
	LUT3 #(
		.INIT('h70)
	) name14346 (
		_w3886_,
		_w11382_,
		_w14379_,
		_w14380_
	);
	LUT4 #(
		.INIT('h95aa)
	) name14347 (
		\a[17] ,
		_w3710_,
		_w12476_,
		_w14380_,
		_w14381_
	);
	LUT4 #(
		.INIT('h010f)
	) name14348 (
		_w14194_,
		_w14196_,
		_w14313_,
		_w14314_,
		_w14382_
	);
	LUT4 #(
		.INIT('h010f)
	) name14349 (
		_w14185_,
		_w14187_,
		_w14304_,
		_w14305_,
		_w14383_
	);
	LUT4 #(
		.INIT('h2228)
	) name14350 (
		_w3214_,
		_w8794_,
		_w8994_,
		_w11267_,
		_w14384_
	);
	LUT4 #(
		.INIT('h007d)
	) name14351 (
		_w3249_,
		_w11268_,
		_w11270_,
		_w14384_,
		_w14385_
	);
	LUT3 #(
		.INIT('h70)
	) name14352 (
		_w3262_,
		_w11394_,
		_w14385_,
		_w14386_
	);
	LUT4 #(
		.INIT('h95aa)
	) name14353 (
		\a[23] ,
		_w37_,
		_w12209_,
		_w14386_,
		_w14387_
	);
	LUT4 #(
		.INIT('h010f)
	) name14354 (
		_w14181_,
		_w14183_,
		_w14301_,
		_w14302_,
		_w14388_
	);
	LUT3 #(
		.INIT('h32)
	) name14355 (
		_w14274_,
		_w14291_,
		_w14292_,
		_w14389_
	);
	LUT3 #(
		.INIT('h82)
	) name14356 (
		_w2549_,
		_w10268_,
		_w11255_,
		_w14390_
	);
	LUT4 #(
		.INIT('h007d)
	) name14357 (
		_w2617_,
		_w11256_,
		_w11258_,
		_w14390_,
		_w14391_
	);
	LUT3 #(
		.INIT('h70)
	) name14358 (
		_w2854_,
		_w11406_,
		_w14391_,
		_w14392_
	);
	LUT4 #(
		.INIT('h95aa)
	) name14359 (
		\a[29] ,
		_w2550_,
		_w11796_,
		_w14392_,
		_w14393_
	);
	LUT4 #(
		.INIT('hf110)
	) name14360 (
		_w14168_,
		_w14170_,
		_w14285_,
		_w14289_,
		_w14394_
	);
	LUT3 #(
		.INIT('h80)
	) name14361 (
		_w978_,
		_w1012_,
		_w1433_,
		_w14395_
	);
	LUT3 #(
		.INIT('h80)
	) name14362 (
		_w7626_,
		_w14028_,
		_w14395_,
		_w14396_
	);
	LUT4 #(
		.INIT('h135f)
	) name14363 (
		_w122_,
		_w110_,
		_w46_,
		_w158_,
		_w14397_
	);
	LUT2 #(
		.INIT('h8)
	) name14364 (
		_w575_,
		_w14397_,
		_w14398_
	);
	LUT3 #(
		.INIT('h80)
	) name14365 (
		_w1603_,
		_w1673_,
		_w3442_,
		_w14399_
	);
	LUT2 #(
		.INIT('h8)
	) name14366 (
		_w14398_,
		_w14399_,
		_w14400_
	);
	LUT4 #(
		.INIT('h135f)
	) name14367 (
		_w55_,
		_w59_,
		_w72_,
		_w43_,
		_w14401_
	);
	LUT4 #(
		.INIT('h8000)
	) name14368 (
		_w663_,
		_w807_,
		_w962_,
		_w14401_,
		_w14402_
	);
	LUT4 #(
		.INIT('h153f)
	) name14369 (
		_w122_,
		_w67_,
		_w72_,
		_w65_,
		_w14403_
	);
	LUT4 #(
		.INIT('h135f)
	) name14370 (
		_w55_,
		_w50_,
		_w166_,
		_w259_,
		_w14404_
	);
	LUT4 #(
		.INIT('h8000)
	) name14371 (
		_w305_,
		_w609_,
		_w14403_,
		_w14404_,
		_w14405_
	);
	LUT4 #(
		.INIT('h8000)
	) name14372 (
		_w14398_,
		_w14399_,
		_w14402_,
		_w14405_,
		_w14406_
	);
	LUT2 #(
		.INIT('h8)
	) name14373 (
		_w14396_,
		_w14406_,
		_w14407_
	);
	LUT3 #(
		.INIT('h80)
	) name14374 (
		_w2085_,
		_w3454_,
		_w7850_,
		_w14408_
	);
	LUT2 #(
		.INIT('h8)
	) name14375 (
		_w14407_,
		_w14408_,
		_w14409_
	);
	LUT2 #(
		.INIT('h8)
	) name14376 (
		_w376_,
		_w11415_,
		_w14410_
	);
	LUT4 #(
		.INIT('h007d)
	) name14377 (
		_w2407_,
		_w10599_,
		_w11253_,
		_w14410_,
		_w14411_
	);
	LUT4 #(
		.INIT('h7d00)
	) name14378 (
		_w2527_,
		_w10580_,
		_w11254_,
		_w14411_,
		_w14412_
	);
	LUT4 #(
		.INIT('h7d00)
	) name14379 (
		_w377_,
		_w11453_,
		_w11455_,
		_w14412_,
		_w14413_
	);
	LUT3 #(
		.INIT('h69)
	) name14380 (
		_w14394_,
		_w14409_,
		_w14413_,
		_w14414_
	);
	LUT2 #(
		.INIT('h4)
	) name14381 (
		_w14393_,
		_w14414_,
		_w14415_
	);
	LUT2 #(
		.INIT('h2)
	) name14382 (
		_w14393_,
		_w14414_,
		_w14416_
	);
	LUT2 #(
		.INIT('h9)
	) name14383 (
		_w14393_,
		_w14414_,
		_w14417_
	);
	LUT2 #(
		.INIT('h9)
	) name14384 (
		_w14389_,
		_w14417_,
		_w14418_
	);
	LUT4 #(
		.INIT('h2228)
	) name14385 (
		_w2874_,
		_w9446_,
		_w9702_,
		_w11261_,
		_w14419_
	);
	LUT4 #(
		.INIT('h007d)
	) name14386 (
		_w2975_,
		_w11262_,
		_w11264_,
		_w14419_,
		_w14420_
	);
	LUT3 #(
		.INIT('h70)
	) name14387 (
		_w2986_,
		_w11400_,
		_w14420_,
		_w14421_
	);
	LUT4 #(
		.INIT('h95aa)
	) name14388 (
		\a[26] ,
		_w2875_,
		_w11967_,
		_w14421_,
		_w14422_
	);
	LUT2 #(
		.INIT('h2)
	) name14389 (
		_w14418_,
		_w14422_,
		_w14423_
	);
	LUT2 #(
		.INIT('h4)
	) name14390 (
		_w14418_,
		_w14422_,
		_w14424_
	);
	LUT2 #(
		.INIT('h9)
	) name14391 (
		_w14418_,
		_w14422_,
		_w14425_
	);
	LUT2 #(
		.INIT('h9)
	) name14392 (
		_w14388_,
		_w14425_,
		_w14426_
	);
	LUT2 #(
		.INIT('h4)
	) name14393 (
		_w14387_,
		_w14426_,
		_w14427_
	);
	LUT2 #(
		.INIT('h2)
	) name14394 (
		_w14387_,
		_w14426_,
		_w14428_
	);
	LUT2 #(
		.INIT('h9)
	) name14395 (
		_w14387_,
		_w14426_,
		_w14429_
	);
	LUT2 #(
		.INIT('h9)
	) name14396 (
		_w14383_,
		_w14429_,
		_w14430_
	);
	LUT4 #(
		.INIT('h2228)
	) name14397 (
		_w3311_,
		_w8466_,
		_w8541_,
		_w11273_,
		_w14431_
	);
	LUT4 #(
		.INIT('h007d)
	) name14398 (
		_w3645_,
		_w11274_,
		_w11276_,
		_w14431_,
		_w14432_
	);
	LUT3 #(
		.INIT('h70)
	) name14399 (
		_w3654_,
		_w11388_,
		_w14432_,
		_w14433_
	);
	LUT4 #(
		.INIT('h95aa)
	) name14400 (
		\a[20] ,
		_w3312_,
		_w12391_,
		_w14433_,
		_w14434_
	);
	LUT2 #(
		.INIT('h2)
	) name14401 (
		_w14430_,
		_w14434_,
		_w14435_
	);
	LUT2 #(
		.INIT('h4)
	) name14402 (
		_w14430_,
		_w14434_,
		_w14436_
	);
	LUT2 #(
		.INIT('h9)
	) name14403 (
		_w14430_,
		_w14434_,
		_w14437_
	);
	LUT2 #(
		.INIT('h9)
	) name14404 (
		_w14382_,
		_w14437_,
		_w14438_
	);
	LUT2 #(
		.INIT('h4)
	) name14405 (
		_w14381_,
		_w14438_,
		_w14439_
	);
	LUT2 #(
		.INIT('h2)
	) name14406 (
		_w14381_,
		_w14438_,
		_w14440_
	);
	LUT2 #(
		.INIT('h9)
	) name14407 (
		_w14381_,
		_w14438_,
		_w14441_
	);
	LUT2 #(
		.INIT('h9)
	) name14408 (
		_w14377_,
		_w14441_,
		_w14442_
	);
	LUT4 #(
		.INIT('h2228)
	) name14409 (
		_w4033_,
		_w7695_,
		_w7750_,
		_w11285_,
		_w14443_
	);
	LUT4 #(
		.INIT('h007d)
	) name14410 (
		_w4367_,
		_w11286_,
		_w11335_,
		_w14443_,
		_w14444_
	);
	LUT3 #(
		.INIT('h70)
	) name14411 (
		_w4382_,
		_w11377_,
		_w14444_,
		_w14445_
	);
	LUT4 #(
		.INIT('h95aa)
	) name14412 (
		\a[14] ,
		_w4034_,
		_w12799_,
		_w14445_,
		_w14446_
	);
	LUT2 #(
		.INIT('h2)
	) name14413 (
		_w14442_,
		_w14446_,
		_w14447_
	);
	LUT2 #(
		.INIT('h4)
	) name14414 (
		_w14442_,
		_w14446_,
		_w14448_
	);
	LUT2 #(
		.INIT('h9)
	) name14415 (
		_w14442_,
		_w14446_,
		_w14449_
	);
	LUT2 #(
		.INIT('h9)
	) name14416 (
		_w14376_,
		_w14449_,
		_w14450_
	);
	LUT2 #(
		.INIT('h4)
	) name14417 (
		_w14375_,
		_w14450_,
		_w14451_
	);
	LUT2 #(
		.INIT('h2)
	) name14418 (
		_w14375_,
		_w14450_,
		_w14452_
	);
	LUT2 #(
		.INIT('h9)
	) name14419 (
		_w14375_,
		_w14450_,
		_w14453_
	);
	LUT2 #(
		.INIT('h9)
	) name14420 (
		_w14371_,
		_w14453_,
		_w14454_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14421 (
		_w4875_,
		_w13243_,
		_w13245_,
		_w13285_,
		_w14455_
	);
	LUT4 #(
		.INIT('h007d)
	) name14422 (
		_w5271_,
		_w13293_,
		_w13322_,
		_w14455_,
		_w14456_
	);
	LUT3 #(
		.INIT('h70)
	) name14423 (
		_w5286_,
		_w13716_,
		_w14456_,
		_w14457_
	);
	LUT4 #(
		.INIT('h95aa)
	) name14424 (
		\a[8] ,
		_w4876_,
		_w13720_,
		_w14457_,
		_w14458_
	);
	LUT2 #(
		.INIT('h2)
	) name14425 (
		_w14454_,
		_w14458_,
		_w14459_
	);
	LUT2 #(
		.INIT('h4)
	) name14426 (
		_w14454_,
		_w14458_,
		_w14460_
	);
	LUT2 #(
		.INIT('h9)
	) name14427 (
		_w14454_,
		_w14458_,
		_w14461_
	);
	LUT2 #(
		.INIT('h9)
	) name14428 (
		_w14370_,
		_w14461_,
		_w14462_
	);
	LUT2 #(
		.INIT('h4)
	) name14429 (
		_w14369_,
		_w14462_,
		_w14463_
	);
	LUT2 #(
		.INIT('h9)
	) name14430 (
		_w14369_,
		_w14462_,
		_w14464_
	);
	LUT4 #(
		.INIT('h6500)
	) name14431 (
		\a[2] ,
		_w14363_,
		_w14365_,
		_w14464_,
		_w14465_
	);
	LUT4 #(
		.INIT('h9a65)
	) name14432 (
		\a[2] ,
		_w14363_,
		_w14365_,
		_w14464_,
		_w14466_
	);
	LUT2 #(
		.INIT('h2)
	) name14433 (
		_w14362_,
		_w14466_,
		_w14467_
	);
	LUT2 #(
		.INIT('h4)
	) name14434 (
		_w14362_,
		_w14466_,
		_w14468_
	);
	LUT2 #(
		.INIT('h9)
	) name14435 (
		_w14362_,
		_w14466_,
		_w14469_
	);
	LUT3 #(
		.INIT('h1e)
	) name14436 (
		_w14356_,
		_w14358_,
		_w14469_,
		_w14470_
	);
	LUT2 #(
		.INIT('h8)
	) name14437 (
		_w14360_,
		_w14470_,
		_w14471_
	);
	LUT2 #(
		.INIT('h6)
	) name14438 (
		_w14360_,
		_w14470_,
		_w14472_
	);
	LUT2 #(
		.INIT('h1)
	) name14439 (
		_w14463_,
		_w14465_,
		_w14473_
	);
	LUT3 #(
		.INIT('h32)
	) name14440 (
		_w14370_,
		_w14459_,
		_w14460_,
		_w14474_
	);
	LUT3 #(
		.INIT('h32)
	) name14441 (
		_w14371_,
		_w14451_,
		_w14452_,
		_w14475_
	);
	LUT3 #(
		.INIT('h32)
	) name14442 (
		_w14376_,
		_w14447_,
		_w14448_,
		_w14476_
	);
	LUT3 #(
		.INIT('h32)
	) name14443 (
		_w14377_,
		_w14439_,
		_w14440_,
		_w14477_
	);
	LUT3 #(
		.INIT('h32)
	) name14444 (
		_w14382_,
		_w14435_,
		_w14436_,
		_w14478_
	);
	LUT3 #(
		.INIT('h32)
	) name14445 (
		_w14383_,
		_w14427_,
		_w14428_,
		_w14479_
	);
	LUT3 #(
		.INIT('h32)
	) name14446 (
		_w14388_,
		_w14423_,
		_w14424_,
		_w14480_
	);
	LUT3 #(
		.INIT('h32)
	) name14447 (
		_w14389_,
		_w14415_,
		_w14416_,
		_w14481_
	);
	LUT3 #(
		.INIT('he8)
	) name14448 (
		_w14394_,
		_w14409_,
		_w14413_,
		_w14482_
	);
	LUT4 #(
		.INIT('h0777)
	) name14449 (
		_w122_,
		_w110_,
		_w78_,
		_w56_,
		_w14483_
	);
	LUT4 #(
		.INIT('h0777)
	) name14450 (
		_w38_,
		_w43_,
		_w65_,
		_w236_,
		_w14484_
	);
	LUT4 #(
		.INIT('h8000)
	) name14451 (
		_w1359_,
		_w1915_,
		_w14483_,
		_w14484_,
		_w14485_
	);
	LUT4 #(
		.INIT('h8000)
	) name14452 (
		_w793_,
		_w902_,
		_w2234_,
		_w7230_,
		_w14486_
	);
	LUT4 #(
		.INIT('h8000)
	) name14453 (
		_w491_,
		_w737_,
		_w2072_,
		_w2136_,
		_w14487_
	);
	LUT4 #(
		.INIT('h8000)
	) name14454 (
		_w4272_,
		_w14487_,
		_w14485_,
		_w14486_,
		_w14488_
	);
	LUT4 #(
		.INIT('h8000)
	) name14455 (
		_w163_,
		_w173_,
		_w1782_,
		_w1786_,
		_w14489_
	);
	LUT4 #(
		.INIT('h8000)
	) name14456 (
		_w2132_,
		_w7205_,
		_w14488_,
		_w14489_,
		_w14490_
	);
	LUT2 #(
		.INIT('h8)
	) name14457 (
		_w587_,
		_w14490_,
		_w14491_
	);
	LUT4 #(
		.INIT('h5ee5)
	) name14458 (
		\a[2] ,
		_w7844_,
		_w14344_,
		_w14347_,
		_w14492_
	);
	LUT3 #(
		.INIT('h82)
	) name14459 (
		_w376_,
		_w10599_,
		_w11253_,
		_w14493_
	);
	LUT4 #(
		.INIT('h007d)
	) name14460 (
		_w2407_,
		_w10580_,
		_w11254_,
		_w14493_,
		_w14494_
	);
	LUT4 #(
		.INIT('h7d00)
	) name14461 (
		_w2527_,
		_w10268_,
		_w11255_,
		_w14494_,
		_w14495_
	);
	LUT4 #(
		.INIT('h7d00)
	) name14462 (
		_w377_,
		_w11456_,
		_w11458_,
		_w14495_,
		_w14496_
	);
	LUT4 #(
		.INIT('h8228)
	) name14463 (
		_w14482_,
		_w14491_,
		_w14492_,
		_w14496_,
		_w14497_
	);
	LUT4 #(
		.INIT('h1441)
	) name14464 (
		_w14482_,
		_w14491_,
		_w14492_,
		_w14496_,
		_w14498_
	);
	LUT4 #(
		.INIT('h6996)
	) name14465 (
		_w14482_,
		_w14491_,
		_w14492_,
		_w14496_,
		_w14499_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14466 (
		_w2550_,
		_w11408_,
		_w11463_,
		_w11464_,
		_w14500_
	);
	LUT4 #(
		.INIT('h2228)
	) name14467 (
		_w2854_,
		_w9446_,
		_w9702_,
		_w11261_,
		_w14501_
	);
	LUT3 #(
		.INIT('h82)
	) name14468 (
		_w2549_,
		_w11256_,
		_w11258_,
		_w14502_
	);
	LUT3 #(
		.INIT('h07)
	) name14469 (
		_w2617_,
		_w11406_,
		_w14502_,
		_w14503_
	);
	LUT2 #(
		.INIT('h4)
	) name14470 (
		_w14501_,
		_w14503_,
		_w14504_
	);
	LUT3 #(
		.INIT('h9a)
	) name14471 (
		\a[29] ,
		_w14500_,
		_w14504_,
		_w14505_
	);
	LUT3 #(
		.INIT('h82)
	) name14472 (
		_w2875_,
		_w11469_,
		_w11471_,
		_w14506_
	);
	LUT4 #(
		.INIT('h2228)
	) name14473 (
		_w2986_,
		_w8794_,
		_w8994_,
		_w11267_,
		_w14507_
	);
	LUT3 #(
		.INIT('h82)
	) name14474 (
		_w2874_,
		_w11262_,
		_w11264_,
		_w14508_
	);
	LUT3 #(
		.INIT('h07)
	) name14475 (
		_w2975_,
		_w11400_,
		_w14508_,
		_w14509_
	);
	LUT2 #(
		.INIT('h4)
	) name14476 (
		_w14507_,
		_w14509_,
		_w14510_
	);
	LUT3 #(
		.INIT('h9a)
	) name14477 (
		\a[26] ,
		_w14506_,
		_w14510_,
		_w14511_
	);
	LUT4 #(
		.INIT('h9669)
	) name14478 (
		_w14481_,
		_w14499_,
		_w14505_,
		_w14511_,
		_w14512_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14479 (
		_w37_,
		_w11396_,
		_w11476_,
		_w11477_,
		_w14513_
	);
	LUT4 #(
		.INIT('h2228)
	) name14480 (
		_w3262_,
		_w8466_,
		_w8541_,
		_w11273_,
		_w14514_
	);
	LUT3 #(
		.INIT('h82)
	) name14481 (
		_w3214_,
		_w11268_,
		_w11270_,
		_w14515_
	);
	LUT3 #(
		.INIT('h07)
	) name14482 (
		_w3249_,
		_w11394_,
		_w14515_,
		_w14516_
	);
	LUT2 #(
		.INIT('h4)
	) name14483 (
		_w14514_,
		_w14516_,
		_w14517_
	);
	LUT3 #(
		.INIT('h9a)
	) name14484 (
		\a[23] ,
		_w14513_,
		_w14517_,
		_w14518_
	);
	LUT4 #(
		.INIT('h2882)
	) name14485 (
		_w14479_,
		_w14480_,
		_w14512_,
		_w14518_,
		_w14519_
	);
	LUT4 #(
		.INIT('h4114)
	) name14486 (
		_w14479_,
		_w14480_,
		_w14512_,
		_w14518_,
		_w14520_
	);
	LUT4 #(
		.INIT('h9669)
	) name14487 (
		_w14479_,
		_w14480_,
		_w14512_,
		_w14518_,
		_w14521_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14488 (
		_w3312_,
		_w11390_,
		_w11482_,
		_w11483_,
		_w14522_
	);
	LUT4 #(
		.INIT('h2228)
	) name14489 (
		_w3654_,
		_w7935_,
		_w8077_,
		_w11279_,
		_w14523_
	);
	LUT3 #(
		.INIT('h82)
	) name14490 (
		_w3311_,
		_w11274_,
		_w11276_,
		_w14524_
	);
	LUT3 #(
		.INIT('h07)
	) name14491 (
		_w3645_,
		_w11388_,
		_w14524_,
		_w14525_
	);
	LUT2 #(
		.INIT('h4)
	) name14492 (
		_w14523_,
		_w14525_,
		_w14526_
	);
	LUT3 #(
		.INIT('h9a)
	) name14493 (
		\a[20] ,
		_w14522_,
		_w14526_,
		_w14527_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14494 (
		_w3710_,
		_w11384_,
		_w11488_,
		_w11489_,
		_w14528_
	);
	LUT4 #(
		.INIT('h2228)
	) name14495 (
		_w3886_,
		_w7695_,
		_w7750_,
		_w11285_,
		_w14529_
	);
	LUT3 #(
		.INIT('h82)
	) name14496 (
		_w3709_,
		_w11280_,
		_w11282_,
		_w14530_
	);
	LUT3 #(
		.INIT('h07)
	) name14497 (
		_w3877_,
		_w11382_,
		_w14530_,
		_w14531_
	);
	LUT2 #(
		.INIT('h4)
	) name14498 (
		_w14529_,
		_w14531_,
		_w14532_
	);
	LUT3 #(
		.INIT('h9a)
	) name14499 (
		\a[17] ,
		_w14528_,
		_w14532_,
		_w14533_
	);
	LUT4 #(
		.INIT('h9669)
	) name14500 (
		_w14478_,
		_w14521_,
		_w14527_,
		_w14533_,
		_w14534_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14501 (
		_w4034_,
		_w11378_,
		_w11494_,
		_w11552_,
		_w14535_
	);
	LUT4 #(
		.INIT('h2228)
	) name14502 (
		_w4382_,
		_w11549_,
		_w11373_,
		_w11375_,
		_w14536_
	);
	LUT3 #(
		.INIT('h82)
	) name14503 (
		_w4033_,
		_w11286_,
		_w11335_,
		_w14537_
	);
	LUT3 #(
		.INIT('h07)
	) name14504 (
		_w4367_,
		_w11377_,
		_w14537_,
		_w14538_
	);
	LUT2 #(
		.INIT('h4)
	) name14505 (
		_w14536_,
		_w14538_,
		_w14539_
	);
	LUT3 #(
		.INIT('h9a)
	) name14506 (
		\a[14] ,
		_w14535_,
		_w14539_,
		_w14540_
	);
	LUT4 #(
		.INIT('h2882)
	) name14507 (
		_w14476_,
		_w14477_,
		_w14534_,
		_w14540_,
		_w14541_
	);
	LUT4 #(
		.INIT('h4114)
	) name14508 (
		_w14476_,
		_w14477_,
		_w14534_,
		_w14540_,
		_w14542_
	);
	LUT4 #(
		.INIT('h9669)
	) name14509 (
		_w14476_,
		_w14477_,
		_w14534_,
		_w14540_,
		_w14543_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14510 (
		_w4459_,
		_w13288_,
		_w13290_,
		_w13291_,
		_w14544_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14511 (
		_w4700_,
		_w13243_,
		_w13245_,
		_w13285_,
		_w14545_
	);
	LUT3 #(
		.INIT('h82)
	) name14512 (
		_w4458_,
		_w13062_,
		_w13099_,
		_w14546_
	);
	LUT3 #(
		.INIT('h07)
	) name14513 (
		_w4684_,
		_w13247_,
		_w14546_,
		_w14547_
	);
	LUT2 #(
		.INIT('h4)
	) name14514 (
		_w14545_,
		_w14547_,
		_w14548_
	);
	LUT3 #(
		.INIT('h9a)
	) name14515 (
		\a[11] ,
		_w14544_,
		_w14548_,
		_w14549_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14516 (
		_w4876_,
		_w13717_,
		_w13719_,
		_w13850_,
		_w14550_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14517 (
		_w5286_,
		_w13712_,
		_w13714_,
		_w13847_,
		_w14551_
	);
	LUT3 #(
		.INIT('h82)
	) name14518 (
		_w4875_,
		_w13293_,
		_w13322_,
		_w14552_
	);
	LUT3 #(
		.INIT('h07)
	) name14519 (
		_w5271_,
		_w13716_,
		_w14552_,
		_w14553_
	);
	LUT2 #(
		.INIT('h4)
	) name14520 (
		_w14551_,
		_w14553_,
		_w14554_
	);
	LUT3 #(
		.INIT('h9a)
	) name14521 (
		\a[8] ,
		_w14550_,
		_w14554_,
		_w14555_
	);
	LUT4 #(
		.INIT('h9669)
	) name14522 (
		_w14475_,
		_w14543_,
		_w14549_,
		_w14555_,
		_w14556_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14523 (
		_w35_,
		_w14113_,
		_w14115_,
		_w14238_,
		_w14557_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14524 (
		_w6324_,
		_w14108_,
		_w14111_,
		_w14235_,
		_w14558_
	);
	LUT3 #(
		.INIT('h82)
	) name14525 (
		_w5524_,
		_w13960_,
		_w13979_,
		_w14559_
	);
	LUT3 #(
		.INIT('h07)
	) name14526 (
		_w6031_,
		_w14112_,
		_w14559_,
		_w14560_
	);
	LUT2 #(
		.INIT('h4)
	) name14527 (
		_w14558_,
		_w14560_,
		_w14561_
	);
	LUT3 #(
		.INIT('h9a)
	) name14528 (
		\a[5] ,
		_w14557_,
		_w14561_,
		_w14562_
	);
	LUT4 #(
		.INIT('h2882)
	) name14529 (
		_w14473_,
		_w14474_,
		_w14556_,
		_w14562_,
		_w14563_
	);
	LUT4 #(
		.INIT('h4114)
	) name14530 (
		_w14473_,
		_w14474_,
		_w14556_,
		_w14562_,
		_w14564_
	);
	LUT4 #(
		.INIT('h9669)
	) name14531 (
		_w14473_,
		_w14474_,
		_w14556_,
		_w14562_,
		_w14565_
	);
	LUT4 #(
		.INIT('h00f1)
	) name14532 (
		_w14356_,
		_w14358_,
		_w14467_,
		_w14468_,
		_w14566_
	);
	LUT3 #(
		.INIT('h82)
	) name14533 (
		_w14471_,
		_w14565_,
		_w14566_,
		_w14567_
	);
	LUT3 #(
		.INIT('h69)
	) name14534 (
		_w14471_,
		_w14565_,
		_w14566_,
		_w14568_
	);
	LUT3 #(
		.INIT('h82)
	) name14535 (
		_w2875_,
		_w11472_,
		_w11474_,
		_w14569_
	);
	LUT3 #(
		.INIT('h82)
	) name14536 (
		_w2986_,
		_w11268_,
		_w11270_,
		_w14570_
	);
	LUT2 #(
		.INIT('h8)
	) name14537 (
		_w2874_,
		_w11400_,
		_w14571_
	);
	LUT4 #(
		.INIT('h2228)
	) name14538 (
		_w2975_,
		_w8794_,
		_w8994_,
		_w11267_,
		_w14572_
	);
	LUT2 #(
		.INIT('h1)
	) name14539 (
		_w14571_,
		_w14572_,
		_w14573_
	);
	LUT2 #(
		.INIT('h4)
	) name14540 (
		_w14570_,
		_w14573_,
		_w14574_
	);
	LUT3 #(
		.INIT('h9a)
	) name14541 (
		\a[26] ,
		_w14569_,
		_w14574_,
		_w14575_
	);
	LUT3 #(
		.INIT('h32)
	) name14542 (
		_w14497_,
		_w14498_,
		_w14505_,
		_w14576_
	);
	LUT4 #(
		.INIT('h153f)
	) name14543 (
		_w122_,
		_w106_,
		_w55_,
		_w47_,
		_w14577_
	);
	LUT4 #(
		.INIT('h8000)
	) name14544 (
		_w225_,
		_w292_,
		_w384_,
		_w14577_,
		_w14578_
	);
	LUT4 #(
		.INIT('h8000)
	) name14545 (
		_w1480_,
		_w1754_,
		_w2060_,
		_w2706_,
		_w14579_
	);
	LUT4 #(
		.INIT('h8000)
	) name14546 (
		_w966_,
		_w1037_,
		_w1221_,
		_w1350_,
		_w14580_
	);
	LUT4 #(
		.INIT('h8000)
	) name14547 (
		_w12419_,
		_w14579_,
		_w14580_,
		_w14578_,
		_w14581_
	);
	LUT4 #(
		.INIT('h153f)
	) name14548 (
		_w52_,
		_w65_,
		_w166_,
		_w430_,
		_w14582_
	);
	LUT3 #(
		.INIT('h40)
	) name14549 (
		_w77_,
		_w81_,
		_w14582_,
		_w14583_
	);
	LUT4 #(
		.INIT('h8000)
	) name14550 (
		_w1443_,
		_w1446_,
		_w8368_,
		_w14583_,
		_w14584_
	);
	LUT4 #(
		.INIT('h8000)
	) name14551 (
		_w1903_,
		_w1914_,
		_w14581_,
		_w14584_,
		_w14585_
	);
	LUT2 #(
		.INIT('h8)
	) name14552 (
		_w8350_,
		_w14585_,
		_w14586_
	);
	LUT4 #(
		.INIT('h24db)
	) name14553 (
		_w14491_,
		_w14492_,
		_w14496_,
		_w14586_,
		_w14587_
	);
	LUT3 #(
		.INIT('h82)
	) name14554 (
		_w376_,
		_w10580_,
		_w11254_,
		_w14588_
	);
	LUT4 #(
		.INIT('h007d)
	) name14555 (
		_w2407_,
		_w10268_,
		_w11255_,
		_w14588_,
		_w14589_
	);
	LUT4 #(
		.INIT('h7d00)
	) name14556 (
		_w2527_,
		_w11256_,
		_w11258_,
		_w14589_,
		_w14590_
	);
	LUT4 #(
		.INIT('h7d00)
	) name14557 (
		_w377_,
		_w11459_,
		_w11461_,
		_w14590_,
		_w14591_
	);
	LUT2 #(
		.INIT('h2)
	) name14558 (
		_w14587_,
		_w14591_,
		_w14592_
	);
	LUT2 #(
		.INIT('h4)
	) name14559 (
		_w14587_,
		_w14591_,
		_w14593_
	);
	LUT2 #(
		.INIT('h9)
	) name14560 (
		_w14587_,
		_w14591_,
		_w14594_
	);
	LUT3 #(
		.INIT('h82)
	) name14561 (
		_w2550_,
		_w11465_,
		_w11467_,
		_w14595_
	);
	LUT3 #(
		.INIT('h82)
	) name14562 (
		_w2854_,
		_w11262_,
		_w11264_,
		_w14596_
	);
	LUT2 #(
		.INIT('h8)
	) name14563 (
		_w2549_,
		_w11406_,
		_w14597_
	);
	LUT4 #(
		.INIT('h2228)
	) name14564 (
		_w2617_,
		_w9446_,
		_w9702_,
		_w11261_,
		_w14598_
	);
	LUT2 #(
		.INIT('h1)
	) name14565 (
		_w14597_,
		_w14598_,
		_w14599_
	);
	LUT2 #(
		.INIT('h4)
	) name14566 (
		_w14596_,
		_w14599_,
		_w14600_
	);
	LUT3 #(
		.INIT('h9a)
	) name14567 (
		\a[29] ,
		_w14595_,
		_w14600_,
		_w14601_
	);
	LUT4 #(
		.INIT('h9669)
	) name14568 (
		_w14575_,
		_w14576_,
		_w14594_,
		_w14601_,
		_w14602_
	);
	LUT4 #(
		.INIT('h41d7)
	) name14569 (
		_w14481_,
		_w14499_,
		_w14505_,
		_w14511_,
		_w14603_
	);
	LUT3 #(
		.INIT('h82)
	) name14570 (
		_w37_,
		_w11478_,
		_w11480_,
		_w14604_
	);
	LUT3 #(
		.INIT('h82)
	) name14571 (
		_w3262_,
		_w11274_,
		_w11276_,
		_w14605_
	);
	LUT2 #(
		.INIT('h8)
	) name14572 (
		_w3214_,
		_w11394_,
		_w14606_
	);
	LUT4 #(
		.INIT('h2228)
	) name14573 (
		_w3249_,
		_w8466_,
		_w8541_,
		_w11273_,
		_w14607_
	);
	LUT2 #(
		.INIT('h1)
	) name14574 (
		_w14606_,
		_w14607_,
		_w14608_
	);
	LUT2 #(
		.INIT('h4)
	) name14575 (
		_w14605_,
		_w14608_,
		_w14609_
	);
	LUT3 #(
		.INIT('h9a)
	) name14576 (
		\a[23] ,
		_w14604_,
		_w14609_,
		_w14610_
	);
	LUT3 #(
		.INIT('h4d)
	) name14577 (
		_w14480_,
		_w14512_,
		_w14518_,
		_w14611_
	);
	LUT4 #(
		.INIT('h0096)
	) name14578 (
		_w14602_,
		_w14603_,
		_w14610_,
		_w14611_,
		_w14612_
	);
	LUT4 #(
		.INIT('h6900)
	) name14579 (
		_w14602_,
		_w14603_,
		_w14610_,
		_w14611_,
		_w14613_
	);
	LUT4 #(
		.INIT('h9669)
	) name14580 (
		_w14602_,
		_w14603_,
		_w14610_,
		_w14611_,
		_w14614_
	);
	LUT3 #(
		.INIT('h82)
	) name14581 (
		_w3312_,
		_w11484_,
		_w11486_,
		_w14615_
	);
	LUT3 #(
		.INIT('h82)
	) name14582 (
		_w3654_,
		_w11280_,
		_w11282_,
		_w14616_
	);
	LUT2 #(
		.INIT('h8)
	) name14583 (
		_w3311_,
		_w11388_,
		_w14617_
	);
	LUT4 #(
		.INIT('h2228)
	) name14584 (
		_w3645_,
		_w7935_,
		_w8077_,
		_w11279_,
		_w14618_
	);
	LUT2 #(
		.INIT('h1)
	) name14585 (
		_w14617_,
		_w14618_,
		_w14619_
	);
	LUT2 #(
		.INIT('h4)
	) name14586 (
		_w14616_,
		_w14619_,
		_w14620_
	);
	LUT3 #(
		.INIT('h9a)
	) name14587 (
		\a[20] ,
		_w14615_,
		_w14620_,
		_w14621_
	);
	LUT3 #(
		.INIT('h45)
	) name14588 (
		_w14519_,
		_w14520_,
		_w14527_,
		_w14622_
	);
	LUT3 #(
		.INIT('h82)
	) name14589 (
		_w3710_,
		_w11490_,
		_w11492_,
		_w14623_
	);
	LUT3 #(
		.INIT('h82)
	) name14590 (
		_w3886_,
		_w11286_,
		_w11335_,
		_w14624_
	);
	LUT2 #(
		.INIT('h8)
	) name14591 (
		_w3709_,
		_w11382_,
		_w14625_
	);
	LUT4 #(
		.INIT('h2228)
	) name14592 (
		_w3877_,
		_w7695_,
		_w7750_,
		_w11285_,
		_w14626_
	);
	LUT2 #(
		.INIT('h1)
	) name14593 (
		_w14625_,
		_w14626_,
		_w14627_
	);
	LUT2 #(
		.INIT('h4)
	) name14594 (
		_w14624_,
		_w14627_,
		_w14628_
	);
	LUT3 #(
		.INIT('h9a)
	) name14595 (
		\a[17] ,
		_w14623_,
		_w14628_,
		_w14629_
	);
	LUT4 #(
		.INIT('h6996)
	) name14596 (
		_w14614_,
		_w14621_,
		_w14622_,
		_w14629_,
		_w14630_
	);
	LUT4 #(
		.INIT('h41d7)
	) name14597 (
		_w14478_,
		_w14521_,
		_w14527_,
		_w14533_,
		_w14631_
	);
	LUT3 #(
		.INIT('h82)
	) name14598 (
		_w4034_,
		_w13061_,
		_w13102_,
		_w14632_
	);
	LUT3 #(
		.INIT('h82)
	) name14599 (
		_w4382_,
		_w13062_,
		_w13099_,
		_w14633_
	);
	LUT2 #(
		.INIT('h8)
	) name14600 (
		_w4033_,
		_w11377_,
		_w14634_
	);
	LUT4 #(
		.INIT('h2228)
	) name14601 (
		_w4367_,
		_w11549_,
		_w11373_,
		_w11375_,
		_w14635_
	);
	LUT2 #(
		.INIT('h1)
	) name14602 (
		_w14634_,
		_w14635_,
		_w14636_
	);
	LUT2 #(
		.INIT('h4)
	) name14603 (
		_w14633_,
		_w14636_,
		_w14637_
	);
	LUT3 #(
		.INIT('h9a)
	) name14604 (
		\a[14] ,
		_w14632_,
		_w14637_,
		_w14638_
	);
	LUT3 #(
		.INIT('h4d)
	) name14605 (
		_w14477_,
		_w14534_,
		_w14540_,
		_w14639_
	);
	LUT4 #(
		.INIT('h0096)
	) name14606 (
		_w14630_,
		_w14631_,
		_w14638_,
		_w14639_,
		_w14640_
	);
	LUT4 #(
		.INIT('h6900)
	) name14607 (
		_w14630_,
		_w14631_,
		_w14638_,
		_w14639_,
		_w14641_
	);
	LUT4 #(
		.INIT('h9669)
	) name14608 (
		_w14630_,
		_w14631_,
		_w14638_,
		_w14639_,
		_w14642_
	);
	LUT3 #(
		.INIT('h82)
	) name14609 (
		_w4459_,
		_w13292_,
		_w13325_,
		_w14643_
	);
	LUT3 #(
		.INIT('h82)
	) name14610 (
		_w4700_,
		_w13293_,
		_w13322_,
		_w14644_
	);
	LUT2 #(
		.INIT('h8)
	) name14611 (
		_w4458_,
		_w13247_,
		_w14645_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14612 (
		_w4684_,
		_w13243_,
		_w13245_,
		_w13285_,
		_w14646_
	);
	LUT2 #(
		.INIT('h1)
	) name14613 (
		_w14645_,
		_w14646_,
		_w14647_
	);
	LUT2 #(
		.INIT('h4)
	) name14614 (
		_w14644_,
		_w14647_,
		_w14648_
	);
	LUT3 #(
		.INIT('h9a)
	) name14615 (
		\a[11] ,
		_w14643_,
		_w14648_,
		_w14649_
	);
	LUT3 #(
		.INIT('h45)
	) name14616 (
		_w14541_,
		_w14542_,
		_w14549_,
		_w14650_
	);
	LUT3 #(
		.INIT('h82)
	) name14617 (
		_w4876_,
		_w13959_,
		_w13982_,
		_w14651_
	);
	LUT3 #(
		.INIT('h82)
	) name14618 (
		_w5286_,
		_w13960_,
		_w13979_,
		_w14652_
	);
	LUT2 #(
		.INIT('h8)
	) name14619 (
		_w4875_,
		_w13716_,
		_w14653_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14620 (
		_w5271_,
		_w13712_,
		_w13714_,
		_w13847_,
		_w14654_
	);
	LUT2 #(
		.INIT('h1)
	) name14621 (
		_w14653_,
		_w14654_,
		_w14655_
	);
	LUT2 #(
		.INIT('h4)
	) name14622 (
		_w14652_,
		_w14655_,
		_w14656_
	);
	LUT3 #(
		.INIT('h9a)
	) name14623 (
		\a[8] ,
		_w14651_,
		_w14656_,
		_w14657_
	);
	LUT4 #(
		.INIT('h6996)
	) name14624 (
		_w14642_,
		_w14649_,
		_w14650_,
		_w14657_,
		_w14658_
	);
	LUT4 #(
		.INIT('h41d7)
	) name14625 (
		_w14475_,
		_w14543_,
		_w14549_,
		_w14555_,
		_w14659_
	);
	LUT3 #(
		.INIT('h82)
	) name14626 (
		_w35_,
		_w14343_,
		_w14349_,
		_w14660_
	);
	LUT3 #(
		.INIT('h28)
	) name14627 (
		_w6324_,
		_w14344_,
		_w14347_,
		_w14661_
	);
	LUT2 #(
		.INIT('h8)
	) name14628 (
		_w5524_,
		_w14112_,
		_w14662_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14629 (
		_w6031_,
		_w14108_,
		_w14111_,
		_w14235_,
		_w14663_
	);
	LUT2 #(
		.INIT('h1)
	) name14630 (
		_w14662_,
		_w14663_,
		_w14664_
	);
	LUT2 #(
		.INIT('h4)
	) name14631 (
		_w14661_,
		_w14664_,
		_w14665_
	);
	LUT3 #(
		.INIT('h9a)
	) name14632 (
		\a[5] ,
		_w14660_,
		_w14665_,
		_w14666_
	);
	LUT3 #(
		.INIT('h4d)
	) name14633 (
		_w14474_,
		_w14556_,
		_w14562_,
		_w14667_
	);
	LUT4 #(
		.INIT('h0096)
	) name14634 (
		_w14658_,
		_w14659_,
		_w14666_,
		_w14667_,
		_w14668_
	);
	LUT4 #(
		.INIT('h6900)
	) name14635 (
		_w14658_,
		_w14659_,
		_w14666_,
		_w14667_,
		_w14669_
	);
	LUT4 #(
		.INIT('h9669)
	) name14636 (
		_w14658_,
		_w14659_,
		_w14666_,
		_w14667_,
		_w14670_
	);
	LUT3 #(
		.INIT('h32)
	) name14637 (
		_w14563_,
		_w14564_,
		_w14566_,
		_w14671_
	);
	LUT3 #(
		.INIT('h82)
	) name14638 (
		_w14567_,
		_w14670_,
		_w14671_,
		_w14672_
	);
	LUT3 #(
		.INIT('h69)
	) name14639 (
		_w14567_,
		_w14670_,
		_w14671_,
		_w14673_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name14640 (
		_w35_,
		_w14343_,
		_w14348_,
		_w14349_,
		_w14674_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14641 (
		_w5524_,
		_w14108_,
		_w14111_,
		_w14235_,
		_w14675_
	);
	LUT4 #(
		.INIT('h00eb)
	) name14642 (
		_w7866_,
		_w14344_,
		_w14347_,
		_w14675_,
		_w14676_
	);
	LUT3 #(
		.INIT('h9a)
	) name14643 (
		\a[5] ,
		_w14674_,
		_w14676_,
		_w14677_
	);
	LUT4 #(
		.INIT('h90f9)
	) name14644 (
		_w14642_,
		_w14649_,
		_w14650_,
		_w14657_,
		_w14678_
	);
	LUT2 #(
		.INIT('h4)
	) name14645 (
		_w14677_,
		_w14678_,
		_w14679_
	);
	LUT2 #(
		.INIT('h2)
	) name14646 (
		_w14677_,
		_w14678_,
		_w14680_
	);
	LUT2 #(
		.INIT('h9)
	) name14647 (
		_w14677_,
		_w14678_,
		_w14681_
	);
	LUT4 #(
		.INIT('hbe28)
	) name14648 (
		_w14575_,
		_w14576_,
		_w14594_,
		_w14601_,
		_w14682_
	);
	LUT4 #(
		.INIT('h2228)
	) name14649 (
		_w2874_,
		_w8794_,
		_w8994_,
		_w11267_,
		_w14683_
	);
	LUT4 #(
		.INIT('h007d)
	) name14650 (
		_w2975_,
		_w11268_,
		_w11270_,
		_w14683_,
		_w14684_
	);
	LUT3 #(
		.INIT('h70)
	) name14651 (
		_w2986_,
		_w11394_,
		_w14684_,
		_w14685_
	);
	LUT4 #(
		.INIT('h95aa)
	) name14652 (
		\a[26] ,
		_w2875_,
		_w12209_,
		_w14685_,
		_w14686_
	);
	LUT4 #(
		.INIT('hecc8)
	) name14653 (
		_w14491_,
		_w14492_,
		_w14496_,
		_w14586_,
		_w14687_
	);
	LUT4 #(
		.INIT('h8000)
	) name14654 (
		_w649_,
		_w1297_,
		_w2073_,
		_w2281_,
		_w14688_
	);
	LUT3 #(
		.INIT('h80)
	) name14655 (
		_w2656_,
		_w7973_,
		_w14688_,
		_w14689_
	);
	LUT4 #(
		.INIT('h153f)
	) name14656 (
		_w56_,
		_w93_,
		_w419_,
		_w378_,
		_w14690_
	);
	LUT4 #(
		.INIT('h153f)
	) name14657 (
		_w67_,
		_w39_,
		_w93_,
		_w236_,
		_w14691_
	);
	LUT4 #(
		.INIT('h4000)
	) name14658 (
		_w431_,
		_w611_,
		_w14691_,
		_w14690_,
		_w14692_
	);
	LUT4 #(
		.INIT('h8000)
	) name14659 (
		_w1038_,
		_w1042_,
		_w2087_,
		_w14692_,
		_w14693_
	);
	LUT3 #(
		.INIT('h80)
	) name14660 (
		_w3541_,
		_w14689_,
		_w14693_,
		_w14694_
	);
	LUT3 #(
		.INIT('h80)
	) name14661 (
		_w1136_,
		_w1939_,
		_w14694_,
		_w14695_
	);
	LUT2 #(
		.INIT('h1)
	) name14662 (
		_w14492_,
		_w14695_,
		_w14696_
	);
	LUT2 #(
		.INIT('h8)
	) name14663 (
		_w14492_,
		_w14695_,
		_w14697_
	);
	LUT2 #(
		.INIT('h6)
	) name14664 (
		_w14492_,
		_w14695_,
		_w14698_
	);
	LUT3 #(
		.INIT('h82)
	) name14665 (
		_w376_,
		_w10268_,
		_w11255_,
		_w14699_
	);
	LUT4 #(
		.INIT('h007d)
	) name14666 (
		_w2407_,
		_w11256_,
		_w11258_,
		_w14699_,
		_w14700_
	);
	LUT3 #(
		.INIT('h70)
	) name14667 (
		_w2527_,
		_w11406_,
		_w14700_,
		_w14701_
	);
	LUT3 #(
		.INIT('h70)
	) name14668 (
		_w377_,
		_w11796_,
		_w14701_,
		_w14702_
	);
	LUT3 #(
		.INIT('h09)
	) name14669 (
		_w14687_,
		_w14698_,
		_w14702_,
		_w14703_
	);
	LUT3 #(
		.INIT('h96)
	) name14670 (
		_w14687_,
		_w14698_,
		_w14702_,
		_w14704_
	);
	LUT4 #(
		.INIT('h4d00)
	) name14671 (
		_w14576_,
		_w14587_,
		_w14591_,
		_w14704_,
		_w14705_
	);
	LUT4 #(
		.INIT('h32cd)
	) name14672 (
		_w14576_,
		_w14592_,
		_w14593_,
		_w14704_,
		_w14706_
	);
	LUT4 #(
		.INIT('h2228)
	) name14673 (
		_w2549_,
		_w9446_,
		_w9702_,
		_w11261_,
		_w14707_
	);
	LUT4 #(
		.INIT('h007d)
	) name14674 (
		_w2617_,
		_w11262_,
		_w11264_,
		_w14707_,
		_w14708_
	);
	LUT3 #(
		.INIT('h70)
	) name14675 (
		_w2854_,
		_w11400_,
		_w14708_,
		_w14709_
	);
	LUT4 #(
		.INIT('h95aa)
	) name14676 (
		\a[29] ,
		_w2550_,
		_w11967_,
		_w14709_,
		_w14710_
	);
	LUT4 #(
		.INIT('h2882)
	) name14677 (
		_w14682_,
		_w14686_,
		_w14706_,
		_w14710_,
		_w14711_
	);
	LUT4 #(
		.INIT('h4114)
	) name14678 (
		_w14682_,
		_w14686_,
		_w14706_,
		_w14710_,
		_w14712_
	);
	LUT4 #(
		.INIT('h9669)
	) name14679 (
		_w14682_,
		_w14686_,
		_w14706_,
		_w14710_,
		_w14713_
	);
	LUT4 #(
		.INIT('h2228)
	) name14680 (
		_w3214_,
		_w8466_,
		_w8541_,
		_w11273_,
		_w14714_
	);
	LUT4 #(
		.INIT('h007d)
	) name14681 (
		_w3249_,
		_w11274_,
		_w11276_,
		_w14714_,
		_w14715_
	);
	LUT3 #(
		.INIT('h70)
	) name14682 (
		_w3262_,
		_w11388_,
		_w14715_,
		_w14716_
	);
	LUT4 #(
		.INIT('h95aa)
	) name14683 (
		\a[23] ,
		_w37_,
		_w12391_,
		_w14716_,
		_w14717_
	);
	LUT3 #(
		.INIT('h8e)
	) name14684 (
		_w14602_,
		_w14603_,
		_w14610_,
		_w14718_
	);
	LUT4 #(
		.INIT('h2228)
	) name14685 (
		_w3311_,
		_w7935_,
		_w8077_,
		_w11279_,
		_w14719_
	);
	LUT4 #(
		.INIT('h007d)
	) name14686 (
		_w3645_,
		_w11280_,
		_w11282_,
		_w14719_,
		_w14720_
	);
	LUT3 #(
		.INIT('h70)
	) name14687 (
		_w3654_,
		_w11382_,
		_w14720_,
		_w14721_
	);
	LUT4 #(
		.INIT('h95aa)
	) name14688 (
		\a[20] ,
		_w3312_,
		_w12476_,
		_w14721_,
		_w14722_
	);
	LUT4 #(
		.INIT('h6996)
	) name14689 (
		_w14713_,
		_w14717_,
		_w14718_,
		_w14722_,
		_w14723_
	);
	LUT3 #(
		.INIT('h45)
	) name14690 (
		_w14612_,
		_w14613_,
		_w14621_,
		_w14724_
	);
	LUT4 #(
		.INIT('h2228)
	) name14691 (
		_w3709_,
		_w7695_,
		_w7750_,
		_w11285_,
		_w14725_
	);
	LUT4 #(
		.INIT('h007d)
	) name14692 (
		_w3877_,
		_w11286_,
		_w11335_,
		_w14725_,
		_w14726_
	);
	LUT3 #(
		.INIT('h70)
	) name14693 (
		_w3886_,
		_w11377_,
		_w14726_,
		_w14727_
	);
	LUT4 #(
		.INIT('h95aa)
	) name14694 (
		\a[17] ,
		_w3710_,
		_w12799_,
		_w14727_,
		_w14728_
	);
	LUT3 #(
		.INIT('h69)
	) name14695 (
		_w14723_,
		_w14724_,
		_w14728_,
		_w14729_
	);
	LUT4 #(
		.INIT('h90f9)
	) name14696 (
		_w14614_,
		_w14621_,
		_w14622_,
		_w14629_,
		_w14730_
	);
	LUT4 #(
		.INIT('h0096)
	) name14697 (
		_w14723_,
		_w14724_,
		_w14728_,
		_w14730_,
		_w14731_
	);
	LUT4 #(
		.INIT('h6900)
	) name14698 (
		_w14723_,
		_w14724_,
		_w14728_,
		_w14730_,
		_w14732_
	);
	LUT4 #(
		.INIT('h9669)
	) name14699 (
		_w14723_,
		_w14724_,
		_w14728_,
		_w14730_,
		_w14733_
	);
	LUT4 #(
		.INIT('h2228)
	) name14700 (
		_w4033_,
		_w11549_,
		_w11373_,
		_w11375_,
		_w14734_
	);
	LUT4 #(
		.INIT('h007d)
	) name14701 (
		_w4367_,
		_w13062_,
		_w13099_,
		_w14734_,
		_w14735_
	);
	LUT3 #(
		.INIT('h70)
	) name14702 (
		_w4382_,
		_w13247_,
		_w14735_,
		_w14736_
	);
	LUT4 #(
		.INIT('h95aa)
	) name14703 (
		\a[14] ,
		_w4034_,
		_w13576_,
		_w14736_,
		_w14737_
	);
	LUT3 #(
		.INIT('h8e)
	) name14704 (
		_w14630_,
		_w14631_,
		_w14638_,
		_w14738_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14705 (
		_w4458_,
		_w13243_,
		_w13245_,
		_w13285_,
		_w14739_
	);
	LUT4 #(
		.INIT('h007d)
	) name14706 (
		_w4684_,
		_w13293_,
		_w13322_,
		_w14739_,
		_w14740_
	);
	LUT3 #(
		.INIT('h70)
	) name14707 (
		_w4700_,
		_w13716_,
		_w14740_,
		_w14741_
	);
	LUT4 #(
		.INIT('h95aa)
	) name14708 (
		\a[11] ,
		_w4459_,
		_w13720_,
		_w14741_,
		_w14742_
	);
	LUT4 #(
		.INIT('h6996)
	) name14709 (
		_w14733_,
		_w14737_,
		_w14738_,
		_w14742_,
		_w14743_
	);
	LUT3 #(
		.INIT('h45)
	) name14710 (
		_w14640_,
		_w14641_,
		_w14649_,
		_w14744_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14711 (
		_w4875_,
		_w13712_,
		_w13714_,
		_w13847_,
		_w14745_
	);
	LUT4 #(
		.INIT('h007d)
	) name14712 (
		_w5271_,
		_w13960_,
		_w13979_,
		_w14745_,
		_w14746_
	);
	LUT3 #(
		.INIT('h70)
	) name14713 (
		_w5286_,
		_w14112_,
		_w14746_,
		_w14747_
	);
	LUT4 #(
		.INIT('h95aa)
	) name14714 (
		\a[8] ,
		_w4876_,
		_w14116_,
		_w14747_,
		_w14748_
	);
	LUT3 #(
		.INIT('h69)
	) name14715 (
		_w14743_,
		_w14744_,
		_w14748_,
		_w14749_
	);
	LUT3 #(
		.INIT('h8e)
	) name14716 (
		_w14658_,
		_w14659_,
		_w14666_,
		_w14750_
	);
	LUT3 #(
		.INIT('h09)
	) name14717 (
		_w14681_,
		_w14749_,
		_w14750_,
		_w14751_
	);
	LUT3 #(
		.INIT('h60)
	) name14718 (
		_w14681_,
		_w14749_,
		_w14750_,
		_w14752_
	);
	LUT3 #(
		.INIT('h96)
	) name14719 (
		_w14681_,
		_w14749_,
		_w14750_,
		_w14753_
	);
	LUT3 #(
		.INIT('h32)
	) name14720 (
		_w14668_,
		_w14669_,
		_w14671_,
		_w14754_
	);
	LUT3 #(
		.INIT('h82)
	) name14721 (
		_w14672_,
		_w14753_,
		_w14754_,
		_w14755_
	);
	LUT3 #(
		.INIT('h69)
	) name14722 (
		_w14672_,
		_w14753_,
		_w14754_,
		_w14756_
	);
	LUT3 #(
		.INIT('h32)
	) name14723 (
		_w14751_,
		_w14752_,
		_w14754_,
		_w14757_
	);
	LUT3 #(
		.INIT('hb2)
	) name14724 (
		_w14686_,
		_w14706_,
		_w14710_,
		_w14758_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14725 (
		_w2875_,
		_w11396_,
		_w11476_,
		_w11477_,
		_w14759_
	);
	LUT4 #(
		.INIT('h2228)
	) name14726 (
		_w2986_,
		_w8466_,
		_w8541_,
		_w11273_,
		_w14760_
	);
	LUT3 #(
		.INIT('h82)
	) name14727 (
		_w2874_,
		_w11268_,
		_w11270_,
		_w14761_
	);
	LUT3 #(
		.INIT('h07)
	) name14728 (
		_w2975_,
		_w11394_,
		_w14761_,
		_w14762_
	);
	LUT2 #(
		.INIT('h4)
	) name14729 (
		_w14760_,
		_w14762_,
		_w14763_
	);
	LUT3 #(
		.INIT('h9a)
	) name14730 (
		\a[26] ,
		_w14759_,
		_w14763_,
		_w14764_
	);
	LUT3 #(
		.INIT('h32)
	) name14731 (
		_w14687_,
		_w14696_,
		_w14697_,
		_w14765_
	);
	LUT4 #(
		.INIT('h5665)
	) name14732 (
		\a[5] ,
		_w7867_,
		_w14344_,
		_w14347_,
		_w14766_
	);
	LUT3 #(
		.INIT('h1f)
	) name14733 (
		_w90_,
		_w56_,
		_w72_,
		_w14767_
	);
	LUT3 #(
		.INIT('h57)
	) name14734 (
		_w38_,
		_w419_,
		_w430_,
		_w14768_
	);
	LUT4 #(
		.INIT('h8000)
	) name14735 (
		_w48_,
		_w150_,
		_w14767_,
		_w14768_,
		_w14769_
	);
	LUT4 #(
		.INIT('h8000)
	) name14736 (
		_w1275_,
		_w1341_,
		_w2125_,
		_w3134_,
		_w14770_
	);
	LUT4 #(
		.INIT('h8000)
	) name14737 (
		_w3450_,
		_w7338_,
		_w14770_,
		_w14769_,
		_w14771_
	);
	LUT4 #(
		.INIT('h8000)
	) name14738 (
		_w2743_,
		_w2751_,
		_w12148_,
		_w14771_,
		_w14772_
	);
	LUT2 #(
		.INIT('h8)
	) name14739 (
		_w1742_,
		_w14772_,
		_w14773_
	);
	LUT3 #(
		.INIT('h69)
	) name14740 (
		_w14492_,
		_w14766_,
		_w14773_,
		_w14774_
	);
	LUT4 #(
		.INIT('h1700)
	) name14741 (
		_w14492_,
		_w14687_,
		_w14695_,
		_w14774_,
		_w14775_
	);
	LUT4 #(
		.INIT('h00e8)
	) name14742 (
		_w14492_,
		_w14687_,
		_w14695_,
		_w14774_,
		_w14776_
	);
	LUT4 #(
		.INIT('h32cd)
	) name14743 (
		_w14687_,
		_w14696_,
		_w14697_,
		_w14774_,
		_w14777_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14744 (
		_w377_,
		_w11408_,
		_w11463_,
		_w11464_,
		_w14778_
	);
	LUT4 #(
		.INIT('h2228)
	) name14745 (
		_w2527_,
		_w9446_,
		_w9702_,
		_w11261_,
		_w14779_
	);
	LUT3 #(
		.INIT('h82)
	) name14746 (
		_w376_,
		_w11256_,
		_w11258_,
		_w14780_
	);
	LUT3 #(
		.INIT('h07)
	) name14747 (
		_w2407_,
		_w11406_,
		_w14780_,
		_w14781_
	);
	LUT2 #(
		.INIT('h4)
	) name14748 (
		_w14779_,
		_w14781_,
		_w14782_
	);
	LUT2 #(
		.INIT('h4)
	) name14749 (
		_w14778_,
		_w14782_,
		_w14783_
	);
	LUT2 #(
		.INIT('h9)
	) name14750 (
		_w14777_,
		_w14783_,
		_w14784_
	);
	LUT3 #(
		.INIT('h82)
	) name14751 (
		_w2550_,
		_w11469_,
		_w11471_,
		_w14785_
	);
	LUT4 #(
		.INIT('h2228)
	) name14752 (
		_w2854_,
		_w8794_,
		_w8994_,
		_w11267_,
		_w14786_
	);
	LUT3 #(
		.INIT('h82)
	) name14753 (
		_w2549_,
		_w11262_,
		_w11264_,
		_w14787_
	);
	LUT3 #(
		.INIT('h07)
	) name14754 (
		_w2617_,
		_w11400_,
		_w14787_,
		_w14788_
	);
	LUT2 #(
		.INIT('h4)
	) name14755 (
		_w14786_,
		_w14788_,
		_w14789_
	);
	LUT3 #(
		.INIT('h9a)
	) name14756 (
		\a[29] ,
		_w14785_,
		_w14789_,
		_w14790_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name14757 (
		_w14703_,
		_w14705_,
		_w14784_,
		_w14790_,
		_w14791_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14758 (
		_w37_,
		_w11390_,
		_w11482_,
		_w11483_,
		_w14792_
	);
	LUT4 #(
		.INIT('h2228)
	) name14759 (
		_w3262_,
		_w7935_,
		_w8077_,
		_w11279_,
		_w14793_
	);
	LUT3 #(
		.INIT('h82)
	) name14760 (
		_w3214_,
		_w11274_,
		_w11276_,
		_w14794_
	);
	LUT3 #(
		.INIT('h07)
	) name14761 (
		_w3249_,
		_w11388_,
		_w14794_,
		_w14795_
	);
	LUT2 #(
		.INIT('h4)
	) name14762 (
		_w14793_,
		_w14795_,
		_w14796_
	);
	LUT3 #(
		.INIT('h9a)
	) name14763 (
		\a[23] ,
		_w14792_,
		_w14796_,
		_w14797_
	);
	LUT4 #(
		.INIT('h0096)
	) name14764 (
		_w14758_,
		_w14764_,
		_w14791_,
		_w14797_,
		_w14798_
	);
	LUT4 #(
		.INIT('h6900)
	) name14765 (
		_w14758_,
		_w14764_,
		_w14791_,
		_w14797_,
		_w14799_
	);
	LUT4 #(
		.INIT('h9669)
	) name14766 (
		_w14758_,
		_w14764_,
		_w14791_,
		_w14797_,
		_w14800_
	);
	LUT3 #(
		.INIT('h45)
	) name14767 (
		_w14711_,
		_w14712_,
		_w14717_,
		_w14801_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14768 (
		_w3312_,
		_w11384_,
		_w11488_,
		_w11489_,
		_w14802_
	);
	LUT4 #(
		.INIT('h2228)
	) name14769 (
		_w3654_,
		_w7695_,
		_w7750_,
		_w11285_,
		_w14803_
	);
	LUT3 #(
		.INIT('h82)
	) name14770 (
		_w3311_,
		_w11280_,
		_w11282_,
		_w14804_
	);
	LUT3 #(
		.INIT('h07)
	) name14771 (
		_w3645_,
		_w11382_,
		_w14804_,
		_w14805_
	);
	LUT2 #(
		.INIT('h4)
	) name14772 (
		_w14803_,
		_w14805_,
		_w14806_
	);
	LUT3 #(
		.INIT('h9a)
	) name14773 (
		\a[20] ,
		_w14802_,
		_w14806_,
		_w14807_
	);
	LUT4 #(
		.INIT('h90f9)
	) name14774 (
		_w14713_,
		_w14717_,
		_w14718_,
		_w14722_,
		_w14808_
	);
	LUT4 #(
		.INIT('h9669)
	) name14775 (
		_w14800_,
		_w14801_,
		_w14807_,
		_w14808_,
		_w14809_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14776 (
		_w3710_,
		_w11378_,
		_w11494_,
		_w11552_,
		_w14810_
	);
	LUT4 #(
		.INIT('h2228)
	) name14777 (
		_w3886_,
		_w11549_,
		_w11373_,
		_w11375_,
		_w14811_
	);
	LUT3 #(
		.INIT('h82)
	) name14778 (
		_w3709_,
		_w11286_,
		_w11335_,
		_w14812_
	);
	LUT3 #(
		.INIT('h07)
	) name14779 (
		_w3877_,
		_w11377_,
		_w14812_,
		_w14813_
	);
	LUT2 #(
		.INIT('h4)
	) name14780 (
		_w14811_,
		_w14813_,
		_w14814_
	);
	LUT3 #(
		.INIT('h9a)
	) name14781 (
		\a[17] ,
		_w14810_,
		_w14814_,
		_w14815_
	);
	LUT3 #(
		.INIT('h8e)
	) name14782 (
		_w14723_,
		_w14724_,
		_w14728_,
		_w14816_
	);
	LUT3 #(
		.INIT('h69)
	) name14783 (
		_w14809_,
		_w14815_,
		_w14816_,
		_w14817_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14784 (
		_w4034_,
		_w13288_,
		_w13290_,
		_w13291_,
		_w14818_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14785 (
		_w4382_,
		_w13243_,
		_w13245_,
		_w13285_,
		_w14819_
	);
	LUT3 #(
		.INIT('h82)
	) name14786 (
		_w4033_,
		_w13062_,
		_w13099_,
		_w14820_
	);
	LUT3 #(
		.INIT('h07)
	) name14787 (
		_w4367_,
		_w13247_,
		_w14820_,
		_w14821_
	);
	LUT2 #(
		.INIT('h4)
	) name14788 (
		_w14819_,
		_w14821_,
		_w14822_
	);
	LUT3 #(
		.INIT('h9a)
	) name14789 (
		\a[14] ,
		_w14818_,
		_w14822_,
		_w14823_
	);
	LUT4 #(
		.INIT('h008e)
	) name14790 (
		_w14729_,
		_w14730_,
		_w14737_,
		_w14823_,
		_w14824_
	);
	LUT4 #(
		.INIT('h7100)
	) name14791 (
		_w14729_,
		_w14730_,
		_w14737_,
		_w14823_,
		_w14825_
	);
	LUT4 #(
		.INIT('h45ba)
	) name14792 (
		_w14731_,
		_w14732_,
		_w14737_,
		_w14823_,
		_w14826_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14793 (
		_w4459_,
		_w13717_,
		_w13719_,
		_w13850_,
		_w14827_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14794 (
		_w4700_,
		_w13712_,
		_w13714_,
		_w13847_,
		_w14828_
	);
	LUT3 #(
		.INIT('h82)
	) name14795 (
		_w4458_,
		_w13293_,
		_w13322_,
		_w14829_
	);
	LUT3 #(
		.INIT('h07)
	) name14796 (
		_w4684_,
		_w13716_,
		_w14829_,
		_w14830_
	);
	LUT2 #(
		.INIT('h4)
	) name14797 (
		_w14828_,
		_w14830_,
		_w14831_
	);
	LUT3 #(
		.INIT('h9a)
	) name14798 (
		\a[11] ,
		_w14827_,
		_w14831_,
		_w14832_
	);
	LUT4 #(
		.INIT('h90f9)
	) name14799 (
		_w14733_,
		_w14737_,
		_w14738_,
		_w14742_,
		_w14833_
	);
	LUT4 #(
		.INIT('h9669)
	) name14800 (
		_w14817_,
		_w14826_,
		_w14832_,
		_w14833_,
		_w14834_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14801 (
		_w4876_,
		_w14113_,
		_w14115_,
		_w14238_,
		_w14835_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14802 (
		_w5286_,
		_w14108_,
		_w14111_,
		_w14235_,
		_w14836_
	);
	LUT3 #(
		.INIT('h82)
	) name14803 (
		_w4875_,
		_w13960_,
		_w13979_,
		_w14837_
	);
	LUT3 #(
		.INIT('h07)
	) name14804 (
		_w5271_,
		_w14112_,
		_w14837_,
		_w14838_
	);
	LUT2 #(
		.INIT('h4)
	) name14805 (
		_w14836_,
		_w14838_,
		_w14839_
	);
	LUT3 #(
		.INIT('h9a)
	) name14806 (
		\a[8] ,
		_w14835_,
		_w14839_,
		_w14840_
	);
	LUT4 #(
		.INIT('h008e)
	) name14807 (
		_w14743_,
		_w14744_,
		_w14748_,
		_w14840_,
		_w14841_
	);
	LUT4 #(
		.INIT('h7100)
	) name14808 (
		_w14743_,
		_w14744_,
		_w14748_,
		_w14840_,
		_w14842_
	);
	LUT4 #(
		.INIT('h8e71)
	) name14809 (
		_w14743_,
		_w14744_,
		_w14748_,
		_w14840_,
		_w14843_
	);
	LUT2 #(
		.INIT('h6)
	) name14810 (
		_w14834_,
		_w14843_,
		_w14844_
	);
	LUT3 #(
		.INIT('h32)
	) name14811 (
		_w14679_,
		_w14680_,
		_w14749_,
		_w14845_
	);
	LUT2 #(
		.INIT('h8)
	) name14812 (
		_w14844_,
		_w14845_,
		_w14846_
	);
	LUT2 #(
		.INIT('h1)
	) name14813 (
		_w14844_,
		_w14845_,
		_w14847_
	);
	LUT2 #(
		.INIT('h6)
	) name14814 (
		_w14844_,
		_w14845_,
		_w14848_
	);
	LUT3 #(
		.INIT('h82)
	) name14815 (
		_w14755_,
		_w14757_,
		_w14848_,
		_w14849_
	);
	LUT3 #(
		.INIT('h69)
	) name14816 (
		_w14755_,
		_w14757_,
		_w14848_,
		_w14850_
	);
	LUT3 #(
		.INIT('h31)
	) name14817 (
		_w14834_,
		_w14841_,
		_w14842_,
		_w14851_
	);
	LUT4 #(
		.INIT('h90f9)
	) name14818 (
		_w14817_,
		_w14826_,
		_w14832_,
		_w14833_,
		_w14852_
	);
	LUT3 #(
		.INIT('h82)
	) name14819 (
		_w4459_,
		_w13959_,
		_w13982_,
		_w14853_
	);
	LUT3 #(
		.INIT('h82)
	) name14820 (
		_w4700_,
		_w13960_,
		_w13979_,
		_w14854_
	);
	LUT2 #(
		.INIT('h8)
	) name14821 (
		_w4458_,
		_w13716_,
		_w14855_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14822 (
		_w4684_,
		_w13712_,
		_w13714_,
		_w13847_,
		_w14856_
	);
	LUT2 #(
		.INIT('h1)
	) name14823 (
		_w14855_,
		_w14856_,
		_w14857_
	);
	LUT2 #(
		.INIT('h4)
	) name14824 (
		_w14854_,
		_w14857_,
		_w14858_
	);
	LUT3 #(
		.INIT('h9a)
	) name14825 (
		\a[11] ,
		_w14853_,
		_w14858_,
		_w14859_
	);
	LUT3 #(
		.INIT('h31)
	) name14826 (
		_w14817_,
		_w14824_,
		_w14825_,
		_w14860_
	);
	LUT3 #(
		.INIT('h4d)
	) name14827 (
		_w14809_,
		_w14815_,
		_w14816_,
		_w14861_
	);
	LUT4 #(
		.INIT('h90f9)
	) name14828 (
		_w14800_,
		_w14801_,
		_w14807_,
		_w14808_,
		_w14862_
	);
	LUT3 #(
		.INIT('h45)
	) name14829 (
		_w14798_,
		_w14799_,
		_w14801_,
		_w14863_
	);
	LUT3 #(
		.INIT('h8e)
	) name14830 (
		_w14758_,
		_w14764_,
		_w14791_,
		_w14864_
	);
	LUT3 #(
		.INIT('h54)
	) name14831 (
		_w14775_,
		_w14776_,
		_w14783_,
		_w14865_
	);
	LUT3 #(
		.INIT('h71)
	) name14832 (
		_w14492_,
		_w14766_,
		_w14773_,
		_w14866_
	);
	LUT3 #(
		.INIT('h80)
	) name14833 (
		_w1221_,
		_w1435_,
		_w1475_,
		_w14867_
	);
	LUT3 #(
		.INIT('h80)
	) name14834 (
		_w3935_,
		_w4271_,
		_w14867_,
		_w14868_
	);
	LUT4 #(
		.INIT('h153f)
	) name14835 (
		_w59_,
		_w46_,
		_w184_,
		_w236_,
		_w14869_
	);
	LUT4 #(
		.INIT('h8000)
	) name14836 (
		_w584_,
		_w652_,
		_w1067_,
		_w14869_,
		_w14870_
	);
	LUT4 #(
		.INIT('h8000)
	) name14837 (
		_w815_,
		_w819_,
		_w1394_,
		_w14870_,
		_w14871_
	);
	LUT2 #(
		.INIT('h8)
	) name14838 (
		_w14868_,
		_w14871_,
		_w14872_
	);
	LUT4 #(
		.INIT('h8000)
	) name14839 (
		_w1575_,
		_w1700_,
		_w2741_,
		_w2809_,
		_w14873_
	);
	LUT3 #(
		.INIT('h80)
	) name14840 (
		_w1090_,
		_w4252_,
		_w14873_,
		_w14874_
	);
	LUT4 #(
		.INIT('h0777)
	) name14841 (
		_w106_,
		_w67_,
		_w78_,
		_w93_,
		_w14875_
	);
	LUT4 #(
		.INIT('h8000)
	) name14842 (
		_w863_,
		_w861_,
		_w909_,
		_w14875_,
		_w14876_
	);
	LUT3 #(
		.INIT('h1f)
	) name14843 (
		_w67_,
		_w90_,
		_w236_,
		_w14877_
	);
	LUT4 #(
		.INIT('h4000)
	) name14844 (
		_w264_,
		_w895_,
		_w2288_,
		_w14877_,
		_w14878_
	);
	LUT4 #(
		.INIT('h8000)
	) name14845 (
		_w1539_,
		_w1543_,
		_w14876_,
		_w14878_,
		_w14879_
	);
	LUT4 #(
		.INIT('h8000)
	) name14846 (
		_w14868_,
		_w14871_,
		_w14874_,
		_w14879_,
		_w14880_
	);
	LUT2 #(
		.INIT('h8)
	) name14847 (
		_w1009_,
		_w14880_,
		_w14881_
	);
	LUT4 #(
		.INIT('h718e)
	) name14848 (
		_w14492_,
		_w14766_,
		_w14773_,
		_w14881_,
		_w14882_
	);
	LUT3 #(
		.INIT('h82)
	) name14849 (
		_w377_,
		_w11465_,
		_w11467_,
		_w14883_
	);
	LUT3 #(
		.INIT('h82)
	) name14850 (
		_w2527_,
		_w11262_,
		_w11264_,
		_w14884_
	);
	LUT2 #(
		.INIT('h8)
	) name14851 (
		_w376_,
		_w11406_,
		_w14885_
	);
	LUT4 #(
		.INIT('h2228)
	) name14852 (
		_w2407_,
		_w9446_,
		_w9702_,
		_w11261_,
		_w14886_
	);
	LUT2 #(
		.INIT('h1)
	) name14853 (
		_w14885_,
		_w14886_,
		_w14887_
	);
	LUT2 #(
		.INIT('h4)
	) name14854 (
		_w14884_,
		_w14887_,
		_w14888_
	);
	LUT2 #(
		.INIT('h4)
	) name14855 (
		_w14883_,
		_w14888_,
		_w14889_
	);
	LUT2 #(
		.INIT('h9)
	) name14856 (
		_w14882_,
		_w14889_,
		_w14890_
	);
	LUT4 #(
		.INIT('h00b2)
	) name14857 (
		_w14765_,
		_w14774_,
		_w14783_,
		_w14890_,
		_w14891_
	);
	LUT4 #(
		.INIT('h4d00)
	) name14858 (
		_w14765_,
		_w14774_,
		_w14783_,
		_w14890_,
		_w14892_
	);
	LUT4 #(
		.INIT('h54ab)
	) name14859 (
		_w14775_,
		_w14776_,
		_w14783_,
		_w14890_,
		_w14893_
	);
	LUT3 #(
		.INIT('h82)
	) name14860 (
		_w2550_,
		_w11472_,
		_w11474_,
		_w14894_
	);
	LUT3 #(
		.INIT('h82)
	) name14861 (
		_w2854_,
		_w11268_,
		_w11270_,
		_w14895_
	);
	LUT2 #(
		.INIT('h8)
	) name14862 (
		_w2549_,
		_w11400_,
		_w14896_
	);
	LUT4 #(
		.INIT('h2228)
	) name14863 (
		_w2617_,
		_w8794_,
		_w8994_,
		_w11267_,
		_w14897_
	);
	LUT2 #(
		.INIT('h1)
	) name14864 (
		_w14896_,
		_w14897_,
		_w14898_
	);
	LUT2 #(
		.INIT('h4)
	) name14865 (
		_w14895_,
		_w14898_,
		_w14899_
	);
	LUT3 #(
		.INIT('h9a)
	) name14866 (
		\a[29] ,
		_w14894_,
		_w14899_,
		_w14900_
	);
	LUT2 #(
		.INIT('h9)
	) name14867 (
		_w14893_,
		_w14900_,
		_w14901_
	);
	LUT4 #(
		.INIT('he0fe)
	) name14868 (
		_w14703_,
		_w14705_,
		_w14784_,
		_w14790_,
		_w14902_
	);
	LUT3 #(
		.INIT('h82)
	) name14869 (
		_w2875_,
		_w11478_,
		_w11480_,
		_w14903_
	);
	LUT3 #(
		.INIT('h82)
	) name14870 (
		_w2986_,
		_w11274_,
		_w11276_,
		_w14904_
	);
	LUT2 #(
		.INIT('h8)
	) name14871 (
		_w2874_,
		_w11394_,
		_w14905_
	);
	LUT4 #(
		.INIT('h2228)
	) name14872 (
		_w2975_,
		_w8466_,
		_w8541_,
		_w11273_,
		_w14906_
	);
	LUT2 #(
		.INIT('h1)
	) name14873 (
		_w14905_,
		_w14906_,
		_w14907_
	);
	LUT2 #(
		.INIT('h4)
	) name14874 (
		_w14904_,
		_w14907_,
		_w14908_
	);
	LUT3 #(
		.INIT('h9a)
	) name14875 (
		\a[26] ,
		_w14903_,
		_w14908_,
		_w14909_
	);
	LUT3 #(
		.INIT('h69)
	) name14876 (
		_w14901_,
		_w14902_,
		_w14909_,
		_w14910_
	);
	LUT3 #(
		.INIT('h82)
	) name14877 (
		_w37_,
		_w11484_,
		_w11486_,
		_w14911_
	);
	LUT3 #(
		.INIT('h82)
	) name14878 (
		_w3262_,
		_w11280_,
		_w11282_,
		_w14912_
	);
	LUT2 #(
		.INIT('h8)
	) name14879 (
		_w3214_,
		_w11388_,
		_w14913_
	);
	LUT4 #(
		.INIT('h2228)
	) name14880 (
		_w3249_,
		_w7935_,
		_w8077_,
		_w11279_,
		_w14914_
	);
	LUT2 #(
		.INIT('h1)
	) name14881 (
		_w14913_,
		_w14914_,
		_w14915_
	);
	LUT2 #(
		.INIT('h4)
	) name14882 (
		_w14912_,
		_w14915_,
		_w14916_
	);
	LUT3 #(
		.INIT('h9a)
	) name14883 (
		\a[23] ,
		_w14911_,
		_w14916_,
		_w14917_
	);
	LUT3 #(
		.INIT('h96)
	) name14884 (
		_w14864_,
		_w14910_,
		_w14917_,
		_w14918_
	);
	LUT3 #(
		.INIT('h82)
	) name14885 (
		_w3312_,
		_w11490_,
		_w11492_,
		_w14919_
	);
	LUT3 #(
		.INIT('h82)
	) name14886 (
		_w3654_,
		_w11286_,
		_w11335_,
		_w14920_
	);
	LUT2 #(
		.INIT('h8)
	) name14887 (
		_w3311_,
		_w11382_,
		_w14921_
	);
	LUT4 #(
		.INIT('h2228)
	) name14888 (
		_w3645_,
		_w7695_,
		_w7750_,
		_w11285_,
		_w14922_
	);
	LUT2 #(
		.INIT('h1)
	) name14889 (
		_w14921_,
		_w14922_,
		_w14923_
	);
	LUT2 #(
		.INIT('h4)
	) name14890 (
		_w14920_,
		_w14923_,
		_w14924_
	);
	LUT3 #(
		.INIT('h9a)
	) name14891 (
		\a[20] ,
		_w14919_,
		_w14924_,
		_w14925_
	);
	LUT4 #(
		.INIT('h2882)
	) name14892 (
		_w14862_,
		_w14863_,
		_w14918_,
		_w14925_,
		_w14926_
	);
	LUT4 #(
		.INIT('h4114)
	) name14893 (
		_w14862_,
		_w14863_,
		_w14918_,
		_w14925_,
		_w14927_
	);
	LUT4 #(
		.INIT('h9669)
	) name14894 (
		_w14862_,
		_w14863_,
		_w14918_,
		_w14925_,
		_w14928_
	);
	LUT3 #(
		.INIT('h82)
	) name14895 (
		_w3710_,
		_w13061_,
		_w13102_,
		_w14929_
	);
	LUT3 #(
		.INIT('h82)
	) name14896 (
		_w3886_,
		_w13062_,
		_w13099_,
		_w14930_
	);
	LUT2 #(
		.INIT('h8)
	) name14897 (
		_w3709_,
		_w11377_,
		_w14931_
	);
	LUT4 #(
		.INIT('h2228)
	) name14898 (
		_w3877_,
		_w11549_,
		_w11373_,
		_w11375_,
		_w14932_
	);
	LUT2 #(
		.INIT('h1)
	) name14899 (
		_w14931_,
		_w14932_,
		_w14933_
	);
	LUT2 #(
		.INIT('h4)
	) name14900 (
		_w14930_,
		_w14933_,
		_w14934_
	);
	LUT3 #(
		.INIT('h9a)
	) name14901 (
		\a[17] ,
		_w14929_,
		_w14934_,
		_w14935_
	);
	LUT3 #(
		.INIT('h82)
	) name14902 (
		_w4034_,
		_w13292_,
		_w13325_,
		_w14936_
	);
	LUT3 #(
		.INIT('h82)
	) name14903 (
		_w4382_,
		_w13293_,
		_w13322_,
		_w14937_
	);
	LUT2 #(
		.INIT('h8)
	) name14904 (
		_w4033_,
		_w13247_,
		_w14938_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14905 (
		_w4367_,
		_w13243_,
		_w13245_,
		_w13285_,
		_w14939_
	);
	LUT2 #(
		.INIT('h1)
	) name14906 (
		_w14938_,
		_w14939_,
		_w14940_
	);
	LUT2 #(
		.INIT('h4)
	) name14907 (
		_w14937_,
		_w14940_,
		_w14941_
	);
	LUT3 #(
		.INIT('h9a)
	) name14908 (
		\a[14] ,
		_w14936_,
		_w14941_,
		_w14942_
	);
	LUT4 #(
		.INIT('h9669)
	) name14909 (
		_w14861_,
		_w14928_,
		_w14935_,
		_w14942_,
		_w14943_
	);
	LUT4 #(
		.INIT('h2882)
	) name14910 (
		_w14852_,
		_w14859_,
		_w14860_,
		_w14943_,
		_w14944_
	);
	LUT4 #(
		.INIT('h4114)
	) name14911 (
		_w14852_,
		_w14859_,
		_w14860_,
		_w14943_,
		_w14945_
	);
	LUT4 #(
		.INIT('h9669)
	) name14912 (
		_w14852_,
		_w14859_,
		_w14860_,
		_w14943_,
		_w14946_
	);
	LUT3 #(
		.INIT('h82)
	) name14913 (
		_w4876_,
		_w14343_,
		_w14349_,
		_w14947_
	);
	LUT3 #(
		.INIT('h28)
	) name14914 (
		_w5286_,
		_w14344_,
		_w14347_,
		_w14948_
	);
	LUT2 #(
		.INIT('h8)
	) name14915 (
		_w4875_,
		_w14112_,
		_w14949_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14916 (
		_w5271_,
		_w14108_,
		_w14111_,
		_w14235_,
		_w14950_
	);
	LUT2 #(
		.INIT('h1)
	) name14917 (
		_w14949_,
		_w14950_,
		_w14951_
	);
	LUT2 #(
		.INIT('h4)
	) name14918 (
		_w14948_,
		_w14951_,
		_w14952_
	);
	LUT3 #(
		.INIT('h9a)
	) name14919 (
		\a[8] ,
		_w14947_,
		_w14952_,
		_w14953_
	);
	LUT3 #(
		.INIT('h41)
	) name14920 (
		_w14851_,
		_w14946_,
		_w14953_,
		_w14954_
	);
	LUT3 #(
		.INIT('h96)
	) name14921 (
		_w14851_,
		_w14946_,
		_w14953_,
		_w14955_
	);
	LUT4 #(
		.INIT('hd400)
	) name14922 (
		_w14757_,
		_w14844_,
		_w14845_,
		_w14955_,
		_w14956_
	);
	LUT4 #(
		.INIT('h32cd)
	) name14923 (
		_w14757_,
		_w14846_,
		_w14847_,
		_w14955_,
		_w14957_
	);
	LUT2 #(
		.INIT('h8)
	) name14924 (
		_w14849_,
		_w14957_,
		_w14958_
	);
	LUT2 #(
		.INIT('h6)
	) name14925 (
		_w14849_,
		_w14957_,
		_w14959_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name14926 (
		_w4876_,
		_w14343_,
		_w14348_,
		_w14349_,
		_w14960_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14927 (
		_w4875_,
		_w14108_,
		_w14111_,
		_w14235_,
		_w14961_
	);
	LUT4 #(
		.INIT('h00d7)
	) name14928 (
		_w8996_,
		_w14344_,
		_w14347_,
		_w14961_,
		_w14962_
	);
	LUT3 #(
		.INIT('h9a)
	) name14929 (
		\a[8] ,
		_w14960_,
		_w14962_,
		_w14963_
	);
	LUT4 #(
		.INIT('h0071)
	) name14930 (
		_w14859_,
		_w14860_,
		_w14943_,
		_w14963_,
		_w14964_
	);
	LUT4 #(
		.INIT('h8e00)
	) name14931 (
		_w14859_,
		_w14860_,
		_w14943_,
		_w14963_,
		_w14965_
	);
	LUT4 #(
		.INIT('h718e)
	) name14932 (
		_w14859_,
		_w14860_,
		_w14943_,
		_w14963_,
		_w14966_
	);
	LUT4 #(
		.INIT('h2228)
	) name14933 (
		_w2874_,
		_w8466_,
		_w8541_,
		_w11273_,
		_w14967_
	);
	LUT4 #(
		.INIT('h007d)
	) name14934 (
		_w2975_,
		_w11274_,
		_w11276_,
		_w14967_,
		_w14968_
	);
	LUT3 #(
		.INIT('h70)
	) name14935 (
		_w2986_,
		_w11388_,
		_w14968_,
		_w14969_
	);
	LUT4 #(
		.INIT('h95aa)
	) name14936 (
		\a[26] ,
		_w2875_,
		_w12391_,
		_w14969_,
		_w14970_
	);
	LUT4 #(
		.INIT('h135f)
	) name14937 (
		_w122_,
		_w93_,
		_w46_,
		_w201_,
		_w14971_
	);
	LUT4 #(
		.INIT('h4000)
	) name14938 (
		_w79_,
		_w348_,
		_w1198_,
		_w14971_,
		_w14972_
	);
	LUT4 #(
		.INIT('h1000)
	) name14939 (
		_w69_,
		_w51_,
		_w2477_,
		_w3109_,
		_w14973_
	);
	LUT3 #(
		.INIT('h80)
	) name14940 (
		_w1688_,
		_w2086_,
		_w2517_,
		_w14974_
	);
	LUT4 #(
		.INIT('h8000)
	) name14941 (
		_w1219_,
		_w14974_,
		_w14972_,
		_w14973_,
		_w14975_
	);
	LUT2 #(
		.INIT('h8)
	) name14942 (
		_w2062_,
		_w14975_,
		_w14976_
	);
	LUT4 #(
		.INIT('h135f)
	) name14943 (
		_w106_,
		_w52_,
		_w90_,
		_w259_,
		_w14977_
	);
	LUT2 #(
		.INIT('h4)
	) name14944 (
		_w398_,
		_w14977_,
		_w14978_
	);
	LUT4 #(
		.INIT('h153f)
	) name14945 (
		_w56_,
		_w43_,
		_w93_,
		_w166_,
		_w14979_
	);
	LUT3 #(
		.INIT('h80)
	) name14946 (
		_w1287_,
		_w2223_,
		_w14979_,
		_w14980_
	);
	LUT2 #(
		.INIT('h8)
	) name14947 (
		_w14978_,
		_w14980_,
		_w14981_
	);
	LUT3 #(
		.INIT('h57)
	) name14948 (
		_w90_,
		_w39_,
		_w201_,
		_w14982_
	);
	LUT4 #(
		.INIT('h135f)
	) name14949 (
		_w52_,
		_w67_,
		_w419_,
		_w430_,
		_w14983_
	);
	LUT4 #(
		.INIT('h8000)
	) name14950 (
		_w138_,
		_w3510_,
		_w14982_,
		_w14983_,
		_w14984_
	);
	LUT4 #(
		.INIT('h4000)
	) name14951 (
		_w390_,
		_w976_,
		_w2654_,
		_w4170_,
		_w14985_
	);
	LUT4 #(
		.INIT('h8000)
	) name14952 (
		_w2730_,
		_w2732_,
		_w14984_,
		_w14985_,
		_w14986_
	);
	LUT3 #(
		.INIT('h80)
	) name14953 (
		_w2693_,
		_w14981_,
		_w14986_,
		_w14987_
	);
	LUT3 #(
		.INIT('h80)
	) name14954 (
		_w7324_,
		_w14976_,
		_w14987_,
		_w14988_
	);
	LUT4 #(
		.INIT('h817e)
	) name14955 (
		_w14866_,
		_w14881_,
		_w14889_,
		_w14988_,
		_w14989_
	);
	LUT4 #(
		.INIT('h2228)
	) name14956 (
		_w376_,
		_w9446_,
		_w9702_,
		_w11261_,
		_w14990_
	);
	LUT4 #(
		.INIT('h007d)
	) name14957 (
		_w2407_,
		_w11262_,
		_w11264_,
		_w14990_,
		_w14991_
	);
	LUT3 #(
		.INIT('h70)
	) name14958 (
		_w2527_,
		_w11400_,
		_w14991_,
		_w14992_
	);
	LUT3 #(
		.INIT('h70)
	) name14959 (
		_w377_,
		_w11967_,
		_w14992_,
		_w14993_
	);
	LUT2 #(
		.INIT('h2)
	) name14960 (
		_w14989_,
		_w14993_,
		_w14994_
	);
	LUT2 #(
		.INIT('h9)
	) name14961 (
		_w14989_,
		_w14993_,
		_w14995_
	);
	LUT4 #(
		.INIT('h4d00)
	) name14962 (
		_w14865_,
		_w14890_,
		_w14900_,
		_w14995_,
		_w14996_
	);
	LUT4 #(
		.INIT('h32cd)
	) name14963 (
		_w14891_,
		_w14892_,
		_w14900_,
		_w14995_,
		_w14997_
	);
	LUT4 #(
		.INIT('h2228)
	) name14964 (
		_w2549_,
		_w8794_,
		_w8994_,
		_w11267_,
		_w14998_
	);
	LUT4 #(
		.INIT('h007d)
	) name14965 (
		_w2617_,
		_w11268_,
		_w11270_,
		_w14998_,
		_w14999_
	);
	LUT3 #(
		.INIT('h70)
	) name14966 (
		_w2854_,
		_w11394_,
		_w14999_,
		_w15000_
	);
	LUT4 #(
		.INIT('h95aa)
	) name14967 (
		\a[29] ,
		_w2550_,
		_w12209_,
		_w15000_,
		_w15001_
	);
	LUT3 #(
		.INIT('h96)
	) name14968 (
		_w14970_,
		_w14997_,
		_w15001_,
		_w15002_
	);
	LUT3 #(
		.INIT('h8e)
	) name14969 (
		_w14901_,
		_w14902_,
		_w14909_,
		_w15003_
	);
	LUT4 #(
		.INIT('h2228)
	) name14970 (
		_w3214_,
		_w7935_,
		_w8077_,
		_w11279_,
		_w15004_
	);
	LUT4 #(
		.INIT('h007d)
	) name14971 (
		_w3249_,
		_w11280_,
		_w11282_,
		_w15004_,
		_w15005_
	);
	LUT3 #(
		.INIT('h70)
	) name14972 (
		_w3262_,
		_w11382_,
		_w15005_,
		_w15006_
	);
	LUT4 #(
		.INIT('h95aa)
	) name14973 (
		\a[23] ,
		_w37_,
		_w12476_,
		_w15006_,
		_w15007_
	);
	LUT3 #(
		.INIT('h69)
	) name14974 (
		_w15002_,
		_w15003_,
		_w15007_,
		_w15008_
	);
	LUT3 #(
		.INIT('h4d)
	) name14975 (
		_w14864_,
		_w14910_,
		_w14917_,
		_w15009_
	);
	LUT4 #(
		.INIT('h2228)
	) name14976 (
		_w3311_,
		_w7695_,
		_w7750_,
		_w11285_,
		_w15010_
	);
	LUT4 #(
		.INIT('h007d)
	) name14977 (
		_w3645_,
		_w11286_,
		_w11335_,
		_w15010_,
		_w15011_
	);
	LUT3 #(
		.INIT('h70)
	) name14978 (
		_w3654_,
		_w11377_,
		_w15011_,
		_w15012_
	);
	LUT4 #(
		.INIT('h95aa)
	) name14979 (
		\a[20] ,
		_w3312_,
		_w12799_,
		_w15012_,
		_w15013_
	);
	LUT3 #(
		.INIT('h69)
	) name14980 (
		_w15008_,
		_w15009_,
		_w15013_,
		_w15014_
	);
	LUT3 #(
		.INIT('h4d)
	) name14981 (
		_w14863_,
		_w14918_,
		_w14925_,
		_w15015_
	);
	LUT4 #(
		.INIT('h2228)
	) name14982 (
		_w3709_,
		_w11549_,
		_w11373_,
		_w11375_,
		_w15016_
	);
	LUT4 #(
		.INIT('h007d)
	) name14983 (
		_w3877_,
		_w13062_,
		_w13099_,
		_w15016_,
		_w15017_
	);
	LUT3 #(
		.INIT('h70)
	) name14984 (
		_w3886_,
		_w13247_,
		_w15017_,
		_w15018_
	);
	LUT4 #(
		.INIT('h95aa)
	) name14985 (
		\a[17] ,
		_w3710_,
		_w13576_,
		_w15018_,
		_w15019_
	);
	LUT3 #(
		.INIT('h69)
	) name14986 (
		_w15014_,
		_w15015_,
		_w15019_,
		_w15020_
	);
	LUT3 #(
		.INIT('h45)
	) name14987 (
		_w14926_,
		_w14927_,
		_w14935_,
		_w15021_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14988 (
		_w4033_,
		_w13243_,
		_w13245_,
		_w13285_,
		_w15022_
	);
	LUT4 #(
		.INIT('h007d)
	) name14989 (
		_w4367_,
		_w13293_,
		_w13322_,
		_w15022_,
		_w15023_
	);
	LUT3 #(
		.INIT('h70)
	) name14990 (
		_w4382_,
		_w13716_,
		_w15023_,
		_w15024_
	);
	LUT4 #(
		.INIT('h95aa)
	) name14991 (
		\a[14] ,
		_w4034_,
		_w13720_,
		_w15024_,
		_w15025_
	);
	LUT3 #(
		.INIT('h69)
	) name14992 (
		_w15020_,
		_w15021_,
		_w15025_,
		_w15026_
	);
	LUT4 #(
		.INIT('h41d7)
	) name14993 (
		_w14861_,
		_w14928_,
		_w14935_,
		_w14942_,
		_w15027_
	);
	LUT4 #(
		.INIT('h0096)
	) name14994 (
		_w15020_,
		_w15021_,
		_w15025_,
		_w15027_,
		_w15028_
	);
	LUT4 #(
		.INIT('h6900)
	) name14995 (
		_w15020_,
		_w15021_,
		_w15025_,
		_w15027_,
		_w15029_
	);
	LUT4 #(
		.INIT('h9669)
	) name14996 (
		_w15020_,
		_w15021_,
		_w15025_,
		_w15027_,
		_w15030_
	);
	LUT4 #(
		.INIT('h02a8)
	) name14997 (
		_w4458_,
		_w13712_,
		_w13714_,
		_w13847_,
		_w15031_
	);
	LUT4 #(
		.INIT('h007d)
	) name14998 (
		_w4684_,
		_w13960_,
		_w13979_,
		_w15031_,
		_w15032_
	);
	LUT3 #(
		.INIT('h70)
	) name14999 (
		_w4700_,
		_w14112_,
		_w15032_,
		_w15033_
	);
	LUT4 #(
		.INIT('h95aa)
	) name15000 (
		\a[11] ,
		_w4459_,
		_w14116_,
		_w15033_,
		_w15034_
	);
	LUT3 #(
		.INIT('h69)
	) name15001 (
		_w14966_,
		_w15030_,
		_w15034_,
		_w15035_
	);
	LUT3 #(
		.INIT('h45)
	) name15002 (
		_w14944_,
		_w14945_,
		_w14953_,
		_w15036_
	);
	LUT2 #(
		.INIT('h8)
	) name15003 (
		_w15035_,
		_w15036_,
		_w15037_
	);
	LUT2 #(
		.INIT('h6)
	) name15004 (
		_w15035_,
		_w15036_,
		_w15038_
	);
	LUT3 #(
		.INIT('h1e)
	) name15005 (
		_w14954_,
		_w14956_,
		_w15038_,
		_w15039_
	);
	LUT2 #(
		.INIT('h6)
	) name15006 (
		_w14958_,
		_w15039_,
		_w15040_
	);
	LUT4 #(
		.INIT('h010f)
	) name15007 (
		_w14954_,
		_w14956_,
		_w15037_,
		_w15038_,
		_w15041_
	);
	LUT3 #(
		.INIT('hb2)
	) name15008 (
		_w14970_,
		_w14997_,
		_w15001_,
		_w15042_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15009 (
		_w2550_,
		_w11396_,
		_w11476_,
		_w11477_,
		_w15043_
	);
	LUT4 #(
		.INIT('h2228)
	) name15010 (
		_w2854_,
		_w8466_,
		_w8541_,
		_w11273_,
		_w15044_
	);
	LUT3 #(
		.INIT('h82)
	) name15011 (
		_w2549_,
		_w11268_,
		_w11270_,
		_w15045_
	);
	LUT3 #(
		.INIT('h07)
	) name15012 (
		_w2617_,
		_w11394_,
		_w15045_,
		_w15046_
	);
	LUT2 #(
		.INIT('h4)
	) name15013 (
		_w15044_,
		_w15046_,
		_w15047_
	);
	LUT3 #(
		.INIT('h9a)
	) name15014 (
		\a[29] ,
		_w15043_,
		_w15047_,
		_w15048_
	);
	LUT4 #(
		.INIT('hb332)
	) name15015 (
		_w14866_,
		_w14881_,
		_w14889_,
		_w14988_,
		_w15049_
	);
	LUT4 #(
		.INIT('h5665)
	) name15016 (
		\a[8] ,
		_w7633_,
		_w14344_,
		_w14347_,
		_w15050_
	);
	LUT4 #(
		.INIT('h4000)
	) name15017 (
		_w186_,
		_w971_,
		_w1523_,
		_w1524_,
		_w15051_
	);
	LUT2 #(
		.INIT('h8)
	) name15018 (
		_w7316_,
		_w15051_,
		_w15052_
	);
	LUT3 #(
		.INIT('h80)
	) name15019 (
		_w760_,
		_w960_,
		_w1275_,
		_w15053_
	);
	LUT4 #(
		.INIT('h135f)
	) name15020 (
		_w122_,
		_w110_,
		_w67_,
		_w378_,
		_w15054_
	);
	LUT4 #(
		.INIT('h8000)
	) name15021 (
		_w260_,
		_w820_,
		_w821_,
		_w15054_,
		_w15055_
	);
	LUT3 #(
		.INIT('h80)
	) name15022 (
		_w7304_,
		_w15053_,
		_w15055_,
		_w15056_
	);
	LUT3 #(
		.INIT('h80)
	) name15023 (
		_w1851_,
		_w15052_,
		_w15056_,
		_w15057_
	);
	LUT4 #(
		.INIT('h8000)
	) name15024 (
		_w881_,
		_w897_,
		_w2269_,
		_w2272_,
		_w15058_
	);
	LUT4 #(
		.INIT('h8000)
	) name15025 (
		_w1009_,
		_w14880_,
		_w15057_,
		_w15058_,
		_w15059_
	);
	LUT4 #(
		.INIT('h0777)
	) name15026 (
		_w1009_,
		_w14880_,
		_w15057_,
		_w15058_,
		_w15060_
	);
	LUT4 #(
		.INIT('h7888)
	) name15027 (
		_w1009_,
		_w14880_,
		_w15057_,
		_w15058_,
		_w15061_
	);
	LUT2 #(
		.INIT('h6)
	) name15028 (
		_w15050_,
		_w15061_,
		_w15062_
	);
	LUT3 #(
		.INIT('h82)
	) name15029 (
		_w377_,
		_w11469_,
		_w11471_,
		_w15063_
	);
	LUT4 #(
		.INIT('h2228)
	) name15030 (
		_w2527_,
		_w8794_,
		_w8994_,
		_w11267_,
		_w15064_
	);
	LUT3 #(
		.INIT('h82)
	) name15031 (
		_w376_,
		_w11262_,
		_w11264_,
		_w15065_
	);
	LUT3 #(
		.INIT('h07)
	) name15032 (
		_w2407_,
		_w11400_,
		_w15065_,
		_w15066_
	);
	LUT2 #(
		.INIT('h4)
	) name15033 (
		_w15064_,
		_w15066_,
		_w15067_
	);
	LUT2 #(
		.INIT('h4)
	) name15034 (
		_w15063_,
		_w15067_,
		_w15068_
	);
	LUT4 #(
		.INIT('h4114)
	) name15035 (
		_w15048_,
		_w15049_,
		_w15062_,
		_w15068_,
		_w15069_
	);
	LUT4 #(
		.INIT('h9669)
	) name15036 (
		_w15048_,
		_w15049_,
		_w15062_,
		_w15068_,
		_w15070_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15037 (
		_w2875_,
		_w11390_,
		_w11482_,
		_w11483_,
		_w15071_
	);
	LUT4 #(
		.INIT('h2228)
	) name15038 (
		_w2986_,
		_w7935_,
		_w8077_,
		_w11279_,
		_w15072_
	);
	LUT3 #(
		.INIT('h82)
	) name15039 (
		_w2874_,
		_w11274_,
		_w11276_,
		_w15073_
	);
	LUT3 #(
		.INIT('h07)
	) name15040 (
		_w2975_,
		_w11388_,
		_w15073_,
		_w15074_
	);
	LUT2 #(
		.INIT('h4)
	) name15041 (
		_w15072_,
		_w15074_,
		_w15075_
	);
	LUT3 #(
		.INIT('h9a)
	) name15042 (
		\a[26] ,
		_w15071_,
		_w15075_,
		_w15076_
	);
	LUT4 #(
		.INIT('h001e)
	) name15043 (
		_w14994_,
		_w14996_,
		_w15070_,
		_w15076_,
		_w15077_
	);
	LUT4 #(
		.INIT('he100)
	) name15044 (
		_w14994_,
		_w14996_,
		_w15070_,
		_w15076_,
		_w15078_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name15045 (
		_w14994_,
		_w14996_,
		_w15070_,
		_w15076_,
		_w15079_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15046 (
		_w37_,
		_w11384_,
		_w11488_,
		_w11489_,
		_w15080_
	);
	LUT4 #(
		.INIT('h2228)
	) name15047 (
		_w3262_,
		_w7695_,
		_w7750_,
		_w11285_,
		_w15081_
	);
	LUT3 #(
		.INIT('h82)
	) name15048 (
		_w3214_,
		_w11280_,
		_w11282_,
		_w15082_
	);
	LUT3 #(
		.INIT('h07)
	) name15049 (
		_w3249_,
		_w11382_,
		_w15082_,
		_w15083_
	);
	LUT2 #(
		.INIT('h4)
	) name15050 (
		_w15081_,
		_w15083_,
		_w15084_
	);
	LUT3 #(
		.INIT('h9a)
	) name15051 (
		\a[23] ,
		_w15080_,
		_w15084_,
		_w15085_
	);
	LUT3 #(
		.INIT('h09)
	) name15052 (
		_w15042_,
		_w15079_,
		_w15085_,
		_w15086_
	);
	LUT3 #(
		.INIT('h60)
	) name15053 (
		_w15042_,
		_w15079_,
		_w15085_,
		_w15087_
	);
	LUT3 #(
		.INIT('h96)
	) name15054 (
		_w15042_,
		_w15079_,
		_w15085_,
		_w15088_
	);
	LUT3 #(
		.INIT('h8e)
	) name15055 (
		_w15002_,
		_w15003_,
		_w15007_,
		_w15089_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15056 (
		_w3312_,
		_w11378_,
		_w11494_,
		_w11552_,
		_w15090_
	);
	LUT4 #(
		.INIT('h2228)
	) name15057 (
		_w3654_,
		_w11549_,
		_w11373_,
		_w11375_,
		_w15091_
	);
	LUT3 #(
		.INIT('h82)
	) name15058 (
		_w3311_,
		_w11286_,
		_w11335_,
		_w15092_
	);
	LUT3 #(
		.INIT('h07)
	) name15059 (
		_w3645_,
		_w11377_,
		_w15092_,
		_w15093_
	);
	LUT2 #(
		.INIT('h4)
	) name15060 (
		_w15091_,
		_w15093_,
		_w15094_
	);
	LUT3 #(
		.INIT('h9a)
	) name15061 (
		\a[20] ,
		_w15090_,
		_w15094_,
		_w15095_
	);
	LUT3 #(
		.INIT('h06)
	) name15062 (
		_w15088_,
		_w15089_,
		_w15095_,
		_w15096_
	);
	LUT3 #(
		.INIT('h90)
	) name15063 (
		_w15088_,
		_w15089_,
		_w15095_,
		_w15097_
	);
	LUT3 #(
		.INIT('h69)
	) name15064 (
		_w15088_,
		_w15089_,
		_w15095_,
		_w15098_
	);
	LUT3 #(
		.INIT('h8e)
	) name15065 (
		_w15008_,
		_w15009_,
		_w15013_,
		_w15099_
	);
	LUT2 #(
		.INIT('h6)
	) name15066 (
		_w15098_,
		_w15099_,
		_w15100_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15067 (
		_w3710_,
		_w13288_,
		_w13290_,
		_w13291_,
		_w15101_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15068 (
		_w3886_,
		_w13243_,
		_w13245_,
		_w13285_,
		_w15102_
	);
	LUT3 #(
		.INIT('h82)
	) name15069 (
		_w3709_,
		_w13062_,
		_w13099_,
		_w15103_
	);
	LUT3 #(
		.INIT('h07)
	) name15070 (
		_w3877_,
		_w13247_,
		_w15103_,
		_w15104_
	);
	LUT2 #(
		.INIT('h4)
	) name15071 (
		_w15102_,
		_w15104_,
		_w15105_
	);
	LUT3 #(
		.INIT('h9a)
	) name15072 (
		\a[17] ,
		_w15101_,
		_w15105_,
		_w15106_
	);
	LUT4 #(
		.INIT('h008e)
	) name15073 (
		_w15014_,
		_w15015_,
		_w15019_,
		_w15106_,
		_w15107_
	);
	LUT4 #(
		.INIT('h7100)
	) name15074 (
		_w15014_,
		_w15015_,
		_w15019_,
		_w15106_,
		_w15108_
	);
	LUT4 #(
		.INIT('h8e71)
	) name15075 (
		_w15014_,
		_w15015_,
		_w15019_,
		_w15106_,
		_w15109_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15076 (
		_w4034_,
		_w13717_,
		_w13719_,
		_w13850_,
		_w15110_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15077 (
		_w4382_,
		_w13712_,
		_w13714_,
		_w13847_,
		_w15111_
	);
	LUT3 #(
		.INIT('h82)
	) name15078 (
		_w4033_,
		_w13293_,
		_w13322_,
		_w15112_
	);
	LUT3 #(
		.INIT('h07)
	) name15079 (
		_w4367_,
		_w13716_,
		_w15112_,
		_w15113_
	);
	LUT2 #(
		.INIT('h4)
	) name15080 (
		_w15111_,
		_w15113_,
		_w15114_
	);
	LUT3 #(
		.INIT('h9a)
	) name15081 (
		\a[14] ,
		_w15110_,
		_w15114_,
		_w15115_
	);
	LUT3 #(
		.INIT('h06)
	) name15082 (
		_w15100_,
		_w15109_,
		_w15115_,
		_w15116_
	);
	LUT3 #(
		.INIT('h90)
	) name15083 (
		_w15100_,
		_w15109_,
		_w15115_,
		_w15117_
	);
	LUT3 #(
		.INIT('h69)
	) name15084 (
		_w15100_,
		_w15109_,
		_w15115_,
		_w15118_
	);
	LUT3 #(
		.INIT('h8e)
	) name15085 (
		_w15020_,
		_w15021_,
		_w15025_,
		_w15119_
	);
	LUT2 #(
		.INIT('h6)
	) name15086 (
		_w15118_,
		_w15119_,
		_w15120_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15087 (
		_w4459_,
		_w14113_,
		_w14115_,
		_w14238_,
		_w15121_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15088 (
		_w4700_,
		_w14108_,
		_w14111_,
		_w14235_,
		_w15122_
	);
	LUT3 #(
		.INIT('h82)
	) name15089 (
		_w4458_,
		_w13960_,
		_w13979_,
		_w15123_
	);
	LUT3 #(
		.INIT('h07)
	) name15090 (
		_w4684_,
		_w14112_,
		_w15123_,
		_w15124_
	);
	LUT2 #(
		.INIT('h4)
	) name15091 (
		_w15122_,
		_w15124_,
		_w15125_
	);
	LUT3 #(
		.INIT('h9a)
	) name15092 (
		\a[11] ,
		_w15121_,
		_w15125_,
		_w15126_
	);
	LUT4 #(
		.INIT('h008e)
	) name15093 (
		_w15026_,
		_w15027_,
		_w15034_,
		_w15126_,
		_w15127_
	);
	LUT4 #(
		.INIT('h7100)
	) name15094 (
		_w15026_,
		_w15027_,
		_w15034_,
		_w15126_,
		_w15128_
	);
	LUT4 #(
		.INIT('h45ba)
	) name15095 (
		_w15028_,
		_w15029_,
		_w15034_,
		_w15126_,
		_w15129_
	);
	LUT4 #(
		.INIT('h3223)
	) name15096 (
		_w14964_,
		_w14965_,
		_w15030_,
		_w15034_,
		_w15130_
	);
	LUT3 #(
		.INIT('h60)
	) name15097 (
		_w15120_,
		_w15129_,
		_w15130_,
		_w15131_
	);
	LUT3 #(
		.INIT('h09)
	) name15098 (
		_w15120_,
		_w15129_,
		_w15130_,
		_w15132_
	);
	LUT3 #(
		.INIT('h96)
	) name15099 (
		_w15120_,
		_w15129_,
		_w15130_,
		_w15133_
	);
	LUT4 #(
		.INIT('h8008)
	) name15100 (
		_w14958_,
		_w15039_,
		_w15041_,
		_w15133_,
		_w15134_
	);
	LUT4 #(
		.INIT('h7887)
	) name15101 (
		_w14958_,
		_w15039_,
		_w15041_,
		_w15133_,
		_w15135_
	);
	LUT3 #(
		.INIT('h31)
	) name15102 (
		_w15120_,
		_w15127_,
		_w15128_,
		_w15136_
	);
	LUT3 #(
		.INIT('h45)
	) name15103 (
		_w15116_,
		_w15117_,
		_w15119_,
		_w15137_
	);
	LUT3 #(
		.INIT('h82)
	) name15104 (
		_w4034_,
		_w13959_,
		_w13982_,
		_w15138_
	);
	LUT3 #(
		.INIT('h82)
	) name15105 (
		_w4382_,
		_w13960_,
		_w13979_,
		_w15139_
	);
	LUT2 #(
		.INIT('h8)
	) name15106 (
		_w4033_,
		_w13716_,
		_w15140_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15107 (
		_w4367_,
		_w13712_,
		_w13714_,
		_w13847_,
		_w15141_
	);
	LUT2 #(
		.INIT('h1)
	) name15108 (
		_w15140_,
		_w15141_,
		_w15142_
	);
	LUT2 #(
		.INIT('h4)
	) name15109 (
		_w15139_,
		_w15142_,
		_w15143_
	);
	LUT3 #(
		.INIT('h9a)
	) name15110 (
		\a[14] ,
		_w15138_,
		_w15143_,
		_w15144_
	);
	LUT3 #(
		.INIT('h31)
	) name15111 (
		_w15100_,
		_w15107_,
		_w15108_,
		_w15145_
	);
	LUT3 #(
		.INIT('h45)
	) name15112 (
		_w15096_,
		_w15097_,
		_w15099_,
		_w15146_
	);
	LUT3 #(
		.INIT('h45)
	) name15113 (
		_w15086_,
		_w15087_,
		_w15089_,
		_w15147_
	);
	LUT3 #(
		.INIT('h32)
	) name15114 (
		_w15042_,
		_w15077_,
		_w15078_,
		_w15148_
	);
	LUT4 #(
		.INIT('h010f)
	) name15115 (
		_w14994_,
		_w14996_,
		_w15069_,
		_w15070_,
		_w15149_
	);
	LUT3 #(
		.INIT('h0d)
	) name15116 (
		_w15050_,
		_w15059_,
		_w15060_,
		_w15150_
	);
	LUT4 #(
		.INIT('h153f)
	) name15117 (
		_w56_,
		_w47_,
		_w39_,
		_w259_,
		_w15151_
	);
	LUT4 #(
		.INIT('h1000)
	) name15118 (
		_w243_,
		_w412_,
		_w502_,
		_w15151_,
		_w15152_
	);
	LUT4 #(
		.INIT('h1000)
	) name15119 (
		_w338_,
		_w426_,
		_w7997_,
		_w8263_,
		_w15153_
	);
	LUT4 #(
		.INIT('h8000)
	) name15120 (
		_w1276_,
		_w1557_,
		_w2198_,
		_w2468_,
		_w15154_
	);
	LUT4 #(
		.INIT('h8000)
	) name15121 (
		_w3334_,
		_w15154_,
		_w15152_,
		_w15153_,
		_w15155_
	);
	LUT4 #(
		.INIT('h8000)
	) name15122 (
		_w730_,
		_w741_,
		_w7535_,
		_w15155_,
		_w15156_
	);
	LUT2 #(
		.INIT('h8)
	) name15123 (
		_w1692_,
		_w15156_,
		_w15157_
	);
	LUT4 #(
		.INIT('h0df2)
	) name15124 (
		_w15050_,
		_w15059_,
		_w15060_,
		_w15157_,
		_w15158_
	);
	LUT3 #(
		.INIT('h82)
	) name15125 (
		_w377_,
		_w11472_,
		_w11474_,
		_w15159_
	);
	LUT3 #(
		.INIT('h82)
	) name15126 (
		_w2527_,
		_w11268_,
		_w11270_,
		_w15160_
	);
	LUT2 #(
		.INIT('h8)
	) name15127 (
		_w376_,
		_w11400_,
		_w15161_
	);
	LUT4 #(
		.INIT('h2228)
	) name15128 (
		_w2407_,
		_w8794_,
		_w8994_,
		_w11267_,
		_w15162_
	);
	LUT2 #(
		.INIT('h1)
	) name15129 (
		_w15161_,
		_w15162_,
		_w15163_
	);
	LUT2 #(
		.INIT('h4)
	) name15130 (
		_w15160_,
		_w15163_,
		_w15164_
	);
	LUT2 #(
		.INIT('h4)
	) name15131 (
		_w15159_,
		_w15164_,
		_w15165_
	);
	LUT2 #(
		.INIT('h9)
	) name15132 (
		_w15158_,
		_w15165_,
		_w15166_
	);
	LUT3 #(
		.INIT('h4d)
	) name15133 (
		_w15049_,
		_w15062_,
		_w15068_,
		_w15167_
	);
	LUT4 #(
		.INIT('h00b2)
	) name15134 (
		_w15049_,
		_w15062_,
		_w15068_,
		_w15166_,
		_w15168_
	);
	LUT4 #(
		.INIT('h4d00)
	) name15135 (
		_w15049_,
		_w15062_,
		_w15068_,
		_w15166_,
		_w15169_
	);
	LUT4 #(
		.INIT('hb24d)
	) name15136 (
		_w15049_,
		_w15062_,
		_w15068_,
		_w15166_,
		_w15170_
	);
	LUT3 #(
		.INIT('h82)
	) name15137 (
		_w2550_,
		_w11478_,
		_w11480_,
		_w15171_
	);
	LUT3 #(
		.INIT('h82)
	) name15138 (
		_w2854_,
		_w11274_,
		_w11276_,
		_w15172_
	);
	LUT2 #(
		.INIT('h8)
	) name15139 (
		_w2549_,
		_w11394_,
		_w15173_
	);
	LUT4 #(
		.INIT('h2228)
	) name15140 (
		_w2617_,
		_w8466_,
		_w8541_,
		_w11273_,
		_w15174_
	);
	LUT2 #(
		.INIT('h1)
	) name15141 (
		_w15173_,
		_w15174_,
		_w15175_
	);
	LUT2 #(
		.INIT('h4)
	) name15142 (
		_w15172_,
		_w15175_,
		_w15176_
	);
	LUT3 #(
		.INIT('h9a)
	) name15143 (
		\a[29] ,
		_w15171_,
		_w15176_,
		_w15177_
	);
	LUT2 #(
		.INIT('h9)
	) name15144 (
		_w15170_,
		_w15177_,
		_w15178_
	);
	LUT3 #(
		.INIT('h82)
	) name15145 (
		_w2875_,
		_w11484_,
		_w11486_,
		_w15179_
	);
	LUT3 #(
		.INIT('h82)
	) name15146 (
		_w2986_,
		_w11280_,
		_w11282_,
		_w15180_
	);
	LUT2 #(
		.INIT('h8)
	) name15147 (
		_w2874_,
		_w11388_,
		_w15181_
	);
	LUT4 #(
		.INIT('h2228)
	) name15148 (
		_w2975_,
		_w7935_,
		_w8077_,
		_w11279_,
		_w15182_
	);
	LUT2 #(
		.INIT('h1)
	) name15149 (
		_w15181_,
		_w15182_,
		_w15183_
	);
	LUT2 #(
		.INIT('h4)
	) name15150 (
		_w15180_,
		_w15183_,
		_w15184_
	);
	LUT3 #(
		.INIT('h9a)
	) name15151 (
		\a[26] ,
		_w15179_,
		_w15184_,
		_w15185_
	);
	LUT3 #(
		.INIT('h96)
	) name15152 (
		_w15149_,
		_w15178_,
		_w15185_,
		_w15186_
	);
	LUT3 #(
		.INIT('h82)
	) name15153 (
		_w37_,
		_w11490_,
		_w11492_,
		_w15187_
	);
	LUT3 #(
		.INIT('h82)
	) name15154 (
		_w3262_,
		_w11286_,
		_w11335_,
		_w15188_
	);
	LUT2 #(
		.INIT('h8)
	) name15155 (
		_w3214_,
		_w11382_,
		_w15189_
	);
	LUT4 #(
		.INIT('h2228)
	) name15156 (
		_w3249_,
		_w7695_,
		_w7750_,
		_w11285_,
		_w15190_
	);
	LUT2 #(
		.INIT('h1)
	) name15157 (
		_w15189_,
		_w15190_,
		_w15191_
	);
	LUT2 #(
		.INIT('h4)
	) name15158 (
		_w15188_,
		_w15191_,
		_w15192_
	);
	LUT3 #(
		.INIT('h9a)
	) name15159 (
		\a[23] ,
		_w15187_,
		_w15192_,
		_w15193_
	);
	LUT3 #(
		.INIT('h96)
	) name15160 (
		_w15148_,
		_w15186_,
		_w15193_,
		_w15194_
	);
	LUT3 #(
		.INIT('h82)
	) name15161 (
		_w3312_,
		_w13061_,
		_w13102_,
		_w15195_
	);
	LUT3 #(
		.INIT('h82)
	) name15162 (
		_w3654_,
		_w13062_,
		_w13099_,
		_w15196_
	);
	LUT2 #(
		.INIT('h8)
	) name15163 (
		_w3311_,
		_w11377_,
		_w15197_
	);
	LUT4 #(
		.INIT('h2228)
	) name15164 (
		_w3645_,
		_w11549_,
		_w11373_,
		_w11375_,
		_w15198_
	);
	LUT2 #(
		.INIT('h1)
	) name15165 (
		_w15197_,
		_w15198_,
		_w15199_
	);
	LUT2 #(
		.INIT('h4)
	) name15166 (
		_w15196_,
		_w15199_,
		_w15200_
	);
	LUT3 #(
		.INIT('h9a)
	) name15167 (
		\a[20] ,
		_w15195_,
		_w15200_,
		_w15201_
	);
	LUT3 #(
		.INIT('h96)
	) name15168 (
		_w15147_,
		_w15194_,
		_w15201_,
		_w15202_
	);
	LUT3 #(
		.INIT('h82)
	) name15169 (
		_w3710_,
		_w13292_,
		_w13325_,
		_w15203_
	);
	LUT3 #(
		.INIT('h82)
	) name15170 (
		_w3886_,
		_w13293_,
		_w13322_,
		_w15204_
	);
	LUT2 #(
		.INIT('h8)
	) name15171 (
		_w3709_,
		_w13247_,
		_w15205_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15172 (
		_w3877_,
		_w13243_,
		_w13245_,
		_w13285_,
		_w15206_
	);
	LUT2 #(
		.INIT('h1)
	) name15173 (
		_w15205_,
		_w15206_,
		_w15207_
	);
	LUT2 #(
		.INIT('h4)
	) name15174 (
		_w15204_,
		_w15207_,
		_w15208_
	);
	LUT3 #(
		.INIT('h9a)
	) name15175 (
		\a[17] ,
		_w15203_,
		_w15208_,
		_w15209_
	);
	LUT3 #(
		.INIT('h96)
	) name15176 (
		_w15146_,
		_w15202_,
		_w15209_,
		_w15210_
	);
	LUT3 #(
		.INIT('h96)
	) name15177 (
		_w15144_,
		_w15145_,
		_w15210_,
		_w15211_
	);
	LUT3 #(
		.INIT('h82)
	) name15178 (
		_w4459_,
		_w14343_,
		_w14349_,
		_w15212_
	);
	LUT3 #(
		.INIT('h28)
	) name15179 (
		_w4700_,
		_w14344_,
		_w14347_,
		_w15213_
	);
	LUT2 #(
		.INIT('h8)
	) name15180 (
		_w4458_,
		_w14112_,
		_w15214_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15181 (
		_w4684_,
		_w14108_,
		_w14111_,
		_w14235_,
		_w15215_
	);
	LUT2 #(
		.INIT('h1)
	) name15182 (
		_w15214_,
		_w15215_,
		_w15216_
	);
	LUT2 #(
		.INIT('h4)
	) name15183 (
		_w15213_,
		_w15216_,
		_w15217_
	);
	LUT3 #(
		.INIT('h9a)
	) name15184 (
		\a[11] ,
		_w15212_,
		_w15217_,
		_w15218_
	);
	LUT3 #(
		.INIT('h96)
	) name15185 (
		_w15137_,
		_w15211_,
		_w15218_,
		_w15219_
	);
	LUT2 #(
		.INIT('h4)
	) name15186 (
		_w15136_,
		_w15219_,
		_w15220_
	);
	LUT2 #(
		.INIT('h9)
	) name15187 (
		_w15136_,
		_w15219_,
		_w15221_
	);
	LUT4 #(
		.INIT('hdc00)
	) name15188 (
		_w15041_,
		_w15131_,
		_w15133_,
		_w15221_,
		_w15222_
	);
	LUT4 #(
		.INIT('h32cd)
	) name15189 (
		_w15041_,
		_w15131_,
		_w15132_,
		_w15221_,
		_w15223_
	);
	LUT2 #(
		.INIT('h8)
	) name15190 (
		_w15134_,
		_w15223_,
		_w15224_
	);
	LUT2 #(
		.INIT('h6)
	) name15191 (
		_w15134_,
		_w15223_,
		_w15225_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name15192 (
		_w4459_,
		_w14343_,
		_w14348_,
		_w14349_,
		_w15226_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15193 (
		_w4458_,
		_w14108_,
		_w14111_,
		_w14235_,
		_w15227_
	);
	LUT4 #(
		.INIT('h00d7)
	) name15194 (
		_w8544_,
		_w14344_,
		_w14347_,
		_w15227_,
		_w15228_
	);
	LUT3 #(
		.INIT('h9a)
	) name15195 (
		\a[11] ,
		_w15226_,
		_w15228_,
		_w15229_
	);
	LUT4 #(
		.INIT('h0071)
	) name15196 (
		_w15144_,
		_w15145_,
		_w15210_,
		_w15229_,
		_w15230_
	);
	LUT4 #(
		.INIT('h8e00)
	) name15197 (
		_w15144_,
		_w15145_,
		_w15210_,
		_w15229_,
		_w15231_
	);
	LUT4 #(
		.INIT('h718e)
	) name15198 (
		_w15144_,
		_w15145_,
		_w15210_,
		_w15229_,
		_w15232_
	);
	LUT3 #(
		.INIT('h32)
	) name15199 (
		_w15168_,
		_w15169_,
		_w15177_,
		_w15233_
	);
	LUT4 #(
		.INIT('h2228)
	) name15200 (
		_w2549_,
		_w8466_,
		_w8541_,
		_w11273_,
		_w15234_
	);
	LUT4 #(
		.INIT('h007d)
	) name15201 (
		_w2617_,
		_w11274_,
		_w11276_,
		_w15234_,
		_w15235_
	);
	LUT3 #(
		.INIT('h70)
	) name15202 (
		_w2854_,
		_w11388_,
		_w15235_,
		_w15236_
	);
	LUT4 #(
		.INIT('h95aa)
	) name15203 (
		\a[29] ,
		_w2550_,
		_w12391_,
		_w15236_,
		_w15237_
	);
	LUT4 #(
		.INIT('h8000)
	) name15204 (
		_w731_,
		_w772_,
		_w1910_,
		_w2252_,
		_w15238_
	);
	LUT4 #(
		.INIT('h8000)
	) name15205 (
		_w1257_,
		_w1333_,
		_w1427_,
		_w2282_,
		_w15239_
	);
	LUT4 #(
		.INIT('h153f)
	) name15206 (
		_w38_,
		_w122_,
		_w44_,
		_w158_,
		_w15240_
	);
	LUT4 #(
		.INIT('h4000)
	) name15207 (
		_w451_,
		_w834_,
		_w1058_,
		_w15240_,
		_w15241_
	);
	LUT4 #(
		.INIT('h8000)
	) name15208 (
		_w8366_,
		_w15239_,
		_w15241_,
		_w15238_,
		_w15242_
	);
	LUT4 #(
		.INIT('h8000)
	) name15209 (
		_w7309_,
		_w7312_,
		_w7987_,
		_w7988_,
		_w15243_
	);
	LUT4 #(
		.INIT('h8000)
	) name15210 (
		_w3563_,
		_w3575_,
		_w15242_,
		_w15243_,
		_w15244_
	);
	LUT2 #(
		.INIT('h8)
	) name15211 (
		_w14872_,
		_w15244_,
		_w15245_
	);
	LUT4 #(
		.INIT('h817e)
	) name15212 (
		_w15150_,
		_w15157_,
		_w15165_,
		_w15245_,
		_w15246_
	);
	LUT4 #(
		.INIT('h2228)
	) name15213 (
		_w376_,
		_w8794_,
		_w8994_,
		_w11267_,
		_w15247_
	);
	LUT4 #(
		.INIT('h007d)
	) name15214 (
		_w2407_,
		_w11268_,
		_w11270_,
		_w15247_,
		_w15248_
	);
	LUT3 #(
		.INIT('h70)
	) name15215 (
		_w2527_,
		_w11394_,
		_w15248_,
		_w15249_
	);
	LUT3 #(
		.INIT('h70)
	) name15216 (
		_w377_,
		_w12209_,
		_w15249_,
		_w15250_
	);
	LUT3 #(
		.INIT('h96)
	) name15217 (
		_w15237_,
		_w15246_,
		_w15250_,
		_w15251_
	);
	LUT4 #(
		.INIT('h8e00)
	) name15218 (
		_w15166_,
		_w15167_,
		_w15177_,
		_w15251_,
		_w15252_
	);
	LUT4 #(
		.INIT('h0071)
	) name15219 (
		_w15166_,
		_w15167_,
		_w15177_,
		_w15251_,
		_w15253_
	);
	LUT4 #(
		.INIT('h32cd)
	) name15220 (
		_w15168_,
		_w15169_,
		_w15177_,
		_w15251_,
		_w15254_
	);
	LUT4 #(
		.INIT('h2228)
	) name15221 (
		_w2874_,
		_w7935_,
		_w8077_,
		_w11279_,
		_w15255_
	);
	LUT4 #(
		.INIT('h007d)
	) name15222 (
		_w2975_,
		_w11280_,
		_w11282_,
		_w15255_,
		_w15256_
	);
	LUT3 #(
		.INIT('h70)
	) name15223 (
		_w2986_,
		_w11382_,
		_w15256_,
		_w15257_
	);
	LUT4 #(
		.INIT('h95aa)
	) name15224 (
		\a[26] ,
		_w2875_,
		_w12476_,
		_w15257_,
		_w15258_
	);
	LUT2 #(
		.INIT('h9)
	) name15225 (
		_w15254_,
		_w15258_,
		_w15259_
	);
	LUT3 #(
		.INIT('h4d)
	) name15226 (
		_w15149_,
		_w15178_,
		_w15185_,
		_w15260_
	);
	LUT4 #(
		.INIT('h00b2)
	) name15227 (
		_w15149_,
		_w15178_,
		_w15185_,
		_w15259_,
		_w15261_
	);
	LUT4 #(
		.INIT('h4d00)
	) name15228 (
		_w15149_,
		_w15178_,
		_w15185_,
		_w15259_,
		_w15262_
	);
	LUT4 #(
		.INIT('hb24d)
	) name15229 (
		_w15149_,
		_w15178_,
		_w15185_,
		_w15259_,
		_w15263_
	);
	LUT4 #(
		.INIT('h2228)
	) name15230 (
		_w3214_,
		_w7695_,
		_w7750_,
		_w11285_,
		_w15264_
	);
	LUT4 #(
		.INIT('h007d)
	) name15231 (
		_w3249_,
		_w11286_,
		_w11335_,
		_w15264_,
		_w15265_
	);
	LUT3 #(
		.INIT('h70)
	) name15232 (
		_w3262_,
		_w11377_,
		_w15265_,
		_w15266_
	);
	LUT4 #(
		.INIT('h95aa)
	) name15233 (
		\a[23] ,
		_w37_,
		_w12799_,
		_w15266_,
		_w15267_
	);
	LUT2 #(
		.INIT('h9)
	) name15234 (
		_w15263_,
		_w15267_,
		_w15268_
	);
	LUT3 #(
		.INIT('h4d)
	) name15235 (
		_w15148_,
		_w15186_,
		_w15193_,
		_w15269_
	);
	LUT4 #(
		.INIT('h2228)
	) name15236 (
		_w3311_,
		_w11549_,
		_w11373_,
		_w11375_,
		_w15270_
	);
	LUT4 #(
		.INIT('h007d)
	) name15237 (
		_w3645_,
		_w13062_,
		_w13099_,
		_w15270_,
		_w15271_
	);
	LUT3 #(
		.INIT('h70)
	) name15238 (
		_w3654_,
		_w13247_,
		_w15271_,
		_w15272_
	);
	LUT4 #(
		.INIT('h95aa)
	) name15239 (
		\a[20] ,
		_w3312_,
		_w13576_,
		_w15272_,
		_w15273_
	);
	LUT3 #(
		.INIT('h69)
	) name15240 (
		_w15268_,
		_w15269_,
		_w15273_,
		_w15274_
	);
	LUT3 #(
		.INIT('h4d)
	) name15241 (
		_w15147_,
		_w15194_,
		_w15201_,
		_w15275_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15242 (
		_w3709_,
		_w13243_,
		_w13245_,
		_w13285_,
		_w15276_
	);
	LUT4 #(
		.INIT('h007d)
	) name15243 (
		_w3877_,
		_w13293_,
		_w13322_,
		_w15276_,
		_w15277_
	);
	LUT3 #(
		.INIT('h70)
	) name15244 (
		_w3886_,
		_w13716_,
		_w15277_,
		_w15278_
	);
	LUT4 #(
		.INIT('h95aa)
	) name15245 (
		\a[17] ,
		_w3710_,
		_w13720_,
		_w15278_,
		_w15279_
	);
	LUT3 #(
		.INIT('h69)
	) name15246 (
		_w15274_,
		_w15275_,
		_w15279_,
		_w15280_
	);
	LUT3 #(
		.INIT('h4d)
	) name15247 (
		_w15146_,
		_w15202_,
		_w15209_,
		_w15281_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15248 (
		_w4033_,
		_w13712_,
		_w13714_,
		_w13847_,
		_w15282_
	);
	LUT4 #(
		.INIT('h007d)
	) name15249 (
		_w4367_,
		_w13960_,
		_w13979_,
		_w15282_,
		_w15283_
	);
	LUT3 #(
		.INIT('h70)
	) name15250 (
		_w4382_,
		_w14112_,
		_w15283_,
		_w15284_
	);
	LUT4 #(
		.INIT('h95aa)
	) name15251 (
		\a[14] ,
		_w4034_,
		_w14116_,
		_w15284_,
		_w15285_
	);
	LUT3 #(
		.INIT('h69)
	) name15252 (
		_w15280_,
		_w15281_,
		_w15285_,
		_w15286_
	);
	LUT2 #(
		.INIT('h6)
	) name15253 (
		_w15232_,
		_w15286_,
		_w15287_
	);
	LUT3 #(
		.INIT('h4d)
	) name15254 (
		_w15137_,
		_w15211_,
		_w15218_,
		_w15288_
	);
	LUT2 #(
		.INIT('h8)
	) name15255 (
		_w15287_,
		_w15288_,
		_w15289_
	);
	LUT2 #(
		.INIT('h6)
	) name15256 (
		_w15287_,
		_w15288_,
		_w15290_
	);
	LUT3 #(
		.INIT('h1e)
	) name15257 (
		_w15220_,
		_w15222_,
		_w15290_,
		_w15291_
	);
	LUT2 #(
		.INIT('h6)
	) name15258 (
		_w15224_,
		_w15291_,
		_w15292_
	);
	LUT4 #(
		.INIT('h010f)
	) name15259 (
		_w15220_,
		_w15222_,
		_w15289_,
		_w15290_,
		_w15293_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15260 (
		_w2875_,
		_w11384_,
		_w11488_,
		_w11489_,
		_w15294_
	);
	LUT4 #(
		.INIT('h2228)
	) name15261 (
		_w2986_,
		_w7695_,
		_w7750_,
		_w11285_,
		_w15295_
	);
	LUT3 #(
		.INIT('h82)
	) name15262 (
		_w2874_,
		_w11280_,
		_w11282_,
		_w15296_
	);
	LUT3 #(
		.INIT('h07)
	) name15263 (
		_w2975_,
		_w11382_,
		_w15296_,
		_w15297_
	);
	LUT2 #(
		.INIT('h4)
	) name15264 (
		_w15295_,
		_w15297_,
		_w15298_
	);
	LUT3 #(
		.INIT('h9a)
	) name15265 (
		\a[26] ,
		_w15294_,
		_w15298_,
		_w15299_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15266 (
		_w2550_,
		_w11390_,
		_w11482_,
		_w11483_,
		_w15300_
	);
	LUT4 #(
		.INIT('h2228)
	) name15267 (
		_w2854_,
		_w7935_,
		_w8077_,
		_w11279_,
		_w15301_
	);
	LUT3 #(
		.INIT('h82)
	) name15268 (
		_w2549_,
		_w11274_,
		_w11276_,
		_w15302_
	);
	LUT3 #(
		.INIT('h07)
	) name15269 (
		_w2617_,
		_w11388_,
		_w15302_,
		_w15303_
	);
	LUT2 #(
		.INIT('h4)
	) name15270 (
		_w15301_,
		_w15303_,
		_w15304_
	);
	LUT3 #(
		.INIT('h9a)
	) name15271 (
		\a[29] ,
		_w15300_,
		_w15304_,
		_w15305_
	);
	LUT3 #(
		.INIT('hb2)
	) name15272 (
		_w15237_,
		_w15246_,
		_w15250_,
		_w15306_
	);
	LUT4 #(
		.INIT('hb332)
	) name15273 (
		_w15150_,
		_w15157_,
		_w15165_,
		_w15245_,
		_w15307_
	);
	LUT4 #(
		.INIT('h5665)
	) name15274 (
		\a[11] ,
		_w7545_,
		_w14344_,
		_w14347_,
		_w15308_
	);
	LUT4 #(
		.INIT('h0777)
	) name15275 (
		_w106_,
		_w55_,
		_w52_,
		_w236_,
		_w15309_
	);
	LUT4 #(
		.INIT('h8000)
	) name15276 (
		_w408_,
		_w522_,
		_w803_,
		_w15309_,
		_w15310_
	);
	LUT4 #(
		.INIT('h4000)
	) name15277 (
		_w457_,
		_w974_,
		_w1401_,
		_w3433_,
		_w15311_
	);
	LUT2 #(
		.INIT('h8)
	) name15278 (
		_w15310_,
		_w15311_,
		_w15312_
	);
	LUT3 #(
		.INIT('h80)
	) name15279 (
		_w1068_,
		_w2160_,
		_w2258_,
		_w15313_
	);
	LUT3 #(
		.INIT('h80)
	) name15280 (
		_w1941_,
		_w3443_,
		_w15313_,
		_w15314_
	);
	LUT3 #(
		.INIT('h80)
	) name15281 (
		_w1488_,
		_w15312_,
		_w15314_,
		_w15315_
	);
	LUT4 #(
		.INIT('h8000)
	) name15282 (
		_w779_,
		_w792_,
		_w1508_,
		_w1517_,
		_w15316_
	);
	LUT2 #(
		.INIT('h8)
	) name15283 (
		_w15315_,
		_w15316_,
		_w15317_
	);
	LUT4 #(
		.INIT('h8000)
	) name15284 (
		_w1692_,
		_w15156_,
		_w15315_,
		_w15316_,
		_w15318_
	);
	LUT4 #(
		.INIT('h0777)
	) name15285 (
		_w1692_,
		_w15156_,
		_w15315_,
		_w15316_,
		_w15319_
	);
	LUT4 #(
		.INIT('h7888)
	) name15286 (
		_w1692_,
		_w15156_,
		_w15315_,
		_w15316_,
		_w15320_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15287 (
		_w377_,
		_w11396_,
		_w11476_,
		_w11477_,
		_w15321_
	);
	LUT4 #(
		.INIT('h2228)
	) name15288 (
		_w2527_,
		_w8466_,
		_w8541_,
		_w11273_,
		_w15322_
	);
	LUT3 #(
		.INIT('h82)
	) name15289 (
		_w376_,
		_w11268_,
		_w11270_,
		_w15323_
	);
	LUT3 #(
		.INIT('h07)
	) name15290 (
		_w2407_,
		_w11394_,
		_w15323_,
		_w15324_
	);
	LUT2 #(
		.INIT('h4)
	) name15291 (
		_w15322_,
		_w15324_,
		_w15325_
	);
	LUT2 #(
		.INIT('h4)
	) name15292 (
		_w15321_,
		_w15325_,
		_w15326_
	);
	LUT3 #(
		.INIT('h06)
	) name15293 (
		_w15308_,
		_w15320_,
		_w15326_,
		_w15327_
	);
	LUT3 #(
		.INIT('h90)
	) name15294 (
		_w15308_,
		_w15320_,
		_w15326_,
		_w15328_
	);
	LUT3 #(
		.INIT('h69)
	) name15295 (
		_w15308_,
		_w15320_,
		_w15326_,
		_w15329_
	);
	LUT2 #(
		.INIT('h9)
	) name15296 (
		_w15307_,
		_w15329_,
		_w15330_
	);
	LUT4 #(
		.INIT('h4114)
	) name15297 (
		_w15299_,
		_w15305_,
		_w15306_,
		_w15330_,
		_w15331_
	);
	LUT4 #(
		.INIT('h9669)
	) name15298 (
		_w15299_,
		_w15305_,
		_w15306_,
		_w15330_,
		_w15332_
	);
	LUT4 #(
		.INIT('h4d00)
	) name15299 (
		_w15233_,
		_w15251_,
		_w15258_,
		_w15332_,
		_w15333_
	);
	LUT4 #(
		.INIT('hdc23)
	) name15300 (
		_w15252_,
		_w15253_,
		_w15258_,
		_w15332_,
		_w15334_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15301 (
		_w37_,
		_w11378_,
		_w11494_,
		_w11552_,
		_w15335_
	);
	LUT4 #(
		.INIT('h2228)
	) name15302 (
		_w3262_,
		_w11549_,
		_w11373_,
		_w11375_,
		_w15336_
	);
	LUT3 #(
		.INIT('h82)
	) name15303 (
		_w3214_,
		_w11286_,
		_w11335_,
		_w15337_
	);
	LUT3 #(
		.INIT('h07)
	) name15304 (
		_w3249_,
		_w11377_,
		_w15337_,
		_w15338_
	);
	LUT2 #(
		.INIT('h4)
	) name15305 (
		_w15336_,
		_w15338_,
		_w15339_
	);
	LUT3 #(
		.INIT('h9a)
	) name15306 (
		\a[23] ,
		_w15335_,
		_w15339_,
		_w15340_
	);
	LUT2 #(
		.INIT('h2)
	) name15307 (
		_w15334_,
		_w15340_,
		_w15341_
	);
	LUT2 #(
		.INIT('h9)
	) name15308 (
		_w15334_,
		_w15340_,
		_w15342_
	);
	LUT4 #(
		.INIT('h8e00)
	) name15309 (
		_w15259_,
		_w15260_,
		_w15267_,
		_w15342_,
		_w15343_
	);
	LUT4 #(
		.INIT('hba45)
	) name15310 (
		_w15261_,
		_w15262_,
		_w15267_,
		_w15342_,
		_w15344_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15311 (
		_w3312_,
		_w13288_,
		_w13290_,
		_w13291_,
		_w15345_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15312 (
		_w3654_,
		_w13243_,
		_w13245_,
		_w13285_,
		_w15346_
	);
	LUT3 #(
		.INIT('h82)
	) name15313 (
		_w3311_,
		_w13062_,
		_w13099_,
		_w15347_
	);
	LUT3 #(
		.INIT('h07)
	) name15314 (
		_w3645_,
		_w13247_,
		_w15347_,
		_w15348_
	);
	LUT2 #(
		.INIT('h4)
	) name15315 (
		_w15346_,
		_w15348_,
		_w15349_
	);
	LUT3 #(
		.INIT('h9a)
	) name15316 (
		\a[20] ,
		_w15345_,
		_w15349_,
		_w15350_
	);
	LUT3 #(
		.INIT('h8e)
	) name15317 (
		_w15268_,
		_w15269_,
		_w15273_,
		_w15351_
	);
	LUT4 #(
		.INIT('h008e)
	) name15318 (
		_w15268_,
		_w15269_,
		_w15273_,
		_w15350_,
		_w15352_
	);
	LUT4 #(
		.INIT('h7100)
	) name15319 (
		_w15268_,
		_w15269_,
		_w15273_,
		_w15350_,
		_w15353_
	);
	LUT4 #(
		.INIT('h8e71)
	) name15320 (
		_w15268_,
		_w15269_,
		_w15273_,
		_w15350_,
		_w15354_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15321 (
		_w3710_,
		_w13717_,
		_w13719_,
		_w13850_,
		_w15355_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15322 (
		_w3886_,
		_w13712_,
		_w13714_,
		_w13847_,
		_w15356_
	);
	LUT3 #(
		.INIT('h82)
	) name15323 (
		_w3709_,
		_w13293_,
		_w13322_,
		_w15357_
	);
	LUT3 #(
		.INIT('h07)
	) name15324 (
		_w3877_,
		_w13716_,
		_w15357_,
		_w15358_
	);
	LUT2 #(
		.INIT('h4)
	) name15325 (
		_w15356_,
		_w15358_,
		_w15359_
	);
	LUT3 #(
		.INIT('h9a)
	) name15326 (
		\a[17] ,
		_w15355_,
		_w15359_,
		_w15360_
	);
	LUT3 #(
		.INIT('h06)
	) name15327 (
		_w15344_,
		_w15354_,
		_w15360_,
		_w15361_
	);
	LUT3 #(
		.INIT('h90)
	) name15328 (
		_w15344_,
		_w15354_,
		_w15360_,
		_w15362_
	);
	LUT3 #(
		.INIT('h69)
	) name15329 (
		_w15344_,
		_w15354_,
		_w15360_,
		_w15363_
	);
	LUT3 #(
		.INIT('h8e)
	) name15330 (
		_w15274_,
		_w15275_,
		_w15279_,
		_w15364_
	);
	LUT2 #(
		.INIT('h6)
	) name15331 (
		_w15363_,
		_w15364_,
		_w15365_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15332 (
		_w4034_,
		_w14113_,
		_w14115_,
		_w14238_,
		_w15366_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15333 (
		_w4382_,
		_w14108_,
		_w14111_,
		_w14235_,
		_w15367_
	);
	LUT3 #(
		.INIT('h82)
	) name15334 (
		_w4033_,
		_w13960_,
		_w13979_,
		_w15368_
	);
	LUT3 #(
		.INIT('h07)
	) name15335 (
		_w4367_,
		_w14112_,
		_w15368_,
		_w15369_
	);
	LUT2 #(
		.INIT('h4)
	) name15336 (
		_w15367_,
		_w15369_,
		_w15370_
	);
	LUT3 #(
		.INIT('h9a)
	) name15337 (
		\a[14] ,
		_w15366_,
		_w15370_,
		_w15371_
	);
	LUT4 #(
		.INIT('h008e)
	) name15338 (
		_w15280_,
		_w15281_,
		_w15285_,
		_w15371_,
		_w15372_
	);
	LUT4 #(
		.INIT('h7100)
	) name15339 (
		_w15280_,
		_w15281_,
		_w15285_,
		_w15371_,
		_w15373_
	);
	LUT4 #(
		.INIT('h8e71)
	) name15340 (
		_w15280_,
		_w15281_,
		_w15285_,
		_w15371_,
		_w15374_
	);
	LUT2 #(
		.INIT('h6)
	) name15341 (
		_w15365_,
		_w15374_,
		_w15375_
	);
	LUT3 #(
		.INIT('h32)
	) name15342 (
		_w15230_,
		_w15231_,
		_w15286_,
		_w15376_
	);
	LUT2 #(
		.INIT('h8)
	) name15343 (
		_w15375_,
		_w15376_,
		_w15377_
	);
	LUT2 #(
		.INIT('h1)
	) name15344 (
		_w15375_,
		_w15376_,
		_w15378_
	);
	LUT2 #(
		.INIT('h6)
	) name15345 (
		_w15375_,
		_w15376_,
		_w15379_
	);
	LUT4 #(
		.INIT('h8008)
	) name15346 (
		_w15224_,
		_w15291_,
		_w15293_,
		_w15379_,
		_w15380_
	);
	LUT4 #(
		.INIT('h7887)
	) name15347 (
		_w15224_,
		_w15291_,
		_w15293_,
		_w15379_,
		_w15381_
	);
	LUT3 #(
		.INIT('h31)
	) name15348 (
		_w15365_,
		_w15372_,
		_w15373_,
		_w15382_
	);
	LUT3 #(
		.INIT('h45)
	) name15349 (
		_w15361_,
		_w15362_,
		_w15364_,
		_w15383_
	);
	LUT3 #(
		.INIT('h82)
	) name15350 (
		_w3710_,
		_w13959_,
		_w13982_,
		_w15384_
	);
	LUT3 #(
		.INIT('h82)
	) name15351 (
		_w3886_,
		_w13960_,
		_w13979_,
		_w15385_
	);
	LUT2 #(
		.INIT('h8)
	) name15352 (
		_w3709_,
		_w13716_,
		_w15386_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15353 (
		_w3877_,
		_w13712_,
		_w13714_,
		_w13847_,
		_w15387_
	);
	LUT2 #(
		.INIT('h1)
	) name15354 (
		_w15386_,
		_w15387_,
		_w15388_
	);
	LUT2 #(
		.INIT('h4)
	) name15355 (
		_w15385_,
		_w15388_,
		_w15389_
	);
	LUT3 #(
		.INIT('h9a)
	) name15356 (
		\a[17] ,
		_w15384_,
		_w15389_,
		_w15390_
	);
	LUT3 #(
		.INIT('h31)
	) name15357 (
		_w15344_,
		_w15352_,
		_w15353_,
		_w15391_
	);
	LUT3 #(
		.INIT('h32)
	) name15358 (
		_w15307_,
		_w15327_,
		_w15328_,
		_w15392_
	);
	LUT3 #(
		.INIT('h0d)
	) name15359 (
		_w15308_,
		_w15318_,
		_w15319_,
		_w15393_
	);
	LUT4 #(
		.INIT('h1000)
	) name15360 (
		_w451_,
		_w476_,
		_w479_,
		_w1181_,
		_w15394_
	);
	LUT4 #(
		.INIT('h4000)
	) name15361 (
		_w335_,
		_w861_,
		_w1514_,
		_w1564_,
		_w15395_
	);
	LUT3 #(
		.INIT('h80)
	) name15362 (
		_w1905_,
		_w2067_,
		_w2369_,
		_w15396_
	);
	LUT4 #(
		.INIT('h8000)
	) name15363 (
		_w7264_,
		_w15396_,
		_w15394_,
		_w15395_,
		_w15397_
	);
	LUT3 #(
		.INIT('h80)
	) name15364 (
		_w14155_,
		_w14400_,
		_w15397_,
		_w15398_
	);
	LUT4 #(
		.INIT('h8000)
	) name15365 (
		_w11304_,
		_w11307_,
		_w7986_,
		_w7989_,
		_w15399_
	);
	LUT2 #(
		.INIT('h8)
	) name15366 (
		_w15398_,
		_w15399_,
		_w15400_
	);
	LUT4 #(
		.INIT('h4d00)
	) name15367 (
		_w15157_,
		_w15308_,
		_w15317_,
		_w15400_,
		_w15401_
	);
	LUT4 #(
		.INIT('h00b2)
	) name15368 (
		_w15157_,
		_w15308_,
		_w15317_,
		_w15400_,
		_w15402_
	);
	LUT4 #(
		.INIT('h0df2)
	) name15369 (
		_w15308_,
		_w15318_,
		_w15319_,
		_w15400_,
		_w15403_
	);
	LUT3 #(
		.INIT('h82)
	) name15370 (
		_w377_,
		_w11478_,
		_w11480_,
		_w15404_
	);
	LUT3 #(
		.INIT('h82)
	) name15371 (
		_w2527_,
		_w11274_,
		_w11276_,
		_w15405_
	);
	LUT2 #(
		.INIT('h8)
	) name15372 (
		_w376_,
		_w11394_,
		_w15406_
	);
	LUT4 #(
		.INIT('h2228)
	) name15373 (
		_w2407_,
		_w8466_,
		_w8541_,
		_w11273_,
		_w15407_
	);
	LUT2 #(
		.INIT('h1)
	) name15374 (
		_w15406_,
		_w15407_,
		_w15408_
	);
	LUT2 #(
		.INIT('h4)
	) name15375 (
		_w15405_,
		_w15408_,
		_w15409_
	);
	LUT2 #(
		.INIT('h4)
	) name15376 (
		_w15404_,
		_w15409_,
		_w15410_
	);
	LUT2 #(
		.INIT('h9)
	) name15377 (
		_w15403_,
		_w15410_,
		_w15411_
	);
	LUT4 #(
		.INIT('h0023)
	) name15378 (
		_w15307_,
		_w15327_,
		_w15329_,
		_w15411_,
		_w15412_
	);
	LUT4 #(
		.INIT('hdc00)
	) name15379 (
		_w15307_,
		_w15327_,
		_w15329_,
		_w15411_,
		_w15413_
	);
	LUT4 #(
		.INIT('h32cd)
	) name15380 (
		_w15307_,
		_w15327_,
		_w15328_,
		_w15411_,
		_w15414_
	);
	LUT3 #(
		.INIT('h82)
	) name15381 (
		_w2550_,
		_w11484_,
		_w11486_,
		_w15415_
	);
	LUT3 #(
		.INIT('h82)
	) name15382 (
		_w2854_,
		_w11280_,
		_w11282_,
		_w15416_
	);
	LUT2 #(
		.INIT('h8)
	) name15383 (
		_w2549_,
		_w11388_,
		_w15417_
	);
	LUT4 #(
		.INIT('h2228)
	) name15384 (
		_w2617_,
		_w7935_,
		_w8077_,
		_w11279_,
		_w15418_
	);
	LUT2 #(
		.INIT('h1)
	) name15385 (
		_w15417_,
		_w15418_,
		_w15419_
	);
	LUT2 #(
		.INIT('h4)
	) name15386 (
		_w15416_,
		_w15419_,
		_w15420_
	);
	LUT3 #(
		.INIT('h9a)
	) name15387 (
		\a[29] ,
		_w15415_,
		_w15420_,
		_w15421_
	);
	LUT2 #(
		.INIT('h9)
	) name15388 (
		_w15414_,
		_w15421_,
		_w15422_
	);
	LUT3 #(
		.INIT('h71)
	) name15389 (
		_w15305_,
		_w15306_,
		_w15330_,
		_w15423_
	);
	LUT3 #(
		.INIT('h82)
	) name15390 (
		_w2875_,
		_w11490_,
		_w11492_,
		_w15424_
	);
	LUT3 #(
		.INIT('h82)
	) name15391 (
		_w2986_,
		_w11286_,
		_w11335_,
		_w15425_
	);
	LUT2 #(
		.INIT('h8)
	) name15392 (
		_w2874_,
		_w11382_,
		_w15426_
	);
	LUT4 #(
		.INIT('h2228)
	) name15393 (
		_w2975_,
		_w7695_,
		_w7750_,
		_w11285_,
		_w15427_
	);
	LUT2 #(
		.INIT('h1)
	) name15394 (
		_w15426_,
		_w15427_,
		_w15428_
	);
	LUT2 #(
		.INIT('h4)
	) name15395 (
		_w15425_,
		_w15428_,
		_w15429_
	);
	LUT3 #(
		.INIT('h9a)
	) name15396 (
		\a[26] ,
		_w15424_,
		_w15429_,
		_w15430_
	);
	LUT3 #(
		.INIT('h69)
	) name15397 (
		_w15422_,
		_w15423_,
		_w15430_,
		_w15431_
	);
	LUT3 #(
		.INIT('h82)
	) name15398 (
		_w37_,
		_w13061_,
		_w13102_,
		_w15432_
	);
	LUT3 #(
		.INIT('h82)
	) name15399 (
		_w3262_,
		_w13062_,
		_w13099_,
		_w15433_
	);
	LUT2 #(
		.INIT('h8)
	) name15400 (
		_w3214_,
		_w11377_,
		_w15434_
	);
	LUT4 #(
		.INIT('h2228)
	) name15401 (
		_w3249_,
		_w11549_,
		_w11373_,
		_w11375_,
		_w15435_
	);
	LUT2 #(
		.INIT('h1)
	) name15402 (
		_w15434_,
		_w15435_,
		_w15436_
	);
	LUT2 #(
		.INIT('h4)
	) name15403 (
		_w15433_,
		_w15436_,
		_w15437_
	);
	LUT3 #(
		.INIT('h9a)
	) name15404 (
		\a[23] ,
		_w15432_,
		_w15437_,
		_w15438_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name15405 (
		_w15331_,
		_w15333_,
		_w15431_,
		_w15438_,
		_w15439_
	);
	LUT3 #(
		.INIT('h82)
	) name15406 (
		_w3312_,
		_w13292_,
		_w13325_,
		_w15440_
	);
	LUT3 #(
		.INIT('h82)
	) name15407 (
		_w3654_,
		_w13293_,
		_w13322_,
		_w15441_
	);
	LUT2 #(
		.INIT('h8)
	) name15408 (
		_w3311_,
		_w13247_,
		_w15442_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15409 (
		_w3645_,
		_w13243_,
		_w13245_,
		_w13285_,
		_w15443_
	);
	LUT2 #(
		.INIT('h1)
	) name15410 (
		_w15442_,
		_w15443_,
		_w15444_
	);
	LUT2 #(
		.INIT('h4)
	) name15411 (
		_w15441_,
		_w15444_,
		_w15445_
	);
	LUT3 #(
		.INIT('h9a)
	) name15412 (
		\a[20] ,
		_w15440_,
		_w15445_,
		_w15446_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name15413 (
		_w15341_,
		_w15343_,
		_w15439_,
		_w15446_,
		_w15447_
	);
	LUT4 #(
		.INIT('hb200)
	) name15414 (
		_w15344_,
		_w15350_,
		_w15351_,
		_w15447_,
		_w15448_
	);
	LUT4 #(
		.INIT('h004d)
	) name15415 (
		_w15344_,
		_w15350_,
		_w15351_,
		_w15447_,
		_w15449_
	);
	LUT4 #(
		.INIT('h31ce)
	) name15416 (
		_w15344_,
		_w15352_,
		_w15353_,
		_w15447_,
		_w15450_
	);
	LUT2 #(
		.INIT('h9)
	) name15417 (
		_w15390_,
		_w15450_,
		_w15451_
	);
	LUT3 #(
		.INIT('h82)
	) name15418 (
		_w4034_,
		_w14343_,
		_w14349_,
		_w15452_
	);
	LUT3 #(
		.INIT('h28)
	) name15419 (
		_w4382_,
		_w14344_,
		_w14347_,
		_w15453_
	);
	LUT2 #(
		.INIT('h8)
	) name15420 (
		_w4033_,
		_w14112_,
		_w15454_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15421 (
		_w4367_,
		_w14108_,
		_w14111_,
		_w14235_,
		_w15455_
	);
	LUT2 #(
		.INIT('h1)
	) name15422 (
		_w15454_,
		_w15455_,
		_w15456_
	);
	LUT2 #(
		.INIT('h4)
	) name15423 (
		_w15453_,
		_w15456_,
		_w15457_
	);
	LUT3 #(
		.INIT('h9a)
	) name15424 (
		\a[14] ,
		_w15452_,
		_w15457_,
		_w15458_
	);
	LUT3 #(
		.INIT('h96)
	) name15425 (
		_w15383_,
		_w15451_,
		_w15458_,
		_w15459_
	);
	LUT2 #(
		.INIT('h4)
	) name15426 (
		_w15382_,
		_w15459_,
		_w15460_
	);
	LUT2 #(
		.INIT('h9)
	) name15427 (
		_w15382_,
		_w15459_,
		_w15461_
	);
	LUT4 #(
		.INIT('hd400)
	) name15428 (
		_w15293_,
		_w15375_,
		_w15376_,
		_w15461_,
		_w15462_
	);
	LUT4 #(
		.INIT('h32cd)
	) name15429 (
		_w15293_,
		_w15377_,
		_w15378_,
		_w15461_,
		_w15463_
	);
	LUT2 #(
		.INIT('h8)
	) name15430 (
		_w15380_,
		_w15463_,
		_w15464_
	);
	LUT2 #(
		.INIT('h6)
	) name15431 (
		_w15380_,
		_w15463_,
		_w15465_
	);
	LUT3 #(
		.INIT('h32)
	) name15432 (
		_w15390_,
		_w15448_,
		_w15449_,
		_w15466_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name15433 (
		_w4034_,
		_w14343_,
		_w14348_,
		_w14349_,
		_w15467_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15434 (
		_w4033_,
		_w14108_,
		_w14111_,
		_w14235_,
		_w15468_
	);
	LUT4 #(
		.INIT('h00eb)
	) name15435 (
		_w8080_,
		_w14344_,
		_w14347_,
		_w15468_,
		_w15469_
	);
	LUT3 #(
		.INIT('h9a)
	) name15436 (
		\a[14] ,
		_w15467_,
		_w15469_,
		_w15470_
	);
	LUT4 #(
		.INIT('h0071)
	) name15437 (
		_w15390_,
		_w15391_,
		_w15447_,
		_w15470_,
		_w15471_
	);
	LUT4 #(
		.INIT('h8e00)
	) name15438 (
		_w15390_,
		_w15391_,
		_w15447_,
		_w15470_,
		_w15472_
	);
	LUT4 #(
		.INIT('hcd32)
	) name15439 (
		_w15390_,
		_w15448_,
		_w15449_,
		_w15470_,
		_w15473_
	);
	LUT4 #(
		.INIT('h2228)
	) name15440 (
		_w2874_,
		_w7695_,
		_w7750_,
		_w11285_,
		_w15474_
	);
	LUT4 #(
		.INIT('h007d)
	) name15441 (
		_w2975_,
		_w11286_,
		_w11335_,
		_w15474_,
		_w15475_
	);
	LUT3 #(
		.INIT('h70)
	) name15442 (
		_w2986_,
		_w11377_,
		_w15475_,
		_w15476_
	);
	LUT4 #(
		.INIT('h95aa)
	) name15443 (
		\a[26] ,
		_w2875_,
		_w12799_,
		_w15476_,
		_w15477_
	);
	LUT4 #(
		.INIT('h8000)
	) name15444 (
		_w628_,
		_w632_,
		_w2371_,
		_w2375_,
		_w15478_
	);
	LUT3 #(
		.INIT('h80)
	) name15445 (
		_w620_,
		_w1099_,
		_w2495_,
		_w15479_
	);
	LUT4 #(
		.INIT('h0777)
	) name15446 (
		_w106_,
		_w59_,
		_w93_,
		_w201_,
		_w15480_
	);
	LUT4 #(
		.INIT('h153f)
	) name15447 (
		_w90_,
		_w46_,
		_w184_,
		_w158_,
		_w15481_
	);
	LUT4 #(
		.INIT('h8000)
	) name15448 (
		_w196_,
		_w442_,
		_w15480_,
		_w15481_,
		_w15482_
	);
	LUT4 #(
		.INIT('h8000)
	) name15449 (
		_w1942_,
		_w2467_,
		_w15479_,
		_w15482_,
		_w15483_
	);
	LUT4 #(
		.INIT('h8000)
	) name15450 (
		_w2110_,
		_w3547_,
		_w15483_,
		_w15478_,
		_w15484_
	);
	LUT4 #(
		.INIT('h40c0)
	) name15451 (
		_w2775_,
		_w15398_,
		_w15399_,
		_w15484_,
		_w15485_
	);
	LUT4 #(
		.INIT('h953f)
	) name15452 (
		_w2775_,
		_w15398_,
		_w15399_,
		_w15484_,
		_w15486_
	);
	LUT4 #(
		.INIT('h2228)
	) name15453 (
		_w376_,
		_w8466_,
		_w8541_,
		_w11273_,
		_w15487_
	);
	LUT4 #(
		.INIT('h007d)
	) name15454 (
		_w2407_,
		_w11274_,
		_w11276_,
		_w15487_,
		_w15488_
	);
	LUT3 #(
		.INIT('h70)
	) name15455 (
		_w2527_,
		_w11388_,
		_w15488_,
		_w15489_
	);
	LUT4 #(
		.INIT('h80f0)
	) name15456 (
		_w377_,
		_w12391_,
		_w15486_,
		_w15489_,
		_w15490_
	);
	LUT4 #(
		.INIT('h780f)
	) name15457 (
		_w377_,
		_w12391_,
		_w15486_,
		_w15489_,
		_w15491_
	);
	LUT4 #(
		.INIT('h4d00)
	) name15458 (
		_w15393_,
		_w15400_,
		_w15410_,
		_w15491_,
		_w15492_
	);
	LUT4 #(
		.INIT('hdc23)
	) name15459 (
		_w15401_,
		_w15402_,
		_w15410_,
		_w15491_,
		_w15493_
	);
	LUT4 #(
		.INIT('h4d00)
	) name15460 (
		_w15392_,
		_w15411_,
		_w15421_,
		_w15493_,
		_w15494_
	);
	LUT4 #(
		.INIT('h32cd)
	) name15461 (
		_w15412_,
		_w15413_,
		_w15421_,
		_w15493_,
		_w15495_
	);
	LUT4 #(
		.INIT('h2228)
	) name15462 (
		_w2549_,
		_w7935_,
		_w8077_,
		_w11279_,
		_w15496_
	);
	LUT4 #(
		.INIT('h007d)
	) name15463 (
		_w2617_,
		_w11280_,
		_w11282_,
		_w15496_,
		_w15497_
	);
	LUT3 #(
		.INIT('h70)
	) name15464 (
		_w2854_,
		_w11382_,
		_w15497_,
		_w15498_
	);
	LUT4 #(
		.INIT('h95aa)
	) name15465 (
		\a[29] ,
		_w2550_,
		_w12476_,
		_w15498_,
		_w15499_
	);
	LUT3 #(
		.INIT('h96)
	) name15466 (
		_w15477_,
		_w15495_,
		_w15499_,
		_w15500_
	);
	LUT3 #(
		.INIT('h8e)
	) name15467 (
		_w15422_,
		_w15423_,
		_w15430_,
		_w15501_
	);
	LUT4 #(
		.INIT('h2228)
	) name15468 (
		_w3214_,
		_w11549_,
		_w11373_,
		_w11375_,
		_w15502_
	);
	LUT4 #(
		.INIT('h007d)
	) name15469 (
		_w3249_,
		_w13062_,
		_w13099_,
		_w15502_,
		_w15503_
	);
	LUT3 #(
		.INIT('h70)
	) name15470 (
		_w3262_,
		_w13247_,
		_w15503_,
		_w15504_
	);
	LUT4 #(
		.INIT('h95aa)
	) name15471 (
		\a[23] ,
		_w37_,
		_w13576_,
		_w15504_,
		_w15505_
	);
	LUT3 #(
		.INIT('h69)
	) name15472 (
		_w15500_,
		_w15501_,
		_w15505_,
		_w15506_
	);
	LUT4 #(
		.INIT('he0fe)
	) name15473 (
		_w15331_,
		_w15333_,
		_w15431_,
		_w15438_,
		_w15507_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15474 (
		_w3311_,
		_w13243_,
		_w13245_,
		_w13285_,
		_w15508_
	);
	LUT4 #(
		.INIT('h007d)
	) name15475 (
		_w3645_,
		_w13293_,
		_w13322_,
		_w15508_,
		_w15509_
	);
	LUT3 #(
		.INIT('h70)
	) name15476 (
		_w3654_,
		_w13716_,
		_w15509_,
		_w15510_
	);
	LUT4 #(
		.INIT('h95aa)
	) name15477 (
		\a[20] ,
		_w3312_,
		_w13720_,
		_w15510_,
		_w15511_
	);
	LUT3 #(
		.INIT('h69)
	) name15478 (
		_w15506_,
		_w15507_,
		_w15511_,
		_w15512_
	);
	LUT4 #(
		.INIT('he0fe)
	) name15479 (
		_w15341_,
		_w15343_,
		_w15439_,
		_w15446_,
		_w15513_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15480 (
		_w3709_,
		_w13712_,
		_w13714_,
		_w13847_,
		_w15514_
	);
	LUT4 #(
		.INIT('h007d)
	) name15481 (
		_w3877_,
		_w13960_,
		_w13979_,
		_w15514_,
		_w15515_
	);
	LUT3 #(
		.INIT('h70)
	) name15482 (
		_w3886_,
		_w14112_,
		_w15515_,
		_w15516_
	);
	LUT4 #(
		.INIT('h95aa)
	) name15483 (
		\a[17] ,
		_w3710_,
		_w14116_,
		_w15516_,
		_w15517_
	);
	LUT3 #(
		.INIT('h69)
	) name15484 (
		_w15512_,
		_w15513_,
		_w15517_,
		_w15518_
	);
	LUT2 #(
		.INIT('h6)
	) name15485 (
		_w15473_,
		_w15518_,
		_w15519_
	);
	LUT3 #(
		.INIT('h4d)
	) name15486 (
		_w15383_,
		_w15451_,
		_w15458_,
		_w15520_
	);
	LUT2 #(
		.INIT('h1)
	) name15487 (
		_w15519_,
		_w15520_,
		_w15521_
	);
	LUT2 #(
		.INIT('h8)
	) name15488 (
		_w15519_,
		_w15520_,
		_w15522_
	);
	LUT2 #(
		.INIT('h6)
	) name15489 (
		_w15519_,
		_w15520_,
		_w15523_
	);
	LUT3 #(
		.INIT('h1e)
	) name15490 (
		_w15460_,
		_w15462_,
		_w15523_,
		_w15524_
	);
	LUT2 #(
		.INIT('h6)
	) name15491 (
		_w15464_,
		_w15524_,
		_w15525_
	);
	LUT4 #(
		.INIT('h00f1)
	) name15492 (
		_w15460_,
		_w15462_,
		_w15521_,
		_w15522_,
		_w15526_
	);
	LUT3 #(
		.INIT('hb2)
	) name15493 (
		_w15477_,
		_w15495_,
		_w15499_,
		_w15527_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15494 (
		_w2550_,
		_w11384_,
		_w11488_,
		_w11489_,
		_w15528_
	);
	LUT4 #(
		.INIT('h2228)
	) name15495 (
		_w2854_,
		_w7695_,
		_w7750_,
		_w11285_,
		_w15529_
	);
	LUT3 #(
		.INIT('h82)
	) name15496 (
		_w2549_,
		_w11280_,
		_w11282_,
		_w15530_
	);
	LUT3 #(
		.INIT('h07)
	) name15497 (
		_w2617_,
		_w11382_,
		_w15530_,
		_w15531_
	);
	LUT2 #(
		.INIT('h4)
	) name15498 (
		_w15529_,
		_w15531_,
		_w15532_
	);
	LUT3 #(
		.INIT('h9a)
	) name15499 (
		\a[29] ,
		_w15528_,
		_w15532_,
		_w15533_
	);
	LUT2 #(
		.INIT('h1)
	) name15500 (
		_w15485_,
		_w15490_,
		_w15534_
	);
	LUT4 #(
		.INIT('h5665)
	) name15501 (
		\a[14] ,
		_w7346_,
		_w14344_,
		_w14347_,
		_w15535_
	);
	LUT4 #(
		.INIT('h2000)
	) name15502 (
		_w172_,
		_w392_,
		_w2143_,
		_w2749_,
		_w15536_
	);
	LUT4 #(
		.INIT('h153f)
	) name15503 (
		_w38_,
		_w122_,
		_w41_,
		_w419_,
		_w15537_
	);
	LUT4 #(
		.INIT('h4000)
	) name15504 (
		_w468_,
		_w882_,
		_w900_,
		_w15537_,
		_w15538_
	);
	LUT4 #(
		.INIT('h8000)
	) name15505 (
		_w7569_,
		_w7834_,
		_w15538_,
		_w15536_,
		_w15539_
	);
	LUT4 #(
		.INIT('h8000)
	) name15506 (
		_w1286_,
		_w1289_,
		_w4275_,
		_w4278_,
		_w15540_
	);
	LUT4 #(
		.INIT('h8000)
	) name15507 (
		_w7436_,
		_w7442_,
		_w15539_,
		_w15540_,
		_w15541_
	);
	LUT4 #(
		.INIT('h8000)
	) name15508 (
		_w1426_,
		_w15398_,
		_w15399_,
		_w15541_,
		_w15542_
	);
	LUT4 #(
		.INIT('h153f)
	) name15509 (
		_w1426_,
		_w15398_,
		_w15399_,
		_w15541_,
		_w15543_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name15510 (
		_w1426_,
		_w15398_,
		_w15399_,
		_w15541_,
		_w15544_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15511 (
		_w377_,
		_w11390_,
		_w11482_,
		_w11483_,
		_w15545_
	);
	LUT4 #(
		.INIT('h2228)
	) name15512 (
		_w2527_,
		_w7935_,
		_w8077_,
		_w11279_,
		_w15546_
	);
	LUT3 #(
		.INIT('h82)
	) name15513 (
		_w376_,
		_w11274_,
		_w11276_,
		_w15547_
	);
	LUT3 #(
		.INIT('h07)
	) name15514 (
		_w2407_,
		_w11388_,
		_w15547_,
		_w15548_
	);
	LUT2 #(
		.INIT('h4)
	) name15515 (
		_w15546_,
		_w15548_,
		_w15549_
	);
	LUT2 #(
		.INIT('h4)
	) name15516 (
		_w15545_,
		_w15549_,
		_w15550_
	);
	LUT4 #(
		.INIT('h6996)
	) name15517 (
		_w15534_,
		_w15535_,
		_w15544_,
		_w15550_,
		_w15551_
	);
	LUT2 #(
		.INIT('h4)
	) name15518 (
		_w15533_,
		_w15551_,
		_w15552_
	);
	LUT2 #(
		.INIT('h2)
	) name15519 (
		_w15533_,
		_w15551_,
		_w15553_
	);
	LUT2 #(
		.INIT('h9)
	) name15520 (
		_w15533_,
		_w15551_,
		_w15554_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15521 (
		_w2875_,
		_w11378_,
		_w11494_,
		_w11552_,
		_w15555_
	);
	LUT4 #(
		.INIT('h2228)
	) name15522 (
		_w2986_,
		_w11549_,
		_w11373_,
		_w11375_,
		_w15556_
	);
	LUT3 #(
		.INIT('h82)
	) name15523 (
		_w2874_,
		_w11286_,
		_w11335_,
		_w15557_
	);
	LUT3 #(
		.INIT('h07)
	) name15524 (
		_w2975_,
		_w11377_,
		_w15557_,
		_w15558_
	);
	LUT2 #(
		.INIT('h4)
	) name15525 (
		_w15556_,
		_w15558_,
		_w15559_
	);
	LUT3 #(
		.INIT('h9a)
	) name15526 (
		\a[26] ,
		_w15555_,
		_w15559_,
		_w15560_
	);
	LUT4 #(
		.INIT('h001e)
	) name15527 (
		_w15492_,
		_w15494_,
		_w15554_,
		_w15560_,
		_w15561_
	);
	LUT4 #(
		.INIT('he100)
	) name15528 (
		_w15492_,
		_w15494_,
		_w15554_,
		_w15560_,
		_w15562_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name15529 (
		_w15492_,
		_w15494_,
		_w15554_,
		_w15560_,
		_w15563_
	);
	LUT2 #(
		.INIT('h9)
	) name15530 (
		_w15527_,
		_w15563_,
		_w15564_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15531 (
		_w37_,
		_w13288_,
		_w13290_,
		_w13291_,
		_w15565_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15532 (
		_w3262_,
		_w13243_,
		_w13245_,
		_w13285_,
		_w15566_
	);
	LUT3 #(
		.INIT('h82)
	) name15533 (
		_w3214_,
		_w13062_,
		_w13099_,
		_w15567_
	);
	LUT3 #(
		.INIT('h07)
	) name15534 (
		_w3249_,
		_w13247_,
		_w15567_,
		_w15568_
	);
	LUT2 #(
		.INIT('h4)
	) name15535 (
		_w15566_,
		_w15568_,
		_w15569_
	);
	LUT3 #(
		.INIT('h9a)
	) name15536 (
		\a[23] ,
		_w15565_,
		_w15569_,
		_w15570_
	);
	LUT4 #(
		.INIT('h008e)
	) name15537 (
		_w15500_,
		_w15501_,
		_w15505_,
		_w15570_,
		_w15571_
	);
	LUT4 #(
		.INIT('h7100)
	) name15538 (
		_w15500_,
		_w15501_,
		_w15505_,
		_w15570_,
		_w15572_
	);
	LUT4 #(
		.INIT('h8e71)
	) name15539 (
		_w15500_,
		_w15501_,
		_w15505_,
		_w15570_,
		_w15573_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15540 (
		_w3312_,
		_w13717_,
		_w13719_,
		_w13850_,
		_w15574_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15541 (
		_w3654_,
		_w13712_,
		_w13714_,
		_w13847_,
		_w15575_
	);
	LUT3 #(
		.INIT('h82)
	) name15542 (
		_w3311_,
		_w13293_,
		_w13322_,
		_w15576_
	);
	LUT3 #(
		.INIT('h07)
	) name15543 (
		_w3645_,
		_w13716_,
		_w15576_,
		_w15577_
	);
	LUT2 #(
		.INIT('h4)
	) name15544 (
		_w15575_,
		_w15577_,
		_w15578_
	);
	LUT3 #(
		.INIT('h9a)
	) name15545 (
		\a[20] ,
		_w15574_,
		_w15578_,
		_w15579_
	);
	LUT3 #(
		.INIT('h06)
	) name15546 (
		_w15564_,
		_w15573_,
		_w15579_,
		_w15580_
	);
	LUT3 #(
		.INIT('h90)
	) name15547 (
		_w15564_,
		_w15573_,
		_w15579_,
		_w15581_
	);
	LUT3 #(
		.INIT('h69)
	) name15548 (
		_w15564_,
		_w15573_,
		_w15579_,
		_w15582_
	);
	LUT3 #(
		.INIT('h8e)
	) name15549 (
		_w15506_,
		_w15507_,
		_w15511_,
		_w15583_
	);
	LUT2 #(
		.INIT('h6)
	) name15550 (
		_w15582_,
		_w15583_,
		_w15584_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15551 (
		_w3710_,
		_w14113_,
		_w14115_,
		_w14238_,
		_w15585_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15552 (
		_w3886_,
		_w14108_,
		_w14111_,
		_w14235_,
		_w15586_
	);
	LUT3 #(
		.INIT('h82)
	) name15553 (
		_w3709_,
		_w13960_,
		_w13979_,
		_w15587_
	);
	LUT3 #(
		.INIT('h07)
	) name15554 (
		_w3877_,
		_w14112_,
		_w15587_,
		_w15588_
	);
	LUT2 #(
		.INIT('h4)
	) name15555 (
		_w15586_,
		_w15588_,
		_w15589_
	);
	LUT3 #(
		.INIT('h9a)
	) name15556 (
		\a[17] ,
		_w15585_,
		_w15589_,
		_w15590_
	);
	LUT3 #(
		.INIT('h8e)
	) name15557 (
		_w15512_,
		_w15513_,
		_w15517_,
		_w15591_
	);
	LUT4 #(
		.INIT('h008e)
	) name15558 (
		_w15512_,
		_w15513_,
		_w15517_,
		_w15590_,
		_w15592_
	);
	LUT4 #(
		.INIT('h7100)
	) name15559 (
		_w15512_,
		_w15513_,
		_w15517_,
		_w15590_,
		_w15593_
	);
	LUT4 #(
		.INIT('h8e71)
	) name15560 (
		_w15512_,
		_w15513_,
		_w15517_,
		_w15590_,
		_w15594_
	);
	LUT2 #(
		.INIT('h6)
	) name15561 (
		_w15584_,
		_w15594_,
		_w15595_
	);
	LUT3 #(
		.INIT('h32)
	) name15562 (
		_w15471_,
		_w15472_,
		_w15518_,
		_w15596_
	);
	LUT4 #(
		.INIT('h7100)
	) name15563 (
		_w15466_,
		_w15470_,
		_w15518_,
		_w15595_,
		_w15597_
	);
	LUT4 #(
		.INIT('h008e)
	) name15564 (
		_w15466_,
		_w15470_,
		_w15518_,
		_w15595_,
		_w15598_
	);
	LUT4 #(
		.INIT('hcd32)
	) name15565 (
		_w15471_,
		_w15472_,
		_w15518_,
		_w15595_,
		_w15599_
	);
	LUT4 #(
		.INIT('h8008)
	) name15566 (
		_w15464_,
		_w15524_,
		_w15526_,
		_w15599_,
		_w15600_
	);
	LUT4 #(
		.INIT('h7887)
	) name15567 (
		_w15464_,
		_w15524_,
		_w15526_,
		_w15599_,
		_w15601_
	);
	LUT3 #(
		.INIT('h45)
	) name15568 (
		_w15580_,
		_w15581_,
		_w15583_,
		_w15602_
	);
	LUT3 #(
		.INIT('h82)
	) name15569 (
		_w3312_,
		_w13959_,
		_w13982_,
		_w15603_
	);
	LUT3 #(
		.INIT('h82)
	) name15570 (
		_w3654_,
		_w13960_,
		_w13979_,
		_w15604_
	);
	LUT2 #(
		.INIT('h8)
	) name15571 (
		_w3311_,
		_w13716_,
		_w15605_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15572 (
		_w3645_,
		_w13712_,
		_w13714_,
		_w13847_,
		_w15606_
	);
	LUT2 #(
		.INIT('h1)
	) name15573 (
		_w15605_,
		_w15606_,
		_w15607_
	);
	LUT2 #(
		.INIT('h4)
	) name15574 (
		_w15604_,
		_w15607_,
		_w15608_
	);
	LUT3 #(
		.INIT('h9a)
	) name15575 (
		\a[20] ,
		_w15603_,
		_w15608_,
		_w15609_
	);
	LUT3 #(
		.INIT('h31)
	) name15576 (
		_w15564_,
		_w15571_,
		_w15572_,
		_w15610_
	);
	LUT3 #(
		.INIT('h32)
	) name15577 (
		_w15527_,
		_w15561_,
		_w15562_,
		_w15611_
	);
	LUT4 #(
		.INIT('h0f01)
	) name15578 (
		_w15492_,
		_w15494_,
		_w15552_,
		_w15553_,
		_w15612_
	);
	LUT3 #(
		.INIT('h0d)
	) name15579 (
		_w15535_,
		_w15542_,
		_w15543_,
		_w15613_
	);
	LUT4 #(
		.INIT('h135f)
	) name15580 (
		_w90_,
		_w41_,
		_w72_,
		_w378_,
		_w15614_
	);
	LUT4 #(
		.INIT('h8000)
	) name15581 (
		_w670_,
		_w687_,
		_w1281_,
		_w15614_,
		_w15615_
	);
	LUT4 #(
		.INIT('h0800)
	) name15582 (
		_w116_,
		_w343_,
		_w360_,
		_w1540_,
		_w15616_
	);
	LUT3 #(
		.INIT('h80)
	) name15583 (
		_w1374_,
		_w1754_,
		_w8343_,
		_w15617_
	);
	LUT4 #(
		.INIT('h8000)
	) name15584 (
		_w644_,
		_w15617_,
		_w15615_,
		_w15616_,
		_w15618_
	);
	LUT4 #(
		.INIT('h8000)
	) name15585 (
		_w3815_,
		_w3816_,
		_w7595_,
		_w7598_,
		_w15619_
	);
	LUT3 #(
		.INIT('h80)
	) name15586 (
		_w3446_,
		_w15618_,
		_w15619_,
		_w15620_
	);
	LUT2 #(
		.INIT('h8)
	) name15587 (
		_w2273_,
		_w15620_,
		_w15621_
	);
	LUT4 #(
		.INIT('h0df2)
	) name15588 (
		_w15535_,
		_w15542_,
		_w15543_,
		_w15621_,
		_w15622_
	);
	LUT3 #(
		.INIT('h82)
	) name15589 (
		_w377_,
		_w11484_,
		_w11486_,
		_w15623_
	);
	LUT3 #(
		.INIT('h82)
	) name15590 (
		_w2527_,
		_w11280_,
		_w11282_,
		_w15624_
	);
	LUT2 #(
		.INIT('h8)
	) name15591 (
		_w376_,
		_w11388_,
		_w15625_
	);
	LUT4 #(
		.INIT('h2228)
	) name15592 (
		_w2407_,
		_w7935_,
		_w8077_,
		_w11279_,
		_w15626_
	);
	LUT2 #(
		.INIT('h1)
	) name15593 (
		_w15625_,
		_w15626_,
		_w15627_
	);
	LUT2 #(
		.INIT('h4)
	) name15594 (
		_w15624_,
		_w15627_,
		_w15628_
	);
	LUT2 #(
		.INIT('h4)
	) name15595 (
		_w15623_,
		_w15628_,
		_w15629_
	);
	LUT4 #(
		.INIT('h147d)
	) name15596 (
		_w15534_,
		_w15535_,
		_w15544_,
		_w15550_,
		_w15630_
	);
	LUT3 #(
		.INIT('h82)
	) name15597 (
		_w2550_,
		_w11490_,
		_w11492_,
		_w15631_
	);
	LUT3 #(
		.INIT('h82)
	) name15598 (
		_w2854_,
		_w11286_,
		_w11335_,
		_w15632_
	);
	LUT2 #(
		.INIT('h8)
	) name15599 (
		_w2549_,
		_w11382_,
		_w15633_
	);
	LUT4 #(
		.INIT('h2228)
	) name15600 (
		_w2617_,
		_w7695_,
		_w7750_,
		_w11285_,
		_w15634_
	);
	LUT2 #(
		.INIT('h1)
	) name15601 (
		_w15633_,
		_w15634_,
		_w15635_
	);
	LUT2 #(
		.INIT('h4)
	) name15602 (
		_w15632_,
		_w15635_,
		_w15636_
	);
	LUT3 #(
		.INIT('h9a)
	) name15603 (
		\a[29] ,
		_w15631_,
		_w15636_,
		_w15637_
	);
	LUT4 #(
		.INIT('h6996)
	) name15604 (
		_w15622_,
		_w15629_,
		_w15630_,
		_w15637_,
		_w15638_
	);
	LUT3 #(
		.INIT('h82)
	) name15605 (
		_w2875_,
		_w13061_,
		_w13102_,
		_w15639_
	);
	LUT3 #(
		.INIT('h82)
	) name15606 (
		_w2986_,
		_w13062_,
		_w13099_,
		_w15640_
	);
	LUT2 #(
		.INIT('h8)
	) name15607 (
		_w2874_,
		_w11377_,
		_w15641_
	);
	LUT4 #(
		.INIT('h2228)
	) name15608 (
		_w2975_,
		_w11549_,
		_w11373_,
		_w11375_,
		_w15642_
	);
	LUT2 #(
		.INIT('h1)
	) name15609 (
		_w15641_,
		_w15642_,
		_w15643_
	);
	LUT2 #(
		.INIT('h4)
	) name15610 (
		_w15640_,
		_w15643_,
		_w15644_
	);
	LUT3 #(
		.INIT('h9a)
	) name15611 (
		\a[26] ,
		_w15639_,
		_w15644_,
		_w15645_
	);
	LUT3 #(
		.INIT('h96)
	) name15612 (
		_w15612_,
		_w15638_,
		_w15645_,
		_w15646_
	);
	LUT3 #(
		.INIT('h82)
	) name15613 (
		_w37_,
		_w13292_,
		_w13325_,
		_w15647_
	);
	LUT3 #(
		.INIT('h82)
	) name15614 (
		_w3262_,
		_w13293_,
		_w13322_,
		_w15648_
	);
	LUT2 #(
		.INIT('h8)
	) name15615 (
		_w3214_,
		_w13247_,
		_w15649_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15616 (
		_w3249_,
		_w13243_,
		_w13245_,
		_w13285_,
		_w15650_
	);
	LUT2 #(
		.INIT('h1)
	) name15617 (
		_w15649_,
		_w15650_,
		_w15651_
	);
	LUT2 #(
		.INIT('h4)
	) name15618 (
		_w15648_,
		_w15651_,
		_w15652_
	);
	LUT3 #(
		.INIT('h9a)
	) name15619 (
		\a[23] ,
		_w15647_,
		_w15652_,
		_w15653_
	);
	LUT3 #(
		.INIT('h96)
	) name15620 (
		_w15611_,
		_w15646_,
		_w15653_,
		_w15654_
	);
	LUT3 #(
		.INIT('h96)
	) name15621 (
		_w15609_,
		_w15610_,
		_w15654_,
		_w15655_
	);
	LUT3 #(
		.INIT('h82)
	) name15622 (
		_w3710_,
		_w14343_,
		_w14349_,
		_w15656_
	);
	LUT3 #(
		.INIT('h28)
	) name15623 (
		_w3886_,
		_w14344_,
		_w14347_,
		_w15657_
	);
	LUT2 #(
		.INIT('h8)
	) name15624 (
		_w3709_,
		_w14112_,
		_w15658_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15625 (
		_w3877_,
		_w14108_,
		_w14111_,
		_w14235_,
		_w15659_
	);
	LUT2 #(
		.INIT('h1)
	) name15626 (
		_w15658_,
		_w15659_,
		_w15660_
	);
	LUT2 #(
		.INIT('h4)
	) name15627 (
		_w15657_,
		_w15660_,
		_w15661_
	);
	LUT3 #(
		.INIT('h9a)
	) name15628 (
		\a[17] ,
		_w15656_,
		_w15661_,
		_w15662_
	);
	LUT3 #(
		.INIT('h96)
	) name15629 (
		_w15602_,
		_w15655_,
		_w15662_,
		_w15663_
	);
	LUT4 #(
		.INIT('hb200)
	) name15630 (
		_w15584_,
		_w15590_,
		_w15591_,
		_w15663_,
		_w15664_
	);
	LUT4 #(
		.INIT('h31ce)
	) name15631 (
		_w15584_,
		_w15592_,
		_w15593_,
		_w15663_,
		_w15665_
	);
	LUT4 #(
		.INIT('hd400)
	) name15632 (
		_w15526_,
		_w15595_,
		_w15596_,
		_w15665_,
		_w15666_
	);
	LUT4 #(
		.INIT('h32cd)
	) name15633 (
		_w15526_,
		_w15597_,
		_w15598_,
		_w15665_,
		_w15667_
	);
	LUT2 #(
		.INIT('h8)
	) name15634 (
		_w15600_,
		_w15667_,
		_w15668_
	);
	LUT2 #(
		.INIT('h6)
	) name15635 (
		_w15600_,
		_w15667_,
		_w15669_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name15636 (
		_w3710_,
		_w14343_,
		_w14348_,
		_w14349_,
		_w15670_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15637 (
		_w3709_,
		_w14108_,
		_w14111_,
		_w14235_,
		_w15671_
	);
	LUT4 #(
		.INIT('h00eb)
	) name15638 (
		_w7753_,
		_w14344_,
		_w14347_,
		_w15671_,
		_w15672_
	);
	LUT3 #(
		.INIT('h9a)
	) name15639 (
		\a[17] ,
		_w15670_,
		_w15672_,
		_w15673_
	);
	LUT4 #(
		.INIT('h0071)
	) name15640 (
		_w15609_,
		_w15610_,
		_w15654_,
		_w15673_,
		_w15674_
	);
	LUT4 #(
		.INIT('h8e00)
	) name15641 (
		_w15609_,
		_w15610_,
		_w15654_,
		_w15673_,
		_w15675_
	);
	LUT4 #(
		.INIT('h718e)
	) name15642 (
		_w15609_,
		_w15610_,
		_w15654_,
		_w15673_,
		_w15676_
	);
	LUT4 #(
		.INIT('h6f06)
	) name15643 (
		_w15622_,
		_w15629_,
		_w15630_,
		_w15637_,
		_w15677_
	);
	LUT4 #(
		.INIT('h2228)
	) name15644 (
		_w2549_,
		_w7695_,
		_w7750_,
		_w11285_,
		_w15678_
	);
	LUT4 #(
		.INIT('h007d)
	) name15645 (
		_w2617_,
		_w11286_,
		_w11335_,
		_w15678_,
		_w15679_
	);
	LUT3 #(
		.INIT('h70)
	) name15646 (
		_w2854_,
		_w11377_,
		_w15679_,
		_w15680_
	);
	LUT4 #(
		.INIT('h95aa)
	) name15647 (
		\a[29] ,
		_w2550_,
		_w12799_,
		_w15680_,
		_w15681_
	);
	LUT4 #(
		.INIT('h135f)
	) name15648 (
		_w52_,
		_w67_,
		_w236_,
		_w378_,
		_w15682_
	);
	LUT2 #(
		.INIT('h8)
	) name15649 (
		_w1403_,
		_w15682_,
		_w15683_
	);
	LUT4 #(
		.INIT('h0777)
	) name15650 (
		_w52_,
		_w72_,
		_w39_,
		_w46_,
		_w15684_
	);
	LUT4 #(
		.INIT('h153f)
	) name15651 (
		_w59_,
		_w78_,
		_w44_,
		_w430_,
		_w15685_
	);
	LUT4 #(
		.INIT('h8000)
	) name15652 (
		_w861_,
		_w1514_,
		_w15684_,
		_w15685_,
		_w15686_
	);
	LUT2 #(
		.INIT('h8)
	) name15653 (
		_w15683_,
		_w15686_,
		_w15687_
	);
	LUT4 #(
		.INIT('h8000)
	) name15654 (
		_w951_,
		_w1001_,
		_w1761_,
		_w1871_,
		_w15688_
	);
	LUT3 #(
		.INIT('h80)
	) name15655 (
		_w581_,
		_w2113_,
		_w15688_,
		_w15689_
	);
	LUT3 #(
		.INIT('h80)
	) name15656 (
		_w2508_,
		_w15687_,
		_w15689_,
		_w15690_
	);
	LUT4 #(
		.INIT('h8000)
	) name15657 (
		_w1336_,
		_w1349_,
		_w3171_,
		_w3556_,
		_w15691_
	);
	LUT2 #(
		.INIT('h8)
	) name15658 (
		_w15690_,
		_w15691_,
		_w15692_
	);
	LUT4 #(
		.INIT('h817e)
	) name15659 (
		_w15613_,
		_w15621_,
		_w15629_,
		_w15692_,
		_w15693_
	);
	LUT4 #(
		.INIT('h2228)
	) name15660 (
		_w376_,
		_w7935_,
		_w8077_,
		_w11279_,
		_w15694_
	);
	LUT4 #(
		.INIT('h007d)
	) name15661 (
		_w2407_,
		_w11280_,
		_w11282_,
		_w15694_,
		_w15695_
	);
	LUT3 #(
		.INIT('h70)
	) name15662 (
		_w2527_,
		_w11382_,
		_w15695_,
		_w15696_
	);
	LUT3 #(
		.INIT('h70)
	) name15663 (
		_w377_,
		_w12476_,
		_w15696_,
		_w15697_
	);
	LUT3 #(
		.INIT('h96)
	) name15664 (
		_w15681_,
		_w15693_,
		_w15697_,
		_w15698_
	);
	LUT4 #(
		.INIT('h4114)
	) name15665 (
		_w15677_,
		_w15681_,
		_w15693_,
		_w15697_,
		_w15699_
	);
	LUT4 #(
		.INIT('h2882)
	) name15666 (
		_w15677_,
		_w15681_,
		_w15693_,
		_w15697_,
		_w15700_
	);
	LUT4 #(
		.INIT('h9669)
	) name15667 (
		_w15677_,
		_w15681_,
		_w15693_,
		_w15697_,
		_w15701_
	);
	LUT4 #(
		.INIT('h2228)
	) name15668 (
		_w2874_,
		_w11549_,
		_w11373_,
		_w11375_,
		_w15702_
	);
	LUT4 #(
		.INIT('h007d)
	) name15669 (
		_w2975_,
		_w13062_,
		_w13099_,
		_w15702_,
		_w15703_
	);
	LUT3 #(
		.INIT('h70)
	) name15670 (
		_w2986_,
		_w13247_,
		_w15703_,
		_w15704_
	);
	LUT4 #(
		.INIT('h95aa)
	) name15671 (
		\a[26] ,
		_w2875_,
		_w13576_,
		_w15704_,
		_w15705_
	);
	LUT2 #(
		.INIT('h9)
	) name15672 (
		_w15701_,
		_w15705_,
		_w15706_
	);
	LUT3 #(
		.INIT('h4d)
	) name15673 (
		_w15612_,
		_w15638_,
		_w15645_,
		_w15707_
	);
	LUT4 #(
		.INIT('h00b2)
	) name15674 (
		_w15612_,
		_w15638_,
		_w15645_,
		_w15706_,
		_w15708_
	);
	LUT4 #(
		.INIT('h4d00)
	) name15675 (
		_w15612_,
		_w15638_,
		_w15645_,
		_w15706_,
		_w15709_
	);
	LUT4 #(
		.INIT('hb24d)
	) name15676 (
		_w15612_,
		_w15638_,
		_w15645_,
		_w15706_,
		_w15710_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15677 (
		_w3214_,
		_w13243_,
		_w13245_,
		_w13285_,
		_w15711_
	);
	LUT4 #(
		.INIT('h007d)
	) name15678 (
		_w3249_,
		_w13293_,
		_w13322_,
		_w15711_,
		_w15712_
	);
	LUT3 #(
		.INIT('h70)
	) name15679 (
		_w3262_,
		_w13716_,
		_w15712_,
		_w15713_
	);
	LUT4 #(
		.INIT('h95aa)
	) name15680 (
		\a[23] ,
		_w37_,
		_w13720_,
		_w15713_,
		_w15714_
	);
	LUT2 #(
		.INIT('h9)
	) name15681 (
		_w15710_,
		_w15714_,
		_w15715_
	);
	LUT3 #(
		.INIT('h4d)
	) name15682 (
		_w15611_,
		_w15646_,
		_w15653_,
		_w15716_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15683 (
		_w3311_,
		_w13712_,
		_w13714_,
		_w13847_,
		_w15717_
	);
	LUT4 #(
		.INIT('h007d)
	) name15684 (
		_w3645_,
		_w13960_,
		_w13979_,
		_w15717_,
		_w15718_
	);
	LUT3 #(
		.INIT('h70)
	) name15685 (
		_w3654_,
		_w14112_,
		_w15718_,
		_w15719_
	);
	LUT4 #(
		.INIT('h95aa)
	) name15686 (
		\a[20] ,
		_w3312_,
		_w14116_,
		_w15719_,
		_w15720_
	);
	LUT3 #(
		.INIT('h69)
	) name15687 (
		_w15715_,
		_w15716_,
		_w15720_,
		_w15721_
	);
	LUT2 #(
		.INIT('h6)
	) name15688 (
		_w15676_,
		_w15721_,
		_w15722_
	);
	LUT3 #(
		.INIT('h4d)
	) name15689 (
		_w15602_,
		_w15655_,
		_w15662_,
		_w15723_
	);
	LUT2 #(
		.INIT('h8)
	) name15690 (
		_w15722_,
		_w15723_,
		_w15724_
	);
	LUT2 #(
		.INIT('h6)
	) name15691 (
		_w15722_,
		_w15723_,
		_w15725_
	);
	LUT3 #(
		.INIT('h1e)
	) name15692 (
		_w15664_,
		_w15666_,
		_w15725_,
		_w15726_
	);
	LUT2 #(
		.INIT('h6)
	) name15693 (
		_w15668_,
		_w15726_,
		_w15727_
	);
	LUT4 #(
		.INIT('h010f)
	) name15694 (
		_w15664_,
		_w15666_,
		_w15724_,
		_w15725_,
		_w15728_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15695 (
		_w37_,
		_w13717_,
		_w13719_,
		_w13850_,
		_w15729_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15696 (
		_w3262_,
		_w13712_,
		_w13714_,
		_w13847_,
		_w15730_
	);
	LUT3 #(
		.INIT('h82)
	) name15697 (
		_w3214_,
		_w13293_,
		_w13322_,
		_w15731_
	);
	LUT3 #(
		.INIT('h07)
	) name15698 (
		_w3249_,
		_w13716_,
		_w15731_,
		_w15732_
	);
	LUT2 #(
		.INIT('h4)
	) name15699 (
		_w15730_,
		_w15732_,
		_w15733_
	);
	LUT3 #(
		.INIT('h9a)
	) name15700 (
		\a[23] ,
		_w15729_,
		_w15733_,
		_w15734_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15701 (
		_w2875_,
		_w13288_,
		_w13290_,
		_w13291_,
		_w15735_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15702 (
		_w2986_,
		_w13243_,
		_w13245_,
		_w13285_,
		_w15736_
	);
	LUT3 #(
		.INIT('h82)
	) name15703 (
		_w2874_,
		_w13062_,
		_w13099_,
		_w15737_
	);
	LUT3 #(
		.INIT('h07)
	) name15704 (
		_w2975_,
		_w13247_,
		_w15737_,
		_w15738_
	);
	LUT2 #(
		.INIT('h4)
	) name15705 (
		_w15736_,
		_w15738_,
		_w15739_
	);
	LUT3 #(
		.INIT('h9a)
	) name15706 (
		\a[26] ,
		_w15735_,
		_w15739_,
		_w15740_
	);
	LUT4 #(
		.INIT('h004d)
	) name15707 (
		_w15677_,
		_w15698_,
		_w15705_,
		_w15740_,
		_w15741_
	);
	LUT4 #(
		.INIT('hb200)
	) name15708 (
		_w15677_,
		_w15698_,
		_w15705_,
		_w15740_,
		_w15742_
	);
	LUT4 #(
		.INIT('h23dc)
	) name15709 (
		_w15699_,
		_w15700_,
		_w15705_,
		_w15740_,
		_w15743_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15710 (
		_w2550_,
		_w11378_,
		_w11494_,
		_w11552_,
		_w15744_
	);
	LUT4 #(
		.INIT('h2228)
	) name15711 (
		_w2854_,
		_w11549_,
		_w11373_,
		_w11375_,
		_w15745_
	);
	LUT3 #(
		.INIT('h82)
	) name15712 (
		_w2549_,
		_w11286_,
		_w11335_,
		_w15746_
	);
	LUT3 #(
		.INIT('h07)
	) name15713 (
		_w2617_,
		_w11377_,
		_w15746_,
		_w15747_
	);
	LUT2 #(
		.INIT('h4)
	) name15714 (
		_w15745_,
		_w15747_,
		_w15748_
	);
	LUT3 #(
		.INIT('h9a)
	) name15715 (
		\a[29] ,
		_w15744_,
		_w15748_,
		_w15749_
	);
	LUT3 #(
		.INIT('hb2)
	) name15716 (
		_w15681_,
		_w15693_,
		_w15697_,
		_w15750_
	);
	LUT4 #(
		.INIT('h80fe)
	) name15717 (
		_w15613_,
		_w15621_,
		_w15629_,
		_w15692_,
		_w15751_
	);
	LUT4 #(
		.INIT('h5665)
	) name15718 (
		\a[17] ,
		_w7245_,
		_w14344_,
		_w14347_,
		_w15752_
	);
	LUT4 #(
		.INIT('h153f)
	) name15719 (
		_w47_,
		_w39_,
		_w46_,
		_w201_,
		_w15753_
	);
	LUT4 #(
		.INIT('h4000)
	) name15720 (
		_w295_,
		_w966_,
		_w1211_,
		_w15753_,
		_w15754_
	);
	LUT4 #(
		.INIT('h8000)
	) name15721 (
		_w584_,
		_w663_,
		_w1352_,
		_w12732_,
		_w15755_
	);
	LUT2 #(
		.INIT('h8)
	) name15722 (
		_w15754_,
		_w15755_,
		_w15756_
	);
	LUT3 #(
		.INIT('h80)
	) name15723 (
		_w1217_,
		_w2278_,
		_w7193_,
		_w15757_
	);
	LUT3 #(
		.INIT('h80)
	) name15724 (
		_w994_,
		_w15756_,
		_w15757_,
		_w15758_
	);
	LUT4 #(
		.INIT('h8000)
	) name15725 (
		_w2900_,
		_w2909_,
		_w3344_,
		_w3348_,
		_w15759_
	);
	LUT2 #(
		.INIT('h8)
	) name15726 (
		_w15758_,
		_w15759_,
		_w15760_
	);
	LUT4 #(
		.INIT('h8000)
	) name15727 (
		_w15690_,
		_w15691_,
		_w15758_,
		_w15759_,
		_w15761_
	);
	LUT4 #(
		.INIT('h0777)
	) name15728 (
		_w15690_,
		_w15691_,
		_w15758_,
		_w15759_,
		_w15762_
	);
	LUT4 #(
		.INIT('h7888)
	) name15729 (
		_w15690_,
		_w15691_,
		_w15758_,
		_w15759_,
		_w15763_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15730 (
		_w377_,
		_w11384_,
		_w11488_,
		_w11489_,
		_w15764_
	);
	LUT4 #(
		.INIT('h2228)
	) name15731 (
		_w2527_,
		_w7695_,
		_w7750_,
		_w11285_,
		_w15765_
	);
	LUT3 #(
		.INIT('h82)
	) name15732 (
		_w376_,
		_w11280_,
		_w11282_,
		_w15766_
	);
	LUT3 #(
		.INIT('h07)
	) name15733 (
		_w2407_,
		_w11382_,
		_w15766_,
		_w15767_
	);
	LUT2 #(
		.INIT('h4)
	) name15734 (
		_w15765_,
		_w15767_,
		_w15768_
	);
	LUT2 #(
		.INIT('h4)
	) name15735 (
		_w15764_,
		_w15768_,
		_w15769_
	);
	LUT3 #(
		.INIT('h06)
	) name15736 (
		_w15752_,
		_w15763_,
		_w15769_,
		_w15770_
	);
	LUT3 #(
		.INIT('h90)
	) name15737 (
		_w15752_,
		_w15763_,
		_w15769_,
		_w15771_
	);
	LUT3 #(
		.INIT('h69)
	) name15738 (
		_w15752_,
		_w15763_,
		_w15769_,
		_w15772_
	);
	LUT2 #(
		.INIT('h9)
	) name15739 (
		_w15751_,
		_w15772_,
		_w15773_
	);
	LUT3 #(
		.INIT('h96)
	) name15740 (
		_w15749_,
		_w15750_,
		_w15773_,
		_w15774_
	);
	LUT3 #(
		.INIT('h14)
	) name15741 (
		_w15734_,
		_w15743_,
		_w15774_,
		_w15775_
	);
	LUT3 #(
		.INIT('h69)
	) name15742 (
		_w15734_,
		_w15743_,
		_w15774_,
		_w15776_
	);
	LUT4 #(
		.INIT('h8e00)
	) name15743 (
		_w15706_,
		_w15707_,
		_w15714_,
		_w15776_,
		_w15777_
	);
	LUT4 #(
		.INIT('hba45)
	) name15744 (
		_w15708_,
		_w15709_,
		_w15714_,
		_w15776_,
		_w15778_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15745 (
		_w3312_,
		_w14113_,
		_w14115_,
		_w14238_,
		_w15779_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15746 (
		_w3654_,
		_w14108_,
		_w14111_,
		_w14235_,
		_w15780_
	);
	LUT3 #(
		.INIT('h82)
	) name15747 (
		_w3311_,
		_w13960_,
		_w13979_,
		_w15781_
	);
	LUT3 #(
		.INIT('h07)
	) name15748 (
		_w3645_,
		_w14112_,
		_w15781_,
		_w15782_
	);
	LUT2 #(
		.INIT('h4)
	) name15749 (
		_w15780_,
		_w15782_,
		_w15783_
	);
	LUT3 #(
		.INIT('h9a)
	) name15750 (
		\a[20] ,
		_w15779_,
		_w15783_,
		_w15784_
	);
	LUT3 #(
		.INIT('h8e)
	) name15751 (
		_w15715_,
		_w15716_,
		_w15720_,
		_w15785_
	);
	LUT4 #(
		.INIT('h008e)
	) name15752 (
		_w15715_,
		_w15716_,
		_w15720_,
		_w15784_,
		_w15786_
	);
	LUT4 #(
		.INIT('h7100)
	) name15753 (
		_w15715_,
		_w15716_,
		_w15720_,
		_w15784_,
		_w15787_
	);
	LUT4 #(
		.INIT('h8e71)
	) name15754 (
		_w15715_,
		_w15716_,
		_w15720_,
		_w15784_,
		_w15788_
	);
	LUT2 #(
		.INIT('h6)
	) name15755 (
		_w15778_,
		_w15788_,
		_w15789_
	);
	LUT3 #(
		.INIT('h32)
	) name15756 (
		_w15674_,
		_w15675_,
		_w15721_,
		_w15790_
	);
	LUT2 #(
		.INIT('h8)
	) name15757 (
		_w15789_,
		_w15790_,
		_w15791_
	);
	LUT2 #(
		.INIT('h1)
	) name15758 (
		_w15789_,
		_w15790_,
		_w15792_
	);
	LUT2 #(
		.INIT('h6)
	) name15759 (
		_w15789_,
		_w15790_,
		_w15793_
	);
	LUT4 #(
		.INIT('h8008)
	) name15760 (
		_w15668_,
		_w15726_,
		_w15728_,
		_w15793_,
		_w15794_
	);
	LUT4 #(
		.INIT('h7887)
	) name15761 (
		_w15668_,
		_w15726_,
		_w15728_,
		_w15793_,
		_w15795_
	);
	LUT3 #(
		.INIT('h82)
	) name15762 (
		_w37_,
		_w13959_,
		_w13982_,
		_w15796_
	);
	LUT3 #(
		.INIT('h82)
	) name15763 (
		_w3262_,
		_w13960_,
		_w13979_,
		_w15797_
	);
	LUT2 #(
		.INIT('h8)
	) name15764 (
		_w3214_,
		_w13716_,
		_w15798_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15765 (
		_w3249_,
		_w13712_,
		_w13714_,
		_w13847_,
		_w15799_
	);
	LUT2 #(
		.INIT('h1)
	) name15766 (
		_w15798_,
		_w15799_,
		_w15800_
	);
	LUT2 #(
		.INIT('h4)
	) name15767 (
		_w15797_,
		_w15800_,
		_w15801_
	);
	LUT3 #(
		.INIT('h9a)
	) name15768 (
		\a[23] ,
		_w15796_,
		_w15801_,
		_w15802_
	);
	LUT3 #(
		.INIT('h45)
	) name15769 (
		_w15741_,
		_w15742_,
		_w15774_,
		_w15803_
	);
	LUT3 #(
		.INIT('h32)
	) name15770 (
		_w15751_,
		_w15770_,
		_w15771_,
		_w15804_
	);
	LUT3 #(
		.INIT('h0d)
	) name15771 (
		_w15752_,
		_w15761_,
		_w15762_,
		_w15805_
	);
	LUT3 #(
		.INIT('h80)
	) name15772 (
		_w997_,
		_w1082_,
		_w3022_,
		_w15806_
	);
	LUT4 #(
		.INIT('h0777)
	) name15773 (
		_w122_,
		_w59_,
		_w50_,
		_w166_,
		_w15807_
	);
	LUT4 #(
		.INIT('h153f)
	) name15774 (
		_w38_,
		_w93_,
		_w166_,
		_w419_,
		_w15808_
	);
	LUT4 #(
		.INIT('h8000)
	) name15775 (
		_w820_,
		_w945_,
		_w15807_,
		_w15808_,
		_w15809_
	);
	LUT4 #(
		.INIT('h4000)
	) name15776 (
		_w304_,
		_w1169_,
		_w1561_,
		_w2205_,
		_w15810_
	);
	LUT3 #(
		.INIT('h80)
	) name15777 (
		_w15806_,
		_w15809_,
		_w15810_,
		_w15811_
	);
	LUT4 #(
		.INIT('h8000)
	) name15778 (
		_w787_,
		_w791_,
		_w2144_,
		_w2147_,
		_w15812_
	);
	LUT4 #(
		.INIT('h8000)
	) name15779 (
		_w1757_,
		_w4147_,
		_w15811_,
		_w15812_,
		_w15813_
	);
	LUT2 #(
		.INIT('h8)
	) name15780 (
		_w14976_,
		_w15813_,
		_w15814_
	);
	LUT4 #(
		.INIT('h4d00)
	) name15781 (
		_w15692_,
		_w15752_,
		_w15760_,
		_w15814_,
		_w15815_
	);
	LUT4 #(
		.INIT('h00b2)
	) name15782 (
		_w15692_,
		_w15752_,
		_w15760_,
		_w15814_,
		_w15816_
	);
	LUT4 #(
		.INIT('h0df2)
	) name15783 (
		_w15752_,
		_w15761_,
		_w15762_,
		_w15814_,
		_w15817_
	);
	LUT3 #(
		.INIT('h82)
	) name15784 (
		_w377_,
		_w11490_,
		_w11492_,
		_w15818_
	);
	LUT3 #(
		.INIT('h82)
	) name15785 (
		_w2527_,
		_w11286_,
		_w11335_,
		_w15819_
	);
	LUT2 #(
		.INIT('h8)
	) name15786 (
		_w376_,
		_w11382_,
		_w15820_
	);
	LUT4 #(
		.INIT('h2228)
	) name15787 (
		_w2407_,
		_w7695_,
		_w7750_,
		_w11285_,
		_w15821_
	);
	LUT2 #(
		.INIT('h1)
	) name15788 (
		_w15820_,
		_w15821_,
		_w15822_
	);
	LUT2 #(
		.INIT('h4)
	) name15789 (
		_w15819_,
		_w15822_,
		_w15823_
	);
	LUT2 #(
		.INIT('h4)
	) name15790 (
		_w15818_,
		_w15823_,
		_w15824_
	);
	LUT2 #(
		.INIT('h9)
	) name15791 (
		_w15817_,
		_w15824_,
		_w15825_
	);
	LUT4 #(
		.INIT('h0023)
	) name15792 (
		_w15751_,
		_w15770_,
		_w15772_,
		_w15825_,
		_w15826_
	);
	LUT4 #(
		.INIT('hdc00)
	) name15793 (
		_w15751_,
		_w15770_,
		_w15772_,
		_w15825_,
		_w15827_
	);
	LUT4 #(
		.INIT('h32cd)
	) name15794 (
		_w15751_,
		_w15770_,
		_w15771_,
		_w15825_,
		_w15828_
	);
	LUT3 #(
		.INIT('h82)
	) name15795 (
		_w2550_,
		_w13061_,
		_w13102_,
		_w15829_
	);
	LUT3 #(
		.INIT('h82)
	) name15796 (
		_w2854_,
		_w13062_,
		_w13099_,
		_w15830_
	);
	LUT2 #(
		.INIT('h8)
	) name15797 (
		_w2549_,
		_w11377_,
		_w15831_
	);
	LUT4 #(
		.INIT('h2228)
	) name15798 (
		_w2617_,
		_w11549_,
		_w11373_,
		_w11375_,
		_w15832_
	);
	LUT2 #(
		.INIT('h1)
	) name15799 (
		_w15831_,
		_w15832_,
		_w15833_
	);
	LUT2 #(
		.INIT('h4)
	) name15800 (
		_w15830_,
		_w15833_,
		_w15834_
	);
	LUT3 #(
		.INIT('h9a)
	) name15801 (
		\a[29] ,
		_w15829_,
		_w15834_,
		_w15835_
	);
	LUT2 #(
		.INIT('h9)
	) name15802 (
		_w15828_,
		_w15835_,
		_w15836_
	);
	LUT3 #(
		.INIT('h71)
	) name15803 (
		_w15749_,
		_w15750_,
		_w15773_,
		_w15837_
	);
	LUT3 #(
		.INIT('h82)
	) name15804 (
		_w2875_,
		_w13292_,
		_w13325_,
		_w15838_
	);
	LUT3 #(
		.INIT('h82)
	) name15805 (
		_w2986_,
		_w13293_,
		_w13322_,
		_w15839_
	);
	LUT2 #(
		.INIT('h8)
	) name15806 (
		_w2874_,
		_w13247_,
		_w15840_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15807 (
		_w2975_,
		_w13243_,
		_w13245_,
		_w13285_,
		_w15841_
	);
	LUT2 #(
		.INIT('h1)
	) name15808 (
		_w15840_,
		_w15841_,
		_w15842_
	);
	LUT2 #(
		.INIT('h4)
	) name15809 (
		_w15839_,
		_w15842_,
		_w15843_
	);
	LUT3 #(
		.INIT('h9a)
	) name15810 (
		\a[26] ,
		_w15838_,
		_w15843_,
		_w15844_
	);
	LUT3 #(
		.INIT('h69)
	) name15811 (
		_w15836_,
		_w15837_,
		_w15844_,
		_w15845_
	);
	LUT3 #(
		.INIT('h69)
	) name15812 (
		_w15802_,
		_w15803_,
		_w15845_,
		_w15846_
	);
	LUT3 #(
		.INIT('h82)
	) name15813 (
		_w3312_,
		_w14343_,
		_w14349_,
		_w15847_
	);
	LUT3 #(
		.INIT('h28)
	) name15814 (
		_w3654_,
		_w14344_,
		_w14347_,
		_w15848_
	);
	LUT2 #(
		.INIT('h8)
	) name15815 (
		_w3311_,
		_w14112_,
		_w15849_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15816 (
		_w3645_,
		_w14108_,
		_w14111_,
		_w14235_,
		_w15850_
	);
	LUT2 #(
		.INIT('h1)
	) name15817 (
		_w15849_,
		_w15850_,
		_w15851_
	);
	LUT2 #(
		.INIT('h4)
	) name15818 (
		_w15848_,
		_w15851_,
		_w15852_
	);
	LUT3 #(
		.INIT('h9a)
	) name15819 (
		\a[20] ,
		_w15847_,
		_w15852_,
		_w15853_
	);
	LUT4 #(
		.INIT('he11e)
	) name15820 (
		_w15775_,
		_w15777_,
		_w15846_,
		_w15853_,
		_w15854_
	);
	LUT4 #(
		.INIT('hb200)
	) name15821 (
		_w15778_,
		_w15784_,
		_w15785_,
		_w15854_,
		_w15855_
	);
	LUT4 #(
		.INIT('h31ce)
	) name15822 (
		_w15778_,
		_w15786_,
		_w15787_,
		_w15854_,
		_w15856_
	);
	LUT4 #(
		.INIT('hd400)
	) name15823 (
		_w15728_,
		_w15789_,
		_w15790_,
		_w15856_,
		_w15857_
	);
	LUT4 #(
		.INIT('h32cd)
	) name15824 (
		_w15728_,
		_w15791_,
		_w15792_,
		_w15856_,
		_w15858_
	);
	LUT2 #(
		.INIT('h8)
	) name15825 (
		_w15794_,
		_w15858_,
		_w15859_
	);
	LUT2 #(
		.INIT('h6)
	) name15826 (
		_w15794_,
		_w15858_,
		_w15860_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name15827 (
		_w3312_,
		_w14343_,
		_w14348_,
		_w14349_,
		_w15861_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15828 (
		_w3311_,
		_w14108_,
		_w14111_,
		_w14235_,
		_w15862_
	);
	LUT4 #(
		.INIT('h00d7)
	) name15829 (
		_w7421_,
		_w14344_,
		_w14347_,
		_w15862_,
		_w15863_
	);
	LUT3 #(
		.INIT('h9a)
	) name15830 (
		\a[20] ,
		_w15861_,
		_w15863_,
		_w15864_
	);
	LUT4 #(
		.INIT('h0071)
	) name15831 (
		_w15802_,
		_w15803_,
		_w15845_,
		_w15864_,
		_w15865_
	);
	LUT4 #(
		.INIT('h8e00)
	) name15832 (
		_w15802_,
		_w15803_,
		_w15845_,
		_w15864_,
		_w15866_
	);
	LUT4 #(
		.INIT('h718e)
	) name15833 (
		_w15802_,
		_w15803_,
		_w15845_,
		_w15864_,
		_w15867_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15834 (
		_w2874_,
		_w13243_,
		_w13245_,
		_w13285_,
		_w15868_
	);
	LUT4 #(
		.INIT('h007d)
	) name15835 (
		_w2975_,
		_w13293_,
		_w13322_,
		_w15868_,
		_w15869_
	);
	LUT3 #(
		.INIT('h70)
	) name15836 (
		_w2986_,
		_w13716_,
		_w15869_,
		_w15870_
	);
	LUT4 #(
		.INIT('h95aa)
	) name15837 (
		\a[26] ,
		_w2875_,
		_w13720_,
		_w15870_,
		_w15871_
	);
	LUT3 #(
		.INIT('h80)
	) name15838 (
		_w976_,
		_w2267_,
		_w7325_,
		_w15872_
	);
	LUT4 #(
		.INIT('h0777)
	) name15839 (
		_w122_,
		_w50_,
		_w44_,
		_w166_,
		_w15873_
	);
	LUT4 #(
		.INIT('h4000)
	) name15840 (
		_w478_,
		_w834_,
		_w7202_,
		_w15873_,
		_w15874_
	);
	LUT3 #(
		.INIT('h80)
	) name15841 (
		_w15683_,
		_w15872_,
		_w15874_,
		_w15875_
	);
	LUT4 #(
		.INIT('h8000)
	) name15842 (
		_w2902_,
		_w2905_,
		_w8368_,
		_w14583_,
		_w15876_
	);
	LUT4 #(
		.INIT('h8000)
	) name15843 (
		_w3168_,
		_w4174_,
		_w15875_,
		_w15876_,
		_w15877_
	);
	LUT4 #(
		.INIT('h40c0)
	) name15844 (
		_w1009_,
		_w14976_,
		_w15813_,
		_w15877_,
		_w15878_
	);
	LUT4 #(
		.INIT('h953f)
	) name15845 (
		_w1009_,
		_w14976_,
		_w15813_,
		_w15877_,
		_w15879_
	);
	LUT4 #(
		.INIT('h2228)
	) name15846 (
		_w376_,
		_w7695_,
		_w7750_,
		_w11285_,
		_w15880_
	);
	LUT4 #(
		.INIT('h007d)
	) name15847 (
		_w2407_,
		_w11286_,
		_w11335_,
		_w15880_,
		_w15881_
	);
	LUT3 #(
		.INIT('h70)
	) name15848 (
		_w2527_,
		_w11377_,
		_w15881_,
		_w15882_
	);
	LUT4 #(
		.INIT('h80f0)
	) name15849 (
		_w377_,
		_w12799_,
		_w15879_,
		_w15882_,
		_w15883_
	);
	LUT4 #(
		.INIT('h780f)
	) name15850 (
		_w377_,
		_w12799_,
		_w15879_,
		_w15882_,
		_w15884_
	);
	LUT4 #(
		.INIT('h4d00)
	) name15851 (
		_w15805_,
		_w15814_,
		_w15824_,
		_w15884_,
		_w15885_
	);
	LUT4 #(
		.INIT('hdc23)
	) name15852 (
		_w15815_,
		_w15816_,
		_w15824_,
		_w15884_,
		_w15886_
	);
	LUT4 #(
		.INIT('h4d00)
	) name15853 (
		_w15804_,
		_w15825_,
		_w15835_,
		_w15886_,
		_w15887_
	);
	LUT4 #(
		.INIT('h32cd)
	) name15854 (
		_w15826_,
		_w15827_,
		_w15835_,
		_w15886_,
		_w15888_
	);
	LUT4 #(
		.INIT('h2228)
	) name15855 (
		_w2549_,
		_w11549_,
		_w11373_,
		_w11375_,
		_w15889_
	);
	LUT4 #(
		.INIT('h007d)
	) name15856 (
		_w2617_,
		_w13062_,
		_w13099_,
		_w15889_,
		_w15890_
	);
	LUT3 #(
		.INIT('h70)
	) name15857 (
		_w2854_,
		_w13247_,
		_w15890_,
		_w15891_
	);
	LUT4 #(
		.INIT('h95aa)
	) name15858 (
		\a[29] ,
		_w2550_,
		_w13576_,
		_w15891_,
		_w15892_
	);
	LUT3 #(
		.INIT('h96)
	) name15859 (
		_w15871_,
		_w15888_,
		_w15892_,
		_w15893_
	);
	LUT3 #(
		.INIT('h8e)
	) name15860 (
		_w15836_,
		_w15837_,
		_w15844_,
		_w15894_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15861 (
		_w3214_,
		_w13712_,
		_w13714_,
		_w13847_,
		_w15895_
	);
	LUT4 #(
		.INIT('h007d)
	) name15862 (
		_w3249_,
		_w13960_,
		_w13979_,
		_w15895_,
		_w15896_
	);
	LUT3 #(
		.INIT('h70)
	) name15863 (
		_w3262_,
		_w14112_,
		_w15896_,
		_w15897_
	);
	LUT4 #(
		.INIT('h95aa)
	) name15864 (
		\a[23] ,
		_w37_,
		_w14116_,
		_w15897_,
		_w15898_
	);
	LUT3 #(
		.INIT('h69)
	) name15865 (
		_w15893_,
		_w15894_,
		_w15898_,
		_w15899_
	);
	LUT2 #(
		.INIT('h6)
	) name15866 (
		_w15867_,
		_w15899_,
		_w15900_
	);
	LUT4 #(
		.INIT('h0eef)
	) name15867 (
		_w15775_,
		_w15777_,
		_w15846_,
		_w15853_,
		_w15901_
	);
	LUT2 #(
		.INIT('h1)
	) name15868 (
		_w15900_,
		_w15901_,
		_w15902_
	);
	LUT2 #(
		.INIT('h8)
	) name15869 (
		_w15900_,
		_w15901_,
		_w15903_
	);
	LUT2 #(
		.INIT('h6)
	) name15870 (
		_w15900_,
		_w15901_,
		_w15904_
	);
	LUT3 #(
		.INIT('h1e)
	) name15871 (
		_w15855_,
		_w15857_,
		_w15904_,
		_w15905_
	);
	LUT2 #(
		.INIT('h6)
	) name15872 (
		_w15859_,
		_w15905_,
		_w15906_
	);
	LUT4 #(
		.INIT('h00f1)
	) name15873 (
		_w15855_,
		_w15857_,
		_w15902_,
		_w15903_,
		_w15907_
	);
	LUT3 #(
		.INIT('hb2)
	) name15874 (
		_w15871_,
		_w15888_,
		_w15892_,
		_w15908_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15875 (
		_w2875_,
		_w13717_,
		_w13719_,
		_w13850_,
		_w15909_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15876 (
		_w2986_,
		_w13712_,
		_w13714_,
		_w13847_,
		_w15910_
	);
	LUT3 #(
		.INIT('h82)
	) name15877 (
		_w2874_,
		_w13293_,
		_w13322_,
		_w15911_
	);
	LUT3 #(
		.INIT('h07)
	) name15878 (
		_w2975_,
		_w13716_,
		_w15911_,
		_w15912_
	);
	LUT2 #(
		.INIT('h4)
	) name15879 (
		_w15910_,
		_w15912_,
		_w15913_
	);
	LUT3 #(
		.INIT('h9a)
	) name15880 (
		\a[26] ,
		_w15909_,
		_w15913_,
		_w15914_
	);
	LUT2 #(
		.INIT('h1)
	) name15881 (
		_w15878_,
		_w15883_,
		_w15915_
	);
	LUT4 #(
		.INIT('h5665)
	) name15882 (
		\a[20] ,
		_w11301_,
		_w14344_,
		_w14347_,
		_w15916_
	);
	LUT3 #(
		.INIT('h80)
	) name15883 (
		_w828_,
		_w1156_,
		_w1310_,
		_w15917_
	);
	LUT4 #(
		.INIT('h135f)
	) name15884 (
		_w122_,
		_w56_,
		_w41_,
		_w236_,
		_w15918_
	);
	LUT4 #(
		.INIT('h135f)
	) name15885 (
		_w56_,
		_w65_,
		_w419_,
		_w430_,
		_w15919_
	);
	LUT4 #(
		.INIT('h8000)
	) name15886 (
		_w737_,
		_w809_,
		_w15918_,
		_w15919_,
		_w15920_
	);
	LUT4 #(
		.INIT('h8000)
	) name15887 (
		_w2113_,
		_w7852_,
		_w15917_,
		_w15920_,
		_w15921_
	);
	LUT3 #(
		.INIT('h20)
	) name15888 (
		_w126_,
		_w451_,
		_w689_,
		_w15922_
	);
	LUT4 #(
		.INIT('h8000)
	) name15889 (
		_w640_,
		_w2243_,
		_w8312_,
		_w15922_,
		_w15923_
	);
	LUT4 #(
		.INIT('h8000)
	) name15890 (
		_w1241_,
		_w1252_,
		_w15921_,
		_w15923_,
		_w15924_
	);
	LUT4 #(
		.INIT('h8000)
	) name15891 (
		_w3106_,
		_w14976_,
		_w15813_,
		_w15924_,
		_w15925_
	);
	LUT4 #(
		.INIT('h153f)
	) name15892 (
		_w3106_,
		_w14976_,
		_w15813_,
		_w15924_,
		_w15926_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name15893 (
		_w3106_,
		_w14976_,
		_w15813_,
		_w15924_,
		_w15927_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15894 (
		_w377_,
		_w11378_,
		_w11494_,
		_w11552_,
		_w15928_
	);
	LUT4 #(
		.INIT('h2228)
	) name15895 (
		_w2527_,
		_w11549_,
		_w11373_,
		_w11375_,
		_w15929_
	);
	LUT3 #(
		.INIT('h82)
	) name15896 (
		_w376_,
		_w11286_,
		_w11335_,
		_w15930_
	);
	LUT3 #(
		.INIT('h07)
	) name15897 (
		_w2407_,
		_w11377_,
		_w15930_,
		_w15931_
	);
	LUT2 #(
		.INIT('h4)
	) name15898 (
		_w15929_,
		_w15931_,
		_w15932_
	);
	LUT2 #(
		.INIT('h4)
	) name15899 (
		_w15928_,
		_w15932_,
		_w15933_
	);
	LUT4 #(
		.INIT('h6996)
	) name15900 (
		_w15915_,
		_w15916_,
		_w15927_,
		_w15933_,
		_w15934_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15901 (
		_w2550_,
		_w13288_,
		_w13290_,
		_w13291_,
		_w15935_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15902 (
		_w2854_,
		_w13243_,
		_w13245_,
		_w13285_,
		_w15936_
	);
	LUT3 #(
		.INIT('h82)
	) name15903 (
		_w2549_,
		_w13062_,
		_w13099_,
		_w15937_
	);
	LUT3 #(
		.INIT('h07)
	) name15904 (
		_w2617_,
		_w13247_,
		_w15937_,
		_w15938_
	);
	LUT2 #(
		.INIT('h4)
	) name15905 (
		_w15936_,
		_w15938_,
		_w15939_
	);
	LUT3 #(
		.INIT('h9a)
	) name15906 (
		\a[29] ,
		_w15935_,
		_w15939_,
		_w15940_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name15907 (
		_w15885_,
		_w15887_,
		_w15934_,
		_w15940_,
		_w15941_
	);
	LUT3 #(
		.INIT('h96)
	) name15908 (
		_w15908_,
		_w15914_,
		_w15941_,
		_w15942_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15909 (
		_w37_,
		_w14113_,
		_w14115_,
		_w14238_,
		_w15943_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15910 (
		_w3262_,
		_w14108_,
		_w14111_,
		_w14235_,
		_w15944_
	);
	LUT3 #(
		.INIT('h82)
	) name15911 (
		_w3214_,
		_w13960_,
		_w13979_,
		_w15945_
	);
	LUT3 #(
		.INIT('h07)
	) name15912 (
		_w3249_,
		_w14112_,
		_w15945_,
		_w15946_
	);
	LUT2 #(
		.INIT('h4)
	) name15913 (
		_w15944_,
		_w15946_,
		_w15947_
	);
	LUT3 #(
		.INIT('h9a)
	) name15914 (
		\a[23] ,
		_w15943_,
		_w15947_,
		_w15948_
	);
	LUT4 #(
		.INIT('h008e)
	) name15915 (
		_w15893_,
		_w15894_,
		_w15898_,
		_w15948_,
		_w15949_
	);
	LUT4 #(
		.INIT('h7100)
	) name15916 (
		_w15893_,
		_w15894_,
		_w15898_,
		_w15948_,
		_w15950_
	);
	LUT4 #(
		.INIT('h8e71)
	) name15917 (
		_w15893_,
		_w15894_,
		_w15898_,
		_w15948_,
		_w15951_
	);
	LUT2 #(
		.INIT('h6)
	) name15918 (
		_w15942_,
		_w15951_,
		_w15952_
	);
	LUT3 #(
		.INIT('h32)
	) name15919 (
		_w15865_,
		_w15866_,
		_w15899_,
		_w15953_
	);
	LUT2 #(
		.INIT('h8)
	) name15920 (
		_w15952_,
		_w15953_,
		_w15954_
	);
	LUT2 #(
		.INIT('h1)
	) name15921 (
		_w15952_,
		_w15953_,
		_w15955_
	);
	LUT2 #(
		.INIT('h6)
	) name15922 (
		_w15952_,
		_w15953_,
		_w15956_
	);
	LUT4 #(
		.INIT('h8008)
	) name15923 (
		_w15859_,
		_w15905_,
		_w15907_,
		_w15956_,
		_w15957_
	);
	LUT4 #(
		.INIT('h7887)
	) name15924 (
		_w15859_,
		_w15905_,
		_w15907_,
		_w15956_,
		_w15958_
	);
	LUT3 #(
		.INIT('h31)
	) name15925 (
		_w15942_,
		_w15949_,
		_w15950_,
		_w15959_
	);
	LUT3 #(
		.INIT('h8e)
	) name15926 (
		_w15908_,
		_w15914_,
		_w15941_,
		_w15960_
	);
	LUT3 #(
		.INIT('h0d)
	) name15927 (
		_w15916_,
		_w15925_,
		_w15926_,
		_w15961_
	);
	LUT4 #(
		.INIT('h0777)
	) name15928 (
		_w122_,
		_w52_,
		_w90_,
		_w236_,
		_w15962_
	);
	LUT4 #(
		.INIT('h4000)
	) name15929 (
		_w407_,
		_w1401_,
		_w1625_,
		_w15962_,
		_w15963_
	);
	LUT3 #(
		.INIT('h80)
	) name15930 (
		_w1704_,
		_w3336_,
		_w3520_,
		_w15964_
	);
	LUT4 #(
		.INIT('h8000)
	) name15931 (
		_w833_,
		_w1646_,
		_w15964_,
		_w15963_,
		_w15965_
	);
	LUT4 #(
		.INIT('h8000)
	) name15932 (
		_w1317_,
		_w2230_,
		_w2742_,
		_w8344_,
		_w15966_
	);
	LUT4 #(
		.INIT('h8000)
	) name15933 (
		_w1672_,
		_w7606_,
		_w15965_,
		_w15966_,
		_w15967_
	);
	LUT2 #(
		.INIT('h8)
	) name15934 (
		_w2910_,
		_w15967_,
		_w15968_
	);
	LUT4 #(
		.INIT('h0df2)
	) name15935 (
		_w15916_,
		_w15925_,
		_w15926_,
		_w15968_,
		_w15969_
	);
	LUT3 #(
		.INIT('h82)
	) name15936 (
		_w377_,
		_w13061_,
		_w13102_,
		_w15970_
	);
	LUT3 #(
		.INIT('h82)
	) name15937 (
		_w2527_,
		_w13062_,
		_w13099_,
		_w15971_
	);
	LUT2 #(
		.INIT('h8)
	) name15938 (
		_w376_,
		_w11377_,
		_w15972_
	);
	LUT4 #(
		.INIT('h2228)
	) name15939 (
		_w2407_,
		_w11549_,
		_w11373_,
		_w11375_,
		_w15973_
	);
	LUT2 #(
		.INIT('h1)
	) name15940 (
		_w15972_,
		_w15973_,
		_w15974_
	);
	LUT2 #(
		.INIT('h4)
	) name15941 (
		_w15971_,
		_w15974_,
		_w15975_
	);
	LUT2 #(
		.INIT('h4)
	) name15942 (
		_w15970_,
		_w15975_,
		_w15976_
	);
	LUT4 #(
		.INIT('h147d)
	) name15943 (
		_w15915_,
		_w15916_,
		_w15927_,
		_w15933_,
		_w15977_
	);
	LUT3 #(
		.INIT('h82)
	) name15944 (
		_w2550_,
		_w13292_,
		_w13325_,
		_w15978_
	);
	LUT3 #(
		.INIT('h82)
	) name15945 (
		_w2854_,
		_w13293_,
		_w13322_,
		_w15979_
	);
	LUT2 #(
		.INIT('h8)
	) name15946 (
		_w2549_,
		_w13247_,
		_w15980_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15947 (
		_w2617_,
		_w13243_,
		_w13245_,
		_w13285_,
		_w15981_
	);
	LUT2 #(
		.INIT('h1)
	) name15948 (
		_w15980_,
		_w15981_,
		_w15982_
	);
	LUT2 #(
		.INIT('h4)
	) name15949 (
		_w15979_,
		_w15982_,
		_w15983_
	);
	LUT3 #(
		.INIT('h9a)
	) name15950 (
		\a[29] ,
		_w15978_,
		_w15983_,
		_w15984_
	);
	LUT4 #(
		.INIT('h6996)
	) name15951 (
		_w15969_,
		_w15976_,
		_w15977_,
		_w15984_,
		_w15985_
	);
	LUT4 #(
		.INIT('he0fe)
	) name15952 (
		_w15885_,
		_w15887_,
		_w15934_,
		_w15940_,
		_w15986_
	);
	LUT3 #(
		.INIT('h82)
	) name15953 (
		_w2875_,
		_w13959_,
		_w13982_,
		_w15987_
	);
	LUT3 #(
		.INIT('h82)
	) name15954 (
		_w2986_,
		_w13960_,
		_w13979_,
		_w15988_
	);
	LUT2 #(
		.INIT('h8)
	) name15955 (
		_w2874_,
		_w13716_,
		_w15989_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15956 (
		_w2975_,
		_w13712_,
		_w13714_,
		_w13847_,
		_w15990_
	);
	LUT2 #(
		.INIT('h1)
	) name15957 (
		_w15989_,
		_w15990_,
		_w15991_
	);
	LUT2 #(
		.INIT('h4)
	) name15958 (
		_w15988_,
		_w15991_,
		_w15992_
	);
	LUT3 #(
		.INIT('h9a)
	) name15959 (
		\a[26] ,
		_w15987_,
		_w15992_,
		_w15993_
	);
	LUT3 #(
		.INIT('h69)
	) name15960 (
		_w15985_,
		_w15986_,
		_w15993_,
		_w15994_
	);
	LUT3 #(
		.INIT('h82)
	) name15961 (
		_w37_,
		_w14343_,
		_w14349_,
		_w15995_
	);
	LUT3 #(
		.INIT('h28)
	) name15962 (
		_w3262_,
		_w14344_,
		_w14347_,
		_w15996_
	);
	LUT2 #(
		.INIT('h8)
	) name15963 (
		_w3214_,
		_w14112_,
		_w15997_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15964 (
		_w3249_,
		_w14108_,
		_w14111_,
		_w14235_,
		_w15998_
	);
	LUT2 #(
		.INIT('h1)
	) name15965 (
		_w15997_,
		_w15998_,
		_w15999_
	);
	LUT2 #(
		.INIT('h4)
	) name15966 (
		_w15996_,
		_w15999_,
		_w16000_
	);
	LUT3 #(
		.INIT('h9a)
	) name15967 (
		\a[23] ,
		_w15995_,
		_w16000_,
		_w16001_
	);
	LUT3 #(
		.INIT('h96)
	) name15968 (
		_w15960_,
		_w15994_,
		_w16001_,
		_w16002_
	);
	LUT2 #(
		.INIT('h4)
	) name15969 (
		_w15959_,
		_w16002_,
		_w16003_
	);
	LUT2 #(
		.INIT('h9)
	) name15970 (
		_w15959_,
		_w16002_,
		_w16004_
	);
	LUT4 #(
		.INIT('hd400)
	) name15971 (
		_w15907_,
		_w15952_,
		_w15953_,
		_w16004_,
		_w16005_
	);
	LUT4 #(
		.INIT('h32cd)
	) name15972 (
		_w15907_,
		_w15954_,
		_w15955_,
		_w16004_,
		_w16006_
	);
	LUT2 #(
		.INIT('h8)
	) name15973 (
		_w15957_,
		_w16006_,
		_w16007_
	);
	LUT2 #(
		.INIT('h6)
	) name15974 (
		_w15957_,
		_w16006_,
		_w16008_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name15975 (
		_w37_,
		_w14343_,
		_w14348_,
		_w14349_,
		_w16009_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15976 (
		_w3214_,
		_w14108_,
		_w14111_,
		_w14235_,
		_w16010_
	);
	LUT4 #(
		.INIT('h00d7)
	) name15977 (
		_w11340_,
		_w14344_,
		_w14347_,
		_w16010_,
		_w16011_
	);
	LUT3 #(
		.INIT('h9a)
	) name15978 (
		\a[23] ,
		_w16009_,
		_w16011_,
		_w16012_
	);
	LUT3 #(
		.INIT('h8e)
	) name15979 (
		_w15985_,
		_w15986_,
		_w15993_,
		_w16013_
	);
	LUT4 #(
		.INIT('h008e)
	) name15980 (
		_w15985_,
		_w15986_,
		_w15993_,
		_w16012_,
		_w16014_
	);
	LUT4 #(
		.INIT('h7100)
	) name15981 (
		_w15985_,
		_w15986_,
		_w15993_,
		_w16012_,
		_w16015_
	);
	LUT4 #(
		.INIT('h8e71)
	) name15982 (
		_w15985_,
		_w15986_,
		_w15993_,
		_w16012_,
		_w16016_
	);
	LUT4 #(
		.INIT('h02a8)
	) name15983 (
		_w2874_,
		_w13712_,
		_w13714_,
		_w13847_,
		_w16017_
	);
	LUT4 #(
		.INIT('h007d)
	) name15984 (
		_w2975_,
		_w13960_,
		_w13979_,
		_w16017_,
		_w16018_
	);
	LUT3 #(
		.INIT('h70)
	) name15985 (
		_w2986_,
		_w14112_,
		_w16018_,
		_w16019_
	);
	LUT4 #(
		.INIT('h95aa)
	) name15986 (
		\a[26] ,
		_w2875_,
		_w14116_,
		_w16019_,
		_w16020_
	);
	LUT4 #(
		.INIT('h6f06)
	) name15987 (
		_w15969_,
		_w15976_,
		_w15977_,
		_w15984_,
		_w16021_
	);
	LUT4 #(
		.INIT('h8000)
	) name15988 (
		_w81_,
		_w834_,
		_w1342_,
		_w1401_,
		_w16022_
	);
	LUT4 #(
		.INIT('h153f)
	) name15989 (
		_w78_,
		_w56_,
		_w72_,
		_w50_,
		_w16023_
	);
	LUT3 #(
		.INIT('h1f)
	) name15990 (
		_w52_,
		_w59_,
		_w166_,
		_w16024_
	);
	LUT4 #(
		.INIT('h8000)
	) name15991 (
		_w956_,
		_w957_,
		_w16023_,
		_w16024_,
		_w16025_
	);
	LUT4 #(
		.INIT('h4000)
	) name15992 (
		_w264_,
		_w2477_,
		_w4172_,
		_w7141_,
		_w16026_
	);
	LUT3 #(
		.INIT('h80)
	) name15993 (
		_w16022_,
		_w16025_,
		_w16026_,
		_w16027_
	);
	LUT4 #(
		.INIT('h8000)
	) name15994 (
		_w13212_,
		_w13213_,
		_w14978_,
		_w14980_,
		_w16028_
	);
	LUT4 #(
		.INIT('h8000)
	) name15995 (
		_w12158_,
		_w12161_,
		_w16027_,
		_w16028_,
		_w16029_
	);
	LUT2 #(
		.INIT('h8)
	) name15996 (
		_w2421_,
		_w16029_,
		_w16030_
	);
	LUT4 #(
		.INIT('h817e)
	) name15997 (
		_w15961_,
		_w15968_,
		_w15976_,
		_w16030_,
		_w16031_
	);
	LUT4 #(
		.INIT('h2228)
	) name15998 (
		_w376_,
		_w11549_,
		_w11373_,
		_w11375_,
		_w16032_
	);
	LUT4 #(
		.INIT('h007d)
	) name15999 (
		_w2407_,
		_w13062_,
		_w13099_,
		_w16032_,
		_w16033_
	);
	LUT3 #(
		.INIT('h70)
	) name16000 (
		_w2527_,
		_w13247_,
		_w16033_,
		_w16034_
	);
	LUT3 #(
		.INIT('h70)
	) name16001 (
		_w377_,
		_w13576_,
		_w16034_,
		_w16035_
	);
	LUT3 #(
		.INIT('h96)
	) name16002 (
		_w16021_,
		_w16031_,
		_w16035_,
		_w16036_
	);
	LUT4 #(
		.INIT('h02a8)
	) name16003 (
		_w2549_,
		_w13243_,
		_w13245_,
		_w13285_,
		_w16037_
	);
	LUT4 #(
		.INIT('h007d)
	) name16004 (
		_w2617_,
		_w13293_,
		_w13322_,
		_w16037_,
		_w16038_
	);
	LUT3 #(
		.INIT('h70)
	) name16005 (
		_w2854_,
		_w13716_,
		_w16038_,
		_w16039_
	);
	LUT4 #(
		.INIT('h95aa)
	) name16006 (
		\a[29] ,
		_w2550_,
		_w13720_,
		_w16039_,
		_w16040_
	);
	LUT4 #(
		.INIT('h0096)
	) name16007 (
		_w16021_,
		_w16031_,
		_w16035_,
		_w16040_,
		_w16041_
	);
	LUT4 #(
		.INIT('h6900)
	) name16008 (
		_w16021_,
		_w16031_,
		_w16035_,
		_w16040_,
		_w16042_
	);
	LUT4 #(
		.INIT('h9669)
	) name16009 (
		_w16021_,
		_w16031_,
		_w16035_,
		_w16040_,
		_w16043_
	);
	LUT2 #(
		.INIT('h9)
	) name16010 (
		_w16020_,
		_w16043_,
		_w16044_
	);
	LUT2 #(
		.INIT('h6)
	) name16011 (
		_w16016_,
		_w16044_,
		_w16045_
	);
	LUT3 #(
		.INIT('h4d)
	) name16012 (
		_w15960_,
		_w15994_,
		_w16001_,
		_w16046_
	);
	LUT2 #(
		.INIT('h1)
	) name16013 (
		_w16045_,
		_w16046_,
		_w16047_
	);
	LUT2 #(
		.INIT('h8)
	) name16014 (
		_w16045_,
		_w16046_,
		_w16048_
	);
	LUT2 #(
		.INIT('h6)
	) name16015 (
		_w16045_,
		_w16046_,
		_w16049_
	);
	LUT3 #(
		.INIT('h1e)
	) name16016 (
		_w16003_,
		_w16005_,
		_w16049_,
		_w16050_
	);
	LUT2 #(
		.INIT('h6)
	) name16017 (
		_w16007_,
		_w16050_,
		_w16051_
	);
	LUT4 #(
		.INIT('h00f1)
	) name16018 (
		_w16003_,
		_w16005_,
		_w16047_,
		_w16048_,
		_w16052_
	);
	LUT4 #(
		.INIT('h02a8)
	) name16019 (
		_w2875_,
		_w14113_,
		_w14115_,
		_w14238_,
		_w16053_
	);
	LUT4 #(
		.INIT('h02a8)
	) name16020 (
		_w2986_,
		_w14108_,
		_w14111_,
		_w14235_,
		_w16054_
	);
	LUT3 #(
		.INIT('h82)
	) name16021 (
		_w2874_,
		_w13960_,
		_w13979_,
		_w16055_
	);
	LUT3 #(
		.INIT('h07)
	) name16022 (
		_w2975_,
		_w14112_,
		_w16055_,
		_w16056_
	);
	LUT2 #(
		.INIT('h4)
	) name16023 (
		_w16054_,
		_w16056_,
		_w16057_
	);
	LUT3 #(
		.INIT('h9a)
	) name16024 (
		\a[26] ,
		_w16053_,
		_w16057_,
		_w16058_
	);
	LUT4 #(
		.INIT('h004d)
	) name16025 (
		_w16020_,
		_w16036_,
		_w16040_,
		_w16058_,
		_w16059_
	);
	LUT4 #(
		.INIT('hb200)
	) name16026 (
		_w16020_,
		_w16036_,
		_w16040_,
		_w16058_,
		_w16060_
	);
	LUT4 #(
		.INIT('hcd32)
	) name16027 (
		_w16020_,
		_w16041_,
		_w16042_,
		_w16058_,
		_w16061_
	);
	LUT3 #(
		.INIT('hb2)
	) name16028 (
		_w16021_,
		_w16031_,
		_w16035_,
		_w16062_
	);
	LUT4 #(
		.INIT('h80fe)
	) name16029 (
		_w15961_,
		_w15968_,
		_w15976_,
		_w16030_,
		_w16063_
	);
	LUT4 #(
		.INIT('h5665)
	) name16030 (
		\a[23] ,
		_w13073_,
		_w14344_,
		_w14347_,
		_w16064_
	);
	LUT3 #(
		.INIT('h57)
	) name16031 (
		_w110_,
		_w158_,
		_w259_,
		_w16065_
	);
	LUT3 #(
		.INIT('h80)
	) name16032 (
		_w66_,
		_w163_,
		_w16065_,
		_w16066_
	);
	LUT3 #(
		.INIT('h80)
	) name16033 (
		_w480_,
		_w857_,
		_w3439_,
		_w16067_
	);
	LUT4 #(
		.INIT('h8000)
	) name16034 (
		_w3349_,
		_w8253_,
		_w16067_,
		_w16066_,
		_w16068_
	);
	LUT3 #(
		.INIT('h80)
	) name16035 (
		_w234_,
		_w405_,
		_w16068_,
		_w16069_
	);
	LUT4 #(
		.INIT('h8000)
	) name16036 (
		_w2394_,
		_w2421_,
		_w16029_,
		_w16069_,
		_w16070_
	);
	LUT4 #(
		.INIT('h153f)
	) name16037 (
		_w2394_,
		_w2421_,
		_w16029_,
		_w16069_,
		_w16071_
	);
	LUT4 #(
		.INIT('h6ac0)
	) name16038 (
		_w2394_,
		_w2421_,
		_w16029_,
		_w16069_,
		_w16072_
	);
	LUT2 #(
		.INIT('h6)
	) name16039 (
		_w16064_,
		_w16072_,
		_w16073_
	);
	LUT4 #(
		.INIT('h02a8)
	) name16040 (
		_w377_,
		_w13288_,
		_w13290_,
		_w13291_,
		_w16074_
	);
	LUT4 #(
		.INIT('h02a8)
	) name16041 (
		_w2527_,
		_w13243_,
		_w13245_,
		_w13285_,
		_w16075_
	);
	LUT3 #(
		.INIT('h82)
	) name16042 (
		_w376_,
		_w13062_,
		_w13099_,
		_w16076_
	);
	LUT3 #(
		.INIT('h07)
	) name16043 (
		_w2407_,
		_w13247_,
		_w16076_,
		_w16077_
	);
	LUT2 #(
		.INIT('h4)
	) name16044 (
		_w16075_,
		_w16077_,
		_w16078_
	);
	LUT2 #(
		.INIT('h4)
	) name16045 (
		_w16074_,
		_w16078_,
		_w16079_
	);
	LUT3 #(
		.INIT('h96)
	) name16046 (
		_w16063_,
		_w16073_,
		_w16079_,
		_w16080_
	);
	LUT4 #(
		.INIT('h02a8)
	) name16047 (
		_w2550_,
		_w13717_,
		_w13719_,
		_w13850_,
		_w16081_
	);
	LUT4 #(
		.INIT('h02a8)
	) name16048 (
		_w2854_,
		_w13712_,
		_w13714_,
		_w13847_,
		_w16082_
	);
	LUT3 #(
		.INIT('h82)
	) name16049 (
		_w2549_,
		_w13293_,
		_w13322_,
		_w16083_
	);
	LUT3 #(
		.INIT('h07)
	) name16050 (
		_w2617_,
		_w13716_,
		_w16083_,
		_w16084_
	);
	LUT2 #(
		.INIT('h4)
	) name16051 (
		_w16082_,
		_w16084_,
		_w16085_
	);
	LUT3 #(
		.INIT('h9a)
	) name16052 (
		\a[29] ,
		_w16081_,
		_w16085_,
		_w16086_
	);
	LUT3 #(
		.INIT('h96)
	) name16053 (
		_w16062_,
		_w16080_,
		_w16086_,
		_w16087_
	);
	LUT2 #(
		.INIT('h6)
	) name16054 (
		_w16061_,
		_w16087_,
		_w16088_
	);
	LUT3 #(
		.INIT('h32)
	) name16055 (
		_w16014_,
		_w16015_,
		_w16044_,
		_w16089_
	);
	LUT4 #(
		.INIT('hd400)
	) name16056 (
		_w16012_,
		_w16013_,
		_w16044_,
		_w16088_,
		_w16090_
	);
	LUT4 #(
		.INIT('h002b)
	) name16057 (
		_w16012_,
		_w16013_,
		_w16044_,
		_w16088_,
		_w16091_
	);
	LUT4 #(
		.INIT('hcd32)
	) name16058 (
		_w16014_,
		_w16015_,
		_w16044_,
		_w16088_,
		_w16092_
	);
	LUT4 #(
		.INIT('h8008)
	) name16059 (
		_w16007_,
		_w16050_,
		_w16052_,
		_w16092_,
		_w16093_
	);
	LUT4 #(
		.INIT('h7887)
	) name16060 (
		_w16007_,
		_w16050_,
		_w16052_,
		_w16092_,
		_w16094_
	);
	LUT3 #(
		.INIT('h45)
	) name16061 (
		_w16059_,
		_w16060_,
		_w16087_,
		_w16095_
	);
	LUT3 #(
		.INIT('h0d)
	) name16062 (
		_w16064_,
		_w16070_,
		_w16071_,
		_w16096_
	);
	LUT3 #(
		.INIT('h80)
	) name16063 (
		_w1519_,
		_w1703_,
		_w2822_,
		_w16097_
	);
	LUT3 #(
		.INIT('h80)
	) name16064 (
		_w4203_,
		_w7835_,
		_w16097_,
		_w16098_
	);
	LUT4 #(
		.INIT('h0777)
	) name16065 (
		_w122_,
		_w52_,
		_w56_,
		_w236_,
		_w16099_
	);
	LUT2 #(
		.INIT('h8)
	) name16066 (
		_w254_,
		_w16099_,
		_w16100_
	);
	LUT4 #(
		.INIT('h8000)
	) name16067 (
		_w676_,
		_w790_,
		_w935_,
		_w1374_,
		_w16101_
	);
	LUT4 #(
		.INIT('h8000)
	) name16068 (
		_w208_,
		_w217_,
		_w16100_,
		_w16101_,
		_w16102_
	);
	LUT3 #(
		.INIT('h80)
	) name16069 (
		_w548_,
		_w16098_,
		_w16102_,
		_w16103_
	);
	LUT3 #(
		.INIT('h80)
	) name16070 (
		_w8260_,
		_w13302_,
		_w16103_,
		_w16104_
	);
	LUT4 #(
		.INIT('h0df2)
	) name16071 (
		_w16064_,
		_w16070_,
		_w16071_,
		_w16104_,
		_w16105_
	);
	LUT3 #(
		.INIT('h82)
	) name16072 (
		_w377_,
		_w13292_,
		_w13325_,
		_w16106_
	);
	LUT3 #(
		.INIT('h82)
	) name16073 (
		_w2527_,
		_w13293_,
		_w13322_,
		_w16107_
	);
	LUT2 #(
		.INIT('h8)
	) name16074 (
		_w376_,
		_w13247_,
		_w16108_
	);
	LUT4 #(
		.INIT('h02a8)
	) name16075 (
		_w2407_,
		_w13243_,
		_w13245_,
		_w13285_,
		_w16109_
	);
	LUT2 #(
		.INIT('h1)
	) name16076 (
		_w16108_,
		_w16109_,
		_w16110_
	);
	LUT2 #(
		.INIT('h4)
	) name16077 (
		_w16107_,
		_w16110_,
		_w16111_
	);
	LUT2 #(
		.INIT('h4)
	) name16078 (
		_w16106_,
		_w16111_,
		_w16112_
	);
	LUT2 #(
		.INIT('h9)
	) name16079 (
		_w16105_,
		_w16112_,
		_w16113_
	);
	LUT3 #(
		.INIT('h4d)
	) name16080 (
		_w16063_,
		_w16073_,
		_w16079_,
		_w16114_
	);
	LUT4 #(
		.INIT('h00b2)
	) name16081 (
		_w16063_,
		_w16073_,
		_w16079_,
		_w16113_,
		_w16115_
	);
	LUT4 #(
		.INIT('h4d00)
	) name16082 (
		_w16063_,
		_w16073_,
		_w16079_,
		_w16113_,
		_w16116_
	);
	LUT4 #(
		.INIT('hb24d)
	) name16083 (
		_w16063_,
		_w16073_,
		_w16079_,
		_w16113_,
		_w16117_
	);
	LUT3 #(
		.INIT('h82)
	) name16084 (
		_w2550_,
		_w13959_,
		_w13982_,
		_w16118_
	);
	LUT3 #(
		.INIT('h82)
	) name16085 (
		_w2854_,
		_w13960_,
		_w13979_,
		_w16119_
	);
	LUT2 #(
		.INIT('h8)
	) name16086 (
		_w2549_,
		_w13716_,
		_w16120_
	);
	LUT4 #(
		.INIT('h02a8)
	) name16087 (
		_w2617_,
		_w13712_,
		_w13714_,
		_w13847_,
		_w16121_
	);
	LUT2 #(
		.INIT('h1)
	) name16088 (
		_w16120_,
		_w16121_,
		_w16122_
	);
	LUT2 #(
		.INIT('h4)
	) name16089 (
		_w16119_,
		_w16122_,
		_w16123_
	);
	LUT3 #(
		.INIT('h9a)
	) name16090 (
		\a[29] ,
		_w16118_,
		_w16123_,
		_w16124_
	);
	LUT2 #(
		.INIT('h9)
	) name16091 (
		_w16117_,
		_w16124_,
		_w16125_
	);
	LUT3 #(
		.INIT('h4d)
	) name16092 (
		_w16062_,
		_w16080_,
		_w16086_,
		_w16126_
	);
	LUT3 #(
		.INIT('h82)
	) name16093 (
		_w2875_,
		_w14343_,
		_w14349_,
		_w16127_
	);
	LUT3 #(
		.INIT('h28)
	) name16094 (
		_w2986_,
		_w14344_,
		_w14347_,
		_w16128_
	);
	LUT2 #(
		.INIT('h8)
	) name16095 (
		_w2874_,
		_w14112_,
		_w16129_
	);
	LUT4 #(
		.INIT('h02a8)
	) name16096 (
		_w2975_,
		_w14108_,
		_w14111_,
		_w14235_,
		_w16130_
	);
	LUT2 #(
		.INIT('h1)
	) name16097 (
		_w16129_,
		_w16130_,
		_w16131_
	);
	LUT2 #(
		.INIT('h4)
	) name16098 (
		_w16128_,
		_w16131_,
		_w16132_
	);
	LUT3 #(
		.INIT('h9a)
	) name16099 (
		\a[26] ,
		_w16127_,
		_w16132_,
		_w16133_
	);
	LUT3 #(
		.INIT('h69)
	) name16100 (
		_w16125_,
		_w16126_,
		_w16133_,
		_w16134_
	);
	LUT2 #(
		.INIT('h4)
	) name16101 (
		_w16095_,
		_w16134_,
		_w16135_
	);
	LUT2 #(
		.INIT('h9)
	) name16102 (
		_w16095_,
		_w16134_,
		_w16136_
	);
	LUT4 #(
		.INIT('hd400)
	) name16103 (
		_w16052_,
		_w16088_,
		_w16089_,
		_w16136_,
		_w16137_
	);
	LUT4 #(
		.INIT('h32cd)
	) name16104 (
		_w16052_,
		_w16090_,
		_w16091_,
		_w16136_,
		_w16138_
	);
	LUT2 #(
		.INIT('h8)
	) name16105 (
		_w16093_,
		_w16138_,
		_w16139_
	);
	LUT2 #(
		.INIT('h6)
	) name16106 (
		_w16093_,
		_w16138_,
		_w16140_
	);
	LUT4 #(
		.INIT('h8000)
	) name16107 (
		_w49_,
		_w63_,
		_w71_,
		_w327_,
		_w16141_
	);
	LUT4 #(
		.INIT('h8000)
	) name16108 (
		_w200_,
		_w307_,
		_w174_,
		_w373_,
		_w16142_
	);
	LUT3 #(
		.INIT('h80)
	) name16109 (
		_w13302_,
		_w16141_,
		_w16142_,
		_w16143_
	);
	LUT4 #(
		.INIT('h817e)
	) name16110 (
		_w16096_,
		_w16104_,
		_w16112_,
		_w16143_,
		_w16144_
	);
	LUT4 #(
		.INIT('h02a8)
	) name16111 (
		_w376_,
		_w13243_,
		_w13245_,
		_w13285_,
		_w16145_
	);
	LUT4 #(
		.INIT('h007d)
	) name16112 (
		_w2407_,
		_w13293_,
		_w13322_,
		_w16145_,
		_w16146_
	);
	LUT3 #(
		.INIT('h70)
	) name16113 (
		_w2527_,
		_w13716_,
		_w16146_,
		_w16147_
	);
	LUT3 #(
		.INIT('h70)
	) name16114 (
		_w377_,
		_w13720_,
		_w16147_,
		_w16148_
	);
	LUT2 #(
		.INIT('h2)
	) name16115 (
		_w16144_,
		_w16148_,
		_w16149_
	);
	LUT2 #(
		.INIT('h9)
	) name16116 (
		_w16144_,
		_w16148_,
		_w16150_
	);
	LUT4 #(
		.INIT('h8e00)
	) name16117 (
		_w16113_,
		_w16114_,
		_w16124_,
		_w16150_,
		_w16151_
	);
	LUT4 #(
		.INIT('h32cd)
	) name16118 (
		_w16115_,
		_w16116_,
		_w16124_,
		_w16150_,
		_w16152_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name16119 (
		_w2875_,
		_w14343_,
		_w14348_,
		_w14349_,
		_w16153_
	);
	LUT4 #(
		.INIT('h02a8)
	) name16120 (
		_w2874_,
		_w14108_,
		_w14111_,
		_w14235_,
		_w16154_
	);
	LUT4 #(
		.INIT('h00eb)
	) name16121 (
		_w13205_,
		_w14344_,
		_w14347_,
		_w16154_,
		_w16155_
	);
	LUT4 #(
		.INIT('h02a8)
	) name16122 (
		_w2549_,
		_w13712_,
		_w13714_,
		_w13847_,
		_w16156_
	);
	LUT4 #(
		.INIT('h007d)
	) name16123 (
		_w2617_,
		_w13960_,
		_w13979_,
		_w16156_,
		_w16157_
	);
	LUT3 #(
		.INIT('h70)
	) name16124 (
		_w2854_,
		_w14112_,
		_w16157_,
		_w16158_
	);
	LUT4 #(
		.INIT('h95aa)
	) name16125 (
		\a[29] ,
		_w2550_,
		_w14116_,
		_w16158_,
		_w16159_
	);
	LUT4 #(
		.INIT('h0065)
	) name16126 (
		\a[26] ,
		_w16153_,
		_w16155_,
		_w16159_,
		_w16160_
	);
	LUT4 #(
		.INIT('h9a00)
	) name16127 (
		\a[26] ,
		_w16153_,
		_w16155_,
		_w16159_,
		_w16161_
	);
	LUT4 #(
		.INIT('h659a)
	) name16128 (
		\a[26] ,
		_w16153_,
		_w16155_,
		_w16159_,
		_w16162_
	);
	LUT2 #(
		.INIT('h6)
	) name16129 (
		_w16152_,
		_w16162_,
		_w16163_
	);
	LUT3 #(
		.INIT('h8e)
	) name16130 (
		_w16125_,
		_w16126_,
		_w16133_,
		_w16164_
	);
	LUT2 #(
		.INIT('h8)
	) name16131 (
		_w16163_,
		_w16164_,
		_w16165_
	);
	LUT2 #(
		.INIT('h1)
	) name16132 (
		_w16163_,
		_w16164_,
		_w16166_
	);
	LUT2 #(
		.INIT('h6)
	) name16133 (
		_w16163_,
		_w16164_,
		_w16167_
	);
	LUT3 #(
		.INIT('h1e)
	) name16134 (
		_w16135_,
		_w16137_,
		_w16167_,
		_w16168_
	);
	LUT2 #(
		.INIT('h6)
	) name16135 (
		_w16139_,
		_w16168_,
		_w16169_
	);
	LUT3 #(
		.INIT('h31)
	) name16136 (
		_w16152_,
		_w16160_,
		_w16161_,
		_w16170_
	);
	LUT4 #(
		.INIT('h0f01)
	) name16137 (
		_w16135_,
		_w16137_,
		_w16165_,
		_w16166_,
		_w16171_
	);
	LUT3 #(
		.INIT('h69)
	) name16138 (
		_w16104_,
		_w16170_,
		_w16171_,
		_w16172_
	);
	LUT3 #(
		.INIT('h14)
	) name16139 (
		_w13300_,
		_w14344_,
		_w14347_,
		_w16173_
	);
	LUT4 #(
		.INIT('hb332)
	) name16140 (
		_w16096_,
		_w16104_,
		_w16112_,
		_w16143_,
		_w16174_
	);
	LUT4 #(
		.INIT('h02a8)
	) name16141 (
		_w377_,
		_w13717_,
		_w13719_,
		_w13850_,
		_w16175_
	);
	LUT4 #(
		.INIT('h02a8)
	) name16142 (
		_w2527_,
		_w13712_,
		_w13714_,
		_w13847_,
		_w16176_
	);
	LUT3 #(
		.INIT('h82)
	) name16143 (
		_w376_,
		_w13293_,
		_w13322_,
		_w16177_
	);
	LUT3 #(
		.INIT('h07)
	) name16144 (
		_w2407_,
		_w13716_,
		_w16177_,
		_w16178_
	);
	LUT2 #(
		.INIT('h4)
	) name16145 (
		_w16176_,
		_w16178_,
		_w16179_
	);
	LUT3 #(
		.INIT('h65)
	) name16146 (
		\a[26] ,
		_w16175_,
		_w16179_,
		_w16180_
	);
	LUT2 #(
		.INIT('h9)
	) name16147 (
		_w16174_,
		_w16180_,
		_w16181_
	);
	LUT4 #(
		.INIT('h9555)
	) name16148 (
		\a[29] ,
		_w121_,
		_w351_,
		_w418_,
		_w16182_
	);
	LUT4 #(
		.INIT('h02a8)
	) name16149 (
		_w2550_,
		_w14113_,
		_w14115_,
		_w14238_,
		_w16183_
	);
	LUT4 #(
		.INIT('h02a8)
	) name16150 (
		_w2854_,
		_w14108_,
		_w14111_,
		_w14235_,
		_w16184_
	);
	LUT3 #(
		.INIT('h82)
	) name16151 (
		_w2549_,
		_w13960_,
		_w13979_,
		_w16185_
	);
	LUT3 #(
		.INIT('h07)
	) name16152 (
		_w2617_,
		_w14112_,
		_w16185_,
		_w16186_
	);
	LUT2 #(
		.INIT('h4)
	) name16153 (
		_w16184_,
		_w16186_,
		_w16187_
	);
	LUT2 #(
		.INIT('h4)
	) name16154 (
		_w16183_,
		_w16187_,
		_w16188_
	);
	LUT4 #(
		.INIT('he11e)
	) name16155 (
		_w16149_,
		_w16151_,
		_w16182_,
		_w16188_,
		_w16189_
	);
	LUT2 #(
		.INIT('h9)
	) name16156 (
		_w16181_,
		_w16189_,
		_w16190_
	);
	LUT4 #(
		.INIT('h8778)
	) name16157 (
		_w16139_,
		_w16168_,
		_w16173_,
		_w16190_,
		_w16191_
	);
	LUT2 #(
		.INIT('h9)
	) name16158 (
		_w16172_,
		_w16191_,
		_w16192_
	);
	assign \result[0]  = _w13730_ ;
	assign \result[1]  = _w13861_ ;
	assign \result[2]  = _w13994_ ;
	assign \result[3]  = _w14125_ ;
	assign \result[4]  = _w14249_ ;
	assign \result[5]  = _w14361_ ;
	assign \result[6]  = _w14472_ ;
	assign \result[7]  = _w14568_ ;
	assign \result[8]  = _w14673_ ;
	assign \result[9]  = _w14756_ ;
	assign \result[10]  = _w14850_ ;
	assign \result[11]  = _w14959_ ;
	assign \result[12]  = _w15040_ ;
	assign \result[13]  = _w15135_ ;
	assign \result[14]  = _w15225_ ;
	assign \result[15]  = _w15292_ ;
	assign \result[16]  = _w15381_ ;
	assign \result[17]  = _w15465_ ;
	assign \result[18]  = _w15525_ ;
	assign \result[19]  = _w15601_ ;
	assign \result[20]  = _w15669_ ;
	assign \result[21]  = _w15727_ ;
	assign \result[22]  = _w15795_ ;
	assign \result[23]  = _w15860_ ;
	assign \result[24]  = _w15906_ ;
	assign \result[25]  = _w15958_ ;
	assign \result[26]  = _w16008_ ;
	assign \result[27]  = _w16051_ ;
	assign \result[28]  = _w16094_ ;
	assign \result[29]  = _w16140_ ;
	assign \result[30]  = _w16169_ ;
	assign \result[31]  = _w16192_ ;
endmodule;