module top( a_pad , b_pad , c_pad , d_pad , e_pad , f_pad , g_pad , h_pad , i_pad , j_pad , k_pad , l_pad );
  input a_pad ;
  input b_pad ;
  input c_pad ;
  input d_pad ;
  input e_pad ;
  input f_pad ;
  input g_pad ;
  input h_pad ;
  input i_pad ;
  input j_pad ;
  input k_pad ;
  output l_pad ;
  wire n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 ;
  assign n13 = ~g_pad & j_pad ;
  assign n12 = ~e_pad & ~j_pad ;
  assign n14 = ~i_pad & ~n12 ;
  assign n15 = ~n13 & n14 ;
  assign n17 = ~h_pad & j_pad ;
  assign n16 = ~f_pad & ~j_pad ;
  assign n18 = i_pad & ~n16 ;
  assign n19 = ~n17 & n18 ;
  assign n20 = ~n15 & ~n19 ;
  assign n21 = k_pad & ~n20 ;
  assign n23 = ~c_pad & j_pad ;
  assign n22 = ~a_pad & ~j_pad ;
  assign n24 = ~i_pad & ~n22 ;
  assign n25 = ~n23 & n24 ;
  assign n27 = ~b_pad & ~j_pad ;
  assign n26 = ~d_pad & j_pad ;
  assign n28 = i_pad & ~n26 ;
  assign n29 = ~n27 & n28 ;
  assign n30 = ~n25 & ~n29 ;
  assign n31 = ~k_pad & ~n30 ;
  assign n32 = ~n21 & ~n31 ;
  assign l_pad = ~n32 ;
endmodule
