module top (\clgen_cnt_reg[0]/NET0131 , \clgen_cnt_reg[10]/NET0131 , \clgen_cnt_reg[11]/NET0131 , \clgen_cnt_reg[12]/NET0131 , \clgen_cnt_reg[13]/NET0131 , \clgen_cnt_reg[14]/NET0131 , \clgen_cnt_reg[15]/NET0131 , \clgen_cnt_reg[1]/NET0131 , \clgen_cnt_reg[2]/NET0131 , \clgen_cnt_reg[3]/NET0131 , \clgen_cnt_reg[4]/NET0131 , \clgen_cnt_reg[5]/NET0131 , \clgen_cnt_reg[6]/NET0131 , \clgen_cnt_reg[7]/NET0131 , \clgen_cnt_reg[8]/NET0131 , \clgen_cnt_reg[9]/NET0131 , \clgen_neg_edge_reg/NET0131 , \clgen_pos_edge_reg/NET0131 , \ctrl_reg[0]/NET0131 , \ctrl_reg[10]/NET0131 , \ctrl_reg[11]/NET0131 , \ctrl_reg[12]/NET0131 , \ctrl_reg[13]/NET0131 , \ctrl_reg[1]/NET0131 , \ctrl_reg[2]/NET0131 , \ctrl_reg[3]/NET0131 , \ctrl_reg[4]/NET0131 , \ctrl_reg[5]/NET0131 , \ctrl_reg[6]/NET0131 , \ctrl_reg[7]/NET0131 , \ctrl_reg[8]/NET0131 , \ctrl_reg[9]/NET0131 , \divider_reg[0]/NET0131 , \divider_reg[10]/NET0131 , \divider_reg[11]/NET0131 , \divider_reg[12]/NET0131 , \divider_reg[13]/NET0131 , \divider_reg[14]/NET0131 , \divider_reg[15]/NET0131 , \divider_reg[1]/NET0131 , \divider_reg[2]/NET0131 , \divider_reg[3]/NET0131 , \divider_reg[4]/NET0131 , \divider_reg[5]/NET0131 , \divider_reg[6]/NET0131 , \divider_reg[7]/NET0131 , \divider_reg[8]/NET0131 , \divider_reg[9]/NET0131 , miso_pad_i_pad, mosi_pad_o_pad, sclk_pad_o_pad, \shift_cnt_reg[0]/NET0131 , \shift_cnt_reg[1]/NET0131 , \shift_cnt_reg[2]/NET0131 , \shift_cnt_reg[3]/NET0131 , \shift_cnt_reg[4]/NET0131 , \shift_cnt_reg[5]/NET0131 , \shift_cnt_reg[6]/NET0131 , \shift_cnt_reg[7]/NET0131 , \shift_data_reg[0]/NET0131 , \shift_data_reg[100]/NET0131 , \shift_data_reg[101]/NET0131 , \shift_data_reg[102]/NET0131 , \shift_data_reg[103]/NET0131 , \shift_data_reg[104]/NET0131 , \shift_data_reg[105]/NET0131 , \shift_data_reg[106]/NET0131 , \shift_data_reg[107]/NET0131 , \shift_data_reg[108]/NET0131 , \shift_data_reg[109]/NET0131 , \shift_data_reg[10]/NET0131 , \shift_data_reg[110]/NET0131 , \shift_data_reg[111]/NET0131 , \shift_data_reg[112]/NET0131 , \shift_data_reg[113]/NET0131 , \shift_data_reg[114]/NET0131 , \shift_data_reg[115]/NET0131 , \shift_data_reg[116]/NET0131 , \shift_data_reg[117]/NET0131 , \shift_data_reg[118]/NET0131 , \shift_data_reg[119]/NET0131 , \shift_data_reg[11]/NET0131 , \shift_data_reg[120]/NET0131 , \shift_data_reg[121]/NET0131 , \shift_data_reg[122]/NET0131 , \shift_data_reg[123]/NET0131 , \shift_data_reg[124]/NET0131 , \shift_data_reg[125]/NET0131 , \shift_data_reg[126]/NET0131 , \shift_data_reg[127]/NET0131 , \shift_data_reg[12]/NET0131 , \shift_data_reg[13]/NET0131 , \shift_data_reg[14]/NET0131 , \shift_data_reg[15]/NET0131 , \shift_data_reg[16]/NET0131 , \shift_data_reg[17]/NET0131 , \shift_data_reg[18]/NET0131 , \shift_data_reg[19]/NET0131 , \shift_data_reg[1]/NET0131 , \shift_data_reg[20]/NET0131 , \shift_data_reg[21]/NET0131 , \shift_data_reg[22]/NET0131 , \shift_data_reg[23]/NET0131 , \shift_data_reg[24]/NET0131 , \shift_data_reg[25]/NET0131 , \shift_data_reg[26]/NET0131 , \shift_data_reg[27]/NET0131 , \shift_data_reg[28]/NET0131 , \shift_data_reg[29]/NET0131 , \shift_data_reg[2]/NET0131 , \shift_data_reg[30]/NET0131 , \shift_data_reg[31]/NET0131 , \shift_data_reg[32]/NET0131 , \shift_data_reg[33]/NET0131 , \shift_data_reg[34]/NET0131 , \shift_data_reg[35]/NET0131 , \shift_data_reg[36]/NET0131 , \shift_data_reg[37]/NET0131 , \shift_data_reg[38]/NET0131 , \shift_data_reg[39]/NET0131 , \shift_data_reg[3]/NET0131 , \shift_data_reg[40]/NET0131 , \shift_data_reg[41]/NET0131 , \shift_data_reg[42]/NET0131 , \shift_data_reg[43]/NET0131 , \shift_data_reg[44]/NET0131 , \shift_data_reg[45]/NET0131 , \shift_data_reg[46]/NET0131 , \shift_data_reg[47]/NET0131 , \shift_data_reg[48]/NET0131 , \shift_data_reg[49]/NET0131 , \shift_data_reg[4]/NET0131 , \shift_data_reg[50]/NET0131 , \shift_data_reg[51]/NET0131 , \shift_data_reg[52]/NET0131 , \shift_data_reg[53]/NET0131 , \shift_data_reg[54]/NET0131 , \shift_data_reg[55]/NET0131 , \shift_data_reg[56]/NET0131 , \shift_data_reg[57]/NET0131 , \shift_data_reg[58]/NET0131 , \shift_data_reg[59]/NET0131 , \shift_data_reg[5]/NET0131 , \shift_data_reg[60]/NET0131 , \shift_data_reg[61]/NET0131 , \shift_data_reg[62]/NET0131 , \shift_data_reg[63]/NET0131 , \shift_data_reg[64]/NET0131 , \shift_data_reg[65]/NET0131 , \shift_data_reg[66]/NET0131 , \shift_data_reg[67]/NET0131 , \shift_data_reg[68]/NET0131 , \shift_data_reg[69]/NET0131 , \shift_data_reg[6]/NET0131 , \shift_data_reg[70]/NET0131 , \shift_data_reg[71]/NET0131 , \shift_data_reg[72]/NET0131 , \shift_data_reg[73]/NET0131 , \shift_data_reg[74]/NET0131 , \shift_data_reg[75]/NET0131 , \shift_data_reg[76]/NET0131 , \shift_data_reg[77]/NET0131 , \shift_data_reg[78]/NET0131 , \shift_data_reg[79]/NET0131 , \shift_data_reg[7]/NET0131 , \shift_data_reg[80]/NET0131 , \shift_data_reg[81]/NET0131 , \shift_data_reg[82]/NET0131 , \shift_data_reg[83]/NET0131 , \shift_data_reg[84]/NET0131 , \shift_data_reg[85]/NET0131 , \shift_data_reg[86]/NET0131 , \shift_data_reg[87]/NET0131 , \shift_data_reg[88]/NET0131 , \shift_data_reg[89]/NET0131 , \shift_data_reg[8]/NET0131 , \shift_data_reg[90]/NET0131 , \shift_data_reg[91]/NET0131 , \shift_data_reg[92]/NET0131 , \shift_data_reg[93]/NET0131 , \shift_data_reg[94]/NET0131 , \shift_data_reg[95]/NET0131 , \shift_data_reg[96]/NET0131 , \shift_data_reg[97]/NET0131 , \shift_data_reg[98]/NET0131 , \shift_data_reg[99]/NET0131 , \shift_data_reg[9]/NET0131 , \shift_tip_reg/NET0131 , \ss_reg[0]/NET0131 , \ss_reg[1]/NET0131 , \ss_reg[2]/NET0131 , \ss_reg[3]/NET0131 , \ss_reg[4]/NET0131 , \ss_reg[5]/NET0131 , \ss_reg[6]/NET0131 , \ss_reg[7]/NET0131 , wb_ack_o_pad, \wb_adr_i[2]_pad , \wb_adr_i[3]_pad , \wb_adr_i[4]_pad , wb_cyc_i_pad, \wb_dat_i[0]_pad , \wb_dat_i[10]_pad , \wb_dat_i[11]_pad , \wb_dat_i[12]_pad , \wb_dat_i[13]_pad , \wb_dat_i[14]_pad , \wb_dat_i[15]_pad , \wb_dat_i[16]_pad , \wb_dat_i[17]_pad , \wb_dat_i[18]_pad , \wb_dat_i[19]_pad , \wb_dat_i[1]_pad , \wb_dat_i[20]_pad , \wb_dat_i[21]_pad , \wb_dat_i[22]_pad , \wb_dat_i[23]_pad , \wb_dat_i[24]_pad , \wb_dat_i[25]_pad , \wb_dat_i[26]_pad , \wb_dat_i[27]_pad , \wb_dat_i[28]_pad , \wb_dat_i[29]_pad , \wb_dat_i[2]_pad , \wb_dat_i[30]_pad , \wb_dat_i[31]_pad , \wb_dat_i[3]_pad , \wb_dat_i[4]_pad , \wb_dat_i[5]_pad , \wb_dat_i[6]_pad , \wb_dat_i[7]_pad , \wb_dat_i[8]_pad , \wb_dat_i[9]_pad , wb_int_o_pad, \wb_sel_i[0]_pad , \wb_sel_i[1]_pad , \wb_sel_i[2]_pad , \wb_sel_i[3]_pad , wb_stb_i_pad, wb_we_i_pad, \_al_n1 , \g10384/_0_ , \g10421/_0_ , \g10487/_0_ , \g10622/_0_ , \g10625/_0_ , \g10631/_3_ , \g10641/_0_ , \g10677/_3_ , \g10695/_0_ , \g10699/_3_ , \g10796/_0_ , \g10814/_00_ , \g10815/_0_ , \g10819/_0_ , \g10821/_0_ , \g10824/_3_ , \g10858/_0_ , \g11042/_00_ , \g11067/_0_ , \g11071/_00_ , \g11074/_0_ , \g11075/_0_ , \g11076/_0_ , \g11077/_0_ , \g11078/_0_ , \g11079/_0_ , \g11080/_0_ , \g11149/_0_ , \g11151/_0_ , \g11190/_00_ , \g11297/_0_ , \g11298/_0_ , \g11300/_0_ , \g11301/_0_ , \g11303/_0_ , \g11346/_0_ , \g11347/_0_ , \g11348/_0_ , \g11358/_0_ , \g11359/_0_ , \g11360/_0_ , \g11361/_0_ , \g11362/_0_ , \g11363/_0_ , \g11470/_0_ , \g11499/_0_ , \g11501/_0_ , \g11502/_0_ , \g11503/_0_ , \g11504/_0_ , \g11505/_0_ , \g11506/_0_ , \g11507/_0_ , \g11508/_0_ , \g11509/_0_ , \g11510/_0_ , \g11511/_0_ , \g11512/_0_ , \g11513/_0_ , \g11514/_0_ , \g11515/_0_ , \g11516/_0_ , \g11517/_0_ , \g11519/_0_ , \g11520/_0_ , \g11521/_0_ , \g11522/_0_ , \g11523/_0_ , \g11524/_0_ , \g11525/_0_ , \g11526/_0_ , \g11527/_0_ , \g11528/_0_ , \g11529/_0_ , \g11530/_0_ , \g11531/_0_ , \g11532/_0_ , \g11533/_0_ , \g11534/_0_ , \g11535/_0_ , \g11536/_0_ , \g11537/_0_ , \g11538/_0_ , \g11539/_0_ , \g11655/_0_ , \g11658/_0_ , \g11659/_0_ , \g11661/_0_ , \g11662/_0_ , \g11680/_0_ , \g11723/_0_ , \g11726/_0_ , \g11730/_0_ , \g11739/_0_ , \g11750/_0_ , \g11759/_0_ , \g11760/_0_ , \g11761/_0_ , \g11764/_0_ , \g11765/_0_ , \g12212/_0_ , \g13497/_0_ , \g13884/_0_ , \g13982/_0_ , \g13999/_0_ , \g9305/_0_ , \g9306/_0_ , \g9307/_0_ , \g9308/_0_ , \g9309/_0_ , \g9310/_0_ , \g9346/_0_ , \g9347/_0_ , \g9348/_0_ , \g9349/_0_ , \g9350/_0_ , \g9351/_0_ , \g9352/_0_ , \g9353/_0_ , \g9354/_0_ , \g9355/_0_ , \g9356/_0_ , \g9357/_0_ , \g9358/_0_ , \g9359/_0_ , \g9360/_0_ , \g9361/_0_ , \g9362/_0_ , \g9363/_0_ , \g9364/_0_ , \g9365/_0_ , \g9366/_0_ , \g9367/_0_ , \g9368/_0_ , \g9369/_0_ , \g9370/_0_ , \g9371/_0_ , \g9372/_0_ , \g9373/_0_ , \g9374/_0_ , \g9375/_0_ , \g9380/_0_ , \g9381/_0_ , \g9382/_0_ , \g9383/_0_ , \g9384/_0_ , \g9385/_0_ , \g9386/_0_ , \g9387/_0_ , \g9388/_0_ , \g9389/_0_ , \g9390/_0_ , \g9391/_0_ , \g9392/_0_ , \g9393/_0_ , \g9394/_0_ , \g9395/_0_ , \g9396/_0_ , \g9397/_0_ , \g9398/_0_ , \g9399/_0_ , \g9400/_0_ , \g9401/_0_ , \g9402/_0_ , \g9403/_0_ , \g9404/_0_ , \g9405/_0_ , \g9406/_0_ , \g9407/_0_ , \g9408/_0_ , \g9409/_0_ , \g9410/_0_ , \g9411/_0_ , \g9439/_0_ , \g9440/_0_ , \g9441/_0_ , \g9442/_0_ , \g9443/_0_ , \g9444/_0_ , \g9445/_0_ , \g9446/_0_ , \g9447/_0_ , \g9448/_0_ , \g9449/_0_ , \g9450/_0_ , \g9451/_0_ , \g9452/_0_ , \g9453/_0_ , \g9454/_0_ , \g9455/_0_ , \g9456/_0_ , \g9457/_0_ , \g9458/_0_ , \g9459/_0_ , \g9461/_0_ , \g9462/_0_ , \g9463/_0_ , \g9464/_0_ , \g9465/_0_ , \g9466/_0_ , \g9529/_0_ , \g9530/_0_ , \g9531/_0_ , \g9532/_0_ , \g9535/_0_ , \g9542/_0_ , \g9543/_0_ , \g9546/_0_ , \g9547/_0_ , \g9548/_0_ , \g9549/_0_ , \g9550/_0_ , \g9551/_0_ , \g9552/_0_ , \g9553/_0_ , \g9559/_0_ , \g9568/_0_ , \g9571/_0_ , \g9573/_0_ , \g9583/_0_ , \g9589/_0_ , \g9590/_0_ , \g9591/_0_ , \g9592/_0_ , \g9593/_0_ , \g9594/_0_ , \g9595/_0_ , \g9596/_0_ , \g9597/_0_ , \ss_pad_o[0]_pad , \ss_pad_o[1]_pad , \ss_pad_o[2]_pad , \ss_pad_o[3]_pad , \ss_pad_o[4]_pad , \ss_pad_o[5]_pad , \ss_pad_o[6]_pad , \ss_pad_o[7]_pad , wb_err_o_pad);
	input \clgen_cnt_reg[0]/NET0131  ;
	input \clgen_cnt_reg[10]/NET0131  ;
	input \clgen_cnt_reg[11]/NET0131  ;
	input \clgen_cnt_reg[12]/NET0131  ;
	input \clgen_cnt_reg[13]/NET0131  ;
	input \clgen_cnt_reg[14]/NET0131  ;
	input \clgen_cnt_reg[15]/NET0131  ;
	input \clgen_cnt_reg[1]/NET0131  ;
	input \clgen_cnt_reg[2]/NET0131  ;
	input \clgen_cnt_reg[3]/NET0131  ;
	input \clgen_cnt_reg[4]/NET0131  ;
	input \clgen_cnt_reg[5]/NET0131  ;
	input \clgen_cnt_reg[6]/NET0131  ;
	input \clgen_cnt_reg[7]/NET0131  ;
	input \clgen_cnt_reg[8]/NET0131  ;
	input \clgen_cnt_reg[9]/NET0131  ;
	input \clgen_neg_edge_reg/NET0131  ;
	input \clgen_pos_edge_reg/NET0131  ;
	input \ctrl_reg[0]/NET0131  ;
	input \ctrl_reg[10]/NET0131  ;
	input \ctrl_reg[11]/NET0131  ;
	input \ctrl_reg[12]/NET0131  ;
	input \ctrl_reg[13]/NET0131  ;
	input \ctrl_reg[1]/NET0131  ;
	input \ctrl_reg[2]/NET0131  ;
	input \ctrl_reg[3]/NET0131  ;
	input \ctrl_reg[4]/NET0131  ;
	input \ctrl_reg[5]/NET0131  ;
	input \ctrl_reg[6]/NET0131  ;
	input \ctrl_reg[7]/NET0131  ;
	input \ctrl_reg[8]/NET0131  ;
	input \ctrl_reg[9]/NET0131  ;
	input \divider_reg[0]/NET0131  ;
	input \divider_reg[10]/NET0131  ;
	input \divider_reg[11]/NET0131  ;
	input \divider_reg[12]/NET0131  ;
	input \divider_reg[13]/NET0131  ;
	input \divider_reg[14]/NET0131  ;
	input \divider_reg[15]/NET0131  ;
	input \divider_reg[1]/NET0131  ;
	input \divider_reg[2]/NET0131  ;
	input \divider_reg[3]/NET0131  ;
	input \divider_reg[4]/NET0131  ;
	input \divider_reg[5]/NET0131  ;
	input \divider_reg[6]/NET0131  ;
	input \divider_reg[7]/NET0131  ;
	input \divider_reg[8]/NET0131  ;
	input \divider_reg[9]/NET0131  ;
	input miso_pad_i_pad ;
	input mosi_pad_o_pad ;
	input sclk_pad_o_pad ;
	input \shift_cnt_reg[0]/NET0131  ;
	input \shift_cnt_reg[1]/NET0131  ;
	input \shift_cnt_reg[2]/NET0131  ;
	input \shift_cnt_reg[3]/NET0131  ;
	input \shift_cnt_reg[4]/NET0131  ;
	input \shift_cnt_reg[5]/NET0131  ;
	input \shift_cnt_reg[6]/NET0131  ;
	input \shift_cnt_reg[7]/NET0131  ;
	input \shift_data_reg[0]/NET0131  ;
	input \shift_data_reg[100]/NET0131  ;
	input \shift_data_reg[101]/NET0131  ;
	input \shift_data_reg[102]/NET0131  ;
	input \shift_data_reg[103]/NET0131  ;
	input \shift_data_reg[104]/NET0131  ;
	input \shift_data_reg[105]/NET0131  ;
	input \shift_data_reg[106]/NET0131  ;
	input \shift_data_reg[107]/NET0131  ;
	input \shift_data_reg[108]/NET0131  ;
	input \shift_data_reg[109]/NET0131  ;
	input \shift_data_reg[10]/NET0131  ;
	input \shift_data_reg[110]/NET0131  ;
	input \shift_data_reg[111]/NET0131  ;
	input \shift_data_reg[112]/NET0131  ;
	input \shift_data_reg[113]/NET0131  ;
	input \shift_data_reg[114]/NET0131  ;
	input \shift_data_reg[115]/NET0131  ;
	input \shift_data_reg[116]/NET0131  ;
	input \shift_data_reg[117]/NET0131  ;
	input \shift_data_reg[118]/NET0131  ;
	input \shift_data_reg[119]/NET0131  ;
	input \shift_data_reg[11]/NET0131  ;
	input \shift_data_reg[120]/NET0131  ;
	input \shift_data_reg[121]/NET0131  ;
	input \shift_data_reg[122]/NET0131  ;
	input \shift_data_reg[123]/NET0131  ;
	input \shift_data_reg[124]/NET0131  ;
	input \shift_data_reg[125]/NET0131  ;
	input \shift_data_reg[126]/NET0131  ;
	input \shift_data_reg[127]/NET0131  ;
	input \shift_data_reg[12]/NET0131  ;
	input \shift_data_reg[13]/NET0131  ;
	input \shift_data_reg[14]/NET0131  ;
	input \shift_data_reg[15]/NET0131  ;
	input \shift_data_reg[16]/NET0131  ;
	input \shift_data_reg[17]/NET0131  ;
	input \shift_data_reg[18]/NET0131  ;
	input \shift_data_reg[19]/NET0131  ;
	input \shift_data_reg[1]/NET0131  ;
	input \shift_data_reg[20]/NET0131  ;
	input \shift_data_reg[21]/NET0131  ;
	input \shift_data_reg[22]/NET0131  ;
	input \shift_data_reg[23]/NET0131  ;
	input \shift_data_reg[24]/NET0131  ;
	input \shift_data_reg[25]/NET0131  ;
	input \shift_data_reg[26]/NET0131  ;
	input \shift_data_reg[27]/NET0131  ;
	input \shift_data_reg[28]/NET0131  ;
	input \shift_data_reg[29]/NET0131  ;
	input \shift_data_reg[2]/NET0131  ;
	input \shift_data_reg[30]/NET0131  ;
	input \shift_data_reg[31]/NET0131  ;
	input \shift_data_reg[32]/NET0131  ;
	input \shift_data_reg[33]/NET0131  ;
	input \shift_data_reg[34]/NET0131  ;
	input \shift_data_reg[35]/NET0131  ;
	input \shift_data_reg[36]/NET0131  ;
	input \shift_data_reg[37]/NET0131  ;
	input \shift_data_reg[38]/NET0131  ;
	input \shift_data_reg[39]/NET0131  ;
	input \shift_data_reg[3]/NET0131  ;
	input \shift_data_reg[40]/NET0131  ;
	input \shift_data_reg[41]/NET0131  ;
	input \shift_data_reg[42]/NET0131  ;
	input \shift_data_reg[43]/NET0131  ;
	input \shift_data_reg[44]/NET0131  ;
	input \shift_data_reg[45]/NET0131  ;
	input \shift_data_reg[46]/NET0131  ;
	input \shift_data_reg[47]/NET0131  ;
	input \shift_data_reg[48]/NET0131  ;
	input \shift_data_reg[49]/NET0131  ;
	input \shift_data_reg[4]/NET0131  ;
	input \shift_data_reg[50]/NET0131  ;
	input \shift_data_reg[51]/NET0131  ;
	input \shift_data_reg[52]/NET0131  ;
	input \shift_data_reg[53]/NET0131  ;
	input \shift_data_reg[54]/NET0131  ;
	input \shift_data_reg[55]/NET0131  ;
	input \shift_data_reg[56]/NET0131  ;
	input \shift_data_reg[57]/NET0131  ;
	input \shift_data_reg[58]/NET0131  ;
	input \shift_data_reg[59]/NET0131  ;
	input \shift_data_reg[5]/NET0131  ;
	input \shift_data_reg[60]/NET0131  ;
	input \shift_data_reg[61]/NET0131  ;
	input \shift_data_reg[62]/NET0131  ;
	input \shift_data_reg[63]/NET0131  ;
	input \shift_data_reg[64]/NET0131  ;
	input \shift_data_reg[65]/NET0131  ;
	input \shift_data_reg[66]/NET0131  ;
	input \shift_data_reg[67]/NET0131  ;
	input \shift_data_reg[68]/NET0131  ;
	input \shift_data_reg[69]/NET0131  ;
	input \shift_data_reg[6]/NET0131  ;
	input \shift_data_reg[70]/NET0131  ;
	input \shift_data_reg[71]/NET0131  ;
	input \shift_data_reg[72]/NET0131  ;
	input \shift_data_reg[73]/NET0131  ;
	input \shift_data_reg[74]/NET0131  ;
	input \shift_data_reg[75]/NET0131  ;
	input \shift_data_reg[76]/NET0131  ;
	input \shift_data_reg[77]/NET0131  ;
	input \shift_data_reg[78]/NET0131  ;
	input \shift_data_reg[79]/NET0131  ;
	input \shift_data_reg[7]/NET0131  ;
	input \shift_data_reg[80]/NET0131  ;
	input \shift_data_reg[81]/NET0131  ;
	input \shift_data_reg[82]/NET0131  ;
	input \shift_data_reg[83]/NET0131  ;
	input \shift_data_reg[84]/NET0131  ;
	input \shift_data_reg[85]/NET0131  ;
	input \shift_data_reg[86]/NET0131  ;
	input \shift_data_reg[87]/NET0131  ;
	input \shift_data_reg[88]/NET0131  ;
	input \shift_data_reg[89]/NET0131  ;
	input \shift_data_reg[8]/NET0131  ;
	input \shift_data_reg[90]/NET0131  ;
	input \shift_data_reg[91]/NET0131  ;
	input \shift_data_reg[92]/NET0131  ;
	input \shift_data_reg[93]/NET0131  ;
	input \shift_data_reg[94]/NET0131  ;
	input \shift_data_reg[95]/NET0131  ;
	input \shift_data_reg[96]/NET0131  ;
	input \shift_data_reg[97]/NET0131  ;
	input \shift_data_reg[98]/NET0131  ;
	input \shift_data_reg[99]/NET0131  ;
	input \shift_data_reg[9]/NET0131  ;
	input \shift_tip_reg/NET0131  ;
	input \ss_reg[0]/NET0131  ;
	input \ss_reg[1]/NET0131  ;
	input \ss_reg[2]/NET0131  ;
	input \ss_reg[3]/NET0131  ;
	input \ss_reg[4]/NET0131  ;
	input \ss_reg[5]/NET0131  ;
	input \ss_reg[6]/NET0131  ;
	input \ss_reg[7]/NET0131  ;
	input wb_ack_o_pad ;
	input \wb_adr_i[2]_pad  ;
	input \wb_adr_i[3]_pad  ;
	input \wb_adr_i[4]_pad  ;
	input wb_cyc_i_pad ;
	input \wb_dat_i[0]_pad  ;
	input \wb_dat_i[10]_pad  ;
	input \wb_dat_i[11]_pad  ;
	input \wb_dat_i[12]_pad  ;
	input \wb_dat_i[13]_pad  ;
	input \wb_dat_i[14]_pad  ;
	input \wb_dat_i[15]_pad  ;
	input \wb_dat_i[16]_pad  ;
	input \wb_dat_i[17]_pad  ;
	input \wb_dat_i[18]_pad  ;
	input \wb_dat_i[19]_pad  ;
	input \wb_dat_i[1]_pad  ;
	input \wb_dat_i[20]_pad  ;
	input \wb_dat_i[21]_pad  ;
	input \wb_dat_i[22]_pad  ;
	input \wb_dat_i[23]_pad  ;
	input \wb_dat_i[24]_pad  ;
	input \wb_dat_i[25]_pad  ;
	input \wb_dat_i[26]_pad  ;
	input \wb_dat_i[27]_pad  ;
	input \wb_dat_i[28]_pad  ;
	input \wb_dat_i[29]_pad  ;
	input \wb_dat_i[2]_pad  ;
	input \wb_dat_i[30]_pad  ;
	input \wb_dat_i[31]_pad  ;
	input \wb_dat_i[3]_pad  ;
	input \wb_dat_i[4]_pad  ;
	input \wb_dat_i[5]_pad  ;
	input \wb_dat_i[6]_pad  ;
	input \wb_dat_i[7]_pad  ;
	input \wb_dat_i[8]_pad  ;
	input \wb_dat_i[9]_pad  ;
	input wb_int_o_pad ;
	input \wb_sel_i[0]_pad  ;
	input \wb_sel_i[1]_pad  ;
	input \wb_sel_i[2]_pad  ;
	input \wb_sel_i[3]_pad  ;
	input wb_stb_i_pad ;
	input wb_we_i_pad ;
	output \_al_n1  ;
	output \g10384/_0_  ;
	output \g10421/_0_  ;
	output \g10487/_0_  ;
	output \g10622/_0_  ;
	output \g10625/_0_  ;
	output \g10631/_3_  ;
	output \g10641/_0_  ;
	output \g10677/_3_  ;
	output \g10695/_0_  ;
	output \g10699/_3_  ;
	output \g10796/_0_  ;
	output \g10814/_00_  ;
	output \g10815/_0_  ;
	output \g10819/_0_  ;
	output \g10821/_0_  ;
	output \g10824/_3_  ;
	output \g10858/_0_  ;
	output \g11042/_00_  ;
	output \g11067/_0_  ;
	output \g11071/_00_  ;
	output \g11074/_0_  ;
	output \g11075/_0_  ;
	output \g11076/_0_  ;
	output \g11077/_0_  ;
	output \g11078/_0_  ;
	output \g11079/_0_  ;
	output \g11080/_0_  ;
	output \g11149/_0_  ;
	output \g11151/_0_  ;
	output \g11190/_00_  ;
	output \g11297/_0_  ;
	output \g11298/_0_  ;
	output \g11300/_0_  ;
	output \g11301/_0_  ;
	output \g11303/_0_  ;
	output \g11346/_0_  ;
	output \g11347/_0_  ;
	output \g11348/_0_  ;
	output \g11358/_0_  ;
	output \g11359/_0_  ;
	output \g11360/_0_  ;
	output \g11361/_0_  ;
	output \g11362/_0_  ;
	output \g11363/_0_  ;
	output \g11470/_0_  ;
	output \g11499/_0_  ;
	output \g11501/_0_  ;
	output \g11502/_0_  ;
	output \g11503/_0_  ;
	output \g11504/_0_  ;
	output \g11505/_0_  ;
	output \g11506/_0_  ;
	output \g11507/_0_  ;
	output \g11508/_0_  ;
	output \g11509/_0_  ;
	output \g11510/_0_  ;
	output \g11511/_0_  ;
	output \g11512/_0_  ;
	output \g11513/_0_  ;
	output \g11514/_0_  ;
	output \g11515/_0_  ;
	output \g11516/_0_  ;
	output \g11517/_0_  ;
	output \g11519/_0_  ;
	output \g11520/_0_  ;
	output \g11521/_0_  ;
	output \g11522/_0_  ;
	output \g11523/_0_  ;
	output \g11524/_0_  ;
	output \g11525/_0_  ;
	output \g11526/_0_  ;
	output \g11527/_0_  ;
	output \g11528/_0_  ;
	output \g11529/_0_  ;
	output \g11530/_0_  ;
	output \g11531/_0_  ;
	output \g11532/_0_  ;
	output \g11533/_0_  ;
	output \g11534/_0_  ;
	output \g11535/_0_  ;
	output \g11536/_0_  ;
	output \g11537/_0_  ;
	output \g11538/_0_  ;
	output \g11539/_0_  ;
	output \g11655/_0_  ;
	output \g11658/_0_  ;
	output \g11659/_0_  ;
	output \g11661/_0_  ;
	output \g11662/_0_  ;
	output \g11680/_0_  ;
	output \g11723/_0_  ;
	output \g11726/_0_  ;
	output \g11730/_0_  ;
	output \g11739/_0_  ;
	output \g11750/_0_  ;
	output \g11759/_0_  ;
	output \g11760/_0_  ;
	output \g11761/_0_  ;
	output \g11764/_0_  ;
	output \g11765/_0_  ;
	output \g12212/_0_  ;
	output \g13497/_0_  ;
	output \g13884/_0_  ;
	output \g13982/_0_  ;
	output \g13999/_0_  ;
	output \g9305/_0_  ;
	output \g9306/_0_  ;
	output \g9307/_0_  ;
	output \g9308/_0_  ;
	output \g9309/_0_  ;
	output \g9310/_0_  ;
	output \g9346/_0_  ;
	output \g9347/_0_  ;
	output \g9348/_0_  ;
	output \g9349/_0_  ;
	output \g9350/_0_  ;
	output \g9351/_0_  ;
	output \g9352/_0_  ;
	output \g9353/_0_  ;
	output \g9354/_0_  ;
	output \g9355/_0_  ;
	output \g9356/_0_  ;
	output \g9357/_0_  ;
	output \g9358/_0_  ;
	output \g9359/_0_  ;
	output \g9360/_0_  ;
	output \g9361/_0_  ;
	output \g9362/_0_  ;
	output \g9363/_0_  ;
	output \g9364/_0_  ;
	output \g9365/_0_  ;
	output \g9366/_0_  ;
	output \g9367/_0_  ;
	output \g9368/_0_  ;
	output \g9369/_0_  ;
	output \g9370/_0_  ;
	output \g9371/_0_  ;
	output \g9372/_0_  ;
	output \g9373/_0_  ;
	output \g9374/_0_  ;
	output \g9375/_0_  ;
	output \g9380/_0_  ;
	output \g9381/_0_  ;
	output \g9382/_0_  ;
	output \g9383/_0_  ;
	output \g9384/_0_  ;
	output \g9385/_0_  ;
	output \g9386/_0_  ;
	output \g9387/_0_  ;
	output \g9388/_0_  ;
	output \g9389/_0_  ;
	output \g9390/_0_  ;
	output \g9391/_0_  ;
	output \g9392/_0_  ;
	output \g9393/_0_  ;
	output \g9394/_0_  ;
	output \g9395/_0_  ;
	output \g9396/_0_  ;
	output \g9397/_0_  ;
	output \g9398/_0_  ;
	output \g9399/_0_  ;
	output \g9400/_0_  ;
	output \g9401/_0_  ;
	output \g9402/_0_  ;
	output \g9403/_0_  ;
	output \g9404/_0_  ;
	output \g9405/_0_  ;
	output \g9406/_0_  ;
	output \g9407/_0_  ;
	output \g9408/_0_  ;
	output \g9409/_0_  ;
	output \g9410/_0_  ;
	output \g9411/_0_  ;
	output \g9439/_0_  ;
	output \g9440/_0_  ;
	output \g9441/_0_  ;
	output \g9442/_0_  ;
	output \g9443/_0_  ;
	output \g9444/_0_  ;
	output \g9445/_0_  ;
	output \g9446/_0_  ;
	output \g9447/_0_  ;
	output \g9448/_0_  ;
	output \g9449/_0_  ;
	output \g9450/_0_  ;
	output \g9451/_0_  ;
	output \g9452/_0_  ;
	output \g9453/_0_  ;
	output \g9454/_0_  ;
	output \g9455/_0_  ;
	output \g9456/_0_  ;
	output \g9457/_0_  ;
	output \g9458/_0_  ;
	output \g9459/_0_  ;
	output \g9461/_0_  ;
	output \g9462/_0_  ;
	output \g9463/_0_  ;
	output \g9464/_0_  ;
	output \g9465/_0_  ;
	output \g9466/_0_  ;
	output \g9529/_0_  ;
	output \g9530/_0_  ;
	output \g9531/_0_  ;
	output \g9532/_0_  ;
	output \g9535/_0_  ;
	output \g9542/_0_  ;
	output \g9543/_0_  ;
	output \g9546/_0_  ;
	output \g9547/_0_  ;
	output \g9548/_0_  ;
	output \g9549/_0_  ;
	output \g9550/_0_  ;
	output \g9551/_0_  ;
	output \g9552/_0_  ;
	output \g9553/_0_  ;
	output \g9559/_0_  ;
	output \g9568/_0_  ;
	output \g9571/_0_  ;
	output \g9573/_0_  ;
	output \g9583/_0_  ;
	output \g9589/_0_  ;
	output \g9590/_0_  ;
	output \g9591/_0_  ;
	output \g9592/_0_  ;
	output \g9593/_0_  ;
	output \g9594/_0_  ;
	output \g9595/_0_  ;
	output \g9596/_0_  ;
	output \g9597/_0_  ;
	output \ss_pad_o[0]_pad  ;
	output \ss_pad_o[1]_pad  ;
	output \ss_pad_o[2]_pad  ;
	output \ss_pad_o[3]_pad  ;
	output \ss_pad_o[4]_pad  ;
	output \ss_pad_o[5]_pad  ;
	output \ss_pad_o[6]_pad  ;
	output \ss_pad_o[7]_pad  ;
	output wb_err_o_pad ;
	wire _w2278_ ;
	wire _w2277_ ;
	wire _w2276_ ;
	wire _w2275_ ;
	wire _w2274_ ;
	wire _w2273_ ;
	wire _w2272_ ;
	wire _w2271_ ;
	wire _w2270_ ;
	wire _w2269_ ;
	wire _w2268_ ;
	wire _w2267_ ;
	wire _w2266_ ;
	wire _w2265_ ;
	wire _w2264_ ;
	wire _w2263_ ;
	wire _w2262_ ;
	wire _w2261_ ;
	wire _w2260_ ;
	wire _w2259_ ;
	wire _w2258_ ;
	wire _w2257_ ;
	wire _w2256_ ;
	wire _w2255_ ;
	wire _w2254_ ;
	wire _w2253_ ;
	wire _w2252_ ;
	wire _w2251_ ;
	wire _w2250_ ;
	wire _w2249_ ;
	wire _w2248_ ;
	wire _w2247_ ;
	wire _w2246_ ;
	wire _w2245_ ;
	wire _w2244_ ;
	wire _w2243_ ;
	wire _w2242_ ;
	wire _w2241_ ;
	wire _w2240_ ;
	wire _w2239_ ;
	wire _w2238_ ;
	wire _w2237_ ;
	wire _w2236_ ;
	wire _w2235_ ;
	wire _w2234_ ;
	wire _w2233_ ;
	wire _w2232_ ;
	wire _w2231_ ;
	wire _w2230_ ;
	wire _w2229_ ;
	wire _w2228_ ;
	wire _w2227_ ;
	wire _w2226_ ;
	wire _w2225_ ;
	wire _w2224_ ;
	wire _w2223_ ;
	wire _w2222_ ;
	wire _w2221_ ;
	wire _w2220_ ;
	wire _w2219_ ;
	wire _w2218_ ;
	wire _w2217_ ;
	wire _w2216_ ;
	wire _w2215_ ;
	wire _w2214_ ;
	wire _w2213_ ;
	wire _w2212_ ;
	wire _w2211_ ;
	wire _w2210_ ;
	wire _w2209_ ;
	wire _w2208_ ;
	wire _w2207_ ;
	wire _w2206_ ;
	wire _w2205_ ;
	wire _w2204_ ;
	wire _w2203_ ;
	wire _w2202_ ;
	wire _w2201_ ;
	wire _w2200_ ;
	wire _w2199_ ;
	wire _w2198_ ;
	wire _w2197_ ;
	wire _w2196_ ;
	wire _w2195_ ;
	wire _w2194_ ;
	wire _w2193_ ;
	wire _w2192_ ;
	wire _w2191_ ;
	wire _w2190_ ;
	wire _w2189_ ;
	wire _w2188_ ;
	wire _w2187_ ;
	wire _w2186_ ;
	wire _w2185_ ;
	wire _w2184_ ;
	wire _w2183_ ;
	wire _w2182_ ;
	wire _w2181_ ;
	wire _w2180_ ;
	wire _w2179_ ;
	wire _w2178_ ;
	wire _w2177_ ;
	wire _w2176_ ;
	wire _w2175_ ;
	wire _w2174_ ;
	wire _w2173_ ;
	wire _w2172_ ;
	wire _w2171_ ;
	wire _w2170_ ;
	wire _w2169_ ;
	wire _w2168_ ;
	wire _w2167_ ;
	wire _w2166_ ;
	wire _w2165_ ;
	wire _w2164_ ;
	wire _w2163_ ;
	wire _w2162_ ;
	wire _w2161_ ;
	wire _w2160_ ;
	wire _w2159_ ;
	wire _w2158_ ;
	wire _w2157_ ;
	wire _w2156_ ;
	wire _w2155_ ;
	wire _w2154_ ;
	wire _w2153_ ;
	wire _w2152_ ;
	wire _w2151_ ;
	wire _w2150_ ;
	wire _w2149_ ;
	wire _w2148_ ;
	wire _w2147_ ;
	wire _w2146_ ;
	wire _w2145_ ;
	wire _w2144_ ;
	wire _w2143_ ;
	wire _w2142_ ;
	wire _w2141_ ;
	wire _w2140_ ;
	wire _w2139_ ;
	wire _w2138_ ;
	wire _w2137_ ;
	wire _w2136_ ;
	wire _w2135_ ;
	wire _w2134_ ;
	wire _w2133_ ;
	wire _w2132_ ;
	wire _w2131_ ;
	wire _w2130_ ;
	wire _w2129_ ;
	wire _w2128_ ;
	wire _w2127_ ;
	wire _w2126_ ;
	wire _w2125_ ;
	wire _w2124_ ;
	wire _w2123_ ;
	wire _w2122_ ;
	wire _w2121_ ;
	wire _w2120_ ;
	wire _w2119_ ;
	wire _w2118_ ;
	wire _w2117_ ;
	wire _w2116_ ;
	wire _w2115_ ;
	wire _w2114_ ;
	wire _w2113_ ;
	wire _w2112_ ;
	wire _w2111_ ;
	wire _w2110_ ;
	wire _w2109_ ;
	wire _w2108_ ;
	wire _w2107_ ;
	wire _w2106_ ;
	wire _w2105_ ;
	wire _w2104_ ;
	wire _w2103_ ;
	wire _w2102_ ;
	wire _w2101_ ;
	wire _w2100_ ;
	wire _w2099_ ;
	wire _w2098_ ;
	wire _w2097_ ;
	wire _w2096_ ;
	wire _w2095_ ;
	wire _w2094_ ;
	wire _w2093_ ;
	wire _w2092_ ;
	wire _w2091_ ;
	wire _w2090_ ;
	wire _w2089_ ;
	wire _w2088_ ;
	wire _w2087_ ;
	wire _w2086_ ;
	wire _w2085_ ;
	wire _w2084_ ;
	wire _w2083_ ;
	wire _w2082_ ;
	wire _w2081_ ;
	wire _w2080_ ;
	wire _w2079_ ;
	wire _w2078_ ;
	wire _w2077_ ;
	wire _w2076_ ;
	wire _w2075_ ;
	wire _w2074_ ;
	wire _w2073_ ;
	wire _w2072_ ;
	wire _w2071_ ;
	wire _w2070_ ;
	wire _w2069_ ;
	wire _w2068_ ;
	wire _w2067_ ;
	wire _w2066_ ;
	wire _w2065_ ;
	wire _w2064_ ;
	wire _w2063_ ;
	wire _w2062_ ;
	wire _w2061_ ;
	wire _w2060_ ;
	wire _w2059_ ;
	wire _w2058_ ;
	wire _w2057_ ;
	wire _w2056_ ;
	wire _w2055_ ;
	wire _w2054_ ;
	wire _w2053_ ;
	wire _w2052_ ;
	wire _w2051_ ;
	wire _w2050_ ;
	wire _w2049_ ;
	wire _w2048_ ;
	wire _w2047_ ;
	wire _w2046_ ;
	wire _w2045_ ;
	wire _w2044_ ;
	wire _w2043_ ;
	wire _w2042_ ;
	wire _w2041_ ;
	wire _w2040_ ;
	wire _w2039_ ;
	wire _w2038_ ;
	wire _w2037_ ;
	wire _w2036_ ;
	wire _w2035_ ;
	wire _w2034_ ;
	wire _w2033_ ;
	wire _w2032_ ;
	wire _w2031_ ;
	wire _w2030_ ;
	wire _w2029_ ;
	wire _w2028_ ;
	wire _w2027_ ;
	wire _w2026_ ;
	wire _w2025_ ;
	wire _w2024_ ;
	wire _w2023_ ;
	wire _w2022_ ;
	wire _w2021_ ;
	wire _w2020_ ;
	wire _w2019_ ;
	wire _w2018_ ;
	wire _w2017_ ;
	wire _w2016_ ;
	wire _w2015_ ;
	wire _w2014_ ;
	wire _w2013_ ;
	wire _w2012_ ;
	wire _w2011_ ;
	wire _w2010_ ;
	wire _w2009_ ;
	wire _w2008_ ;
	wire _w2007_ ;
	wire _w2006_ ;
	wire _w2005_ ;
	wire _w2004_ ;
	wire _w2003_ ;
	wire _w2002_ ;
	wire _w2001_ ;
	wire _w2000_ ;
	wire _w1999_ ;
	wire _w1998_ ;
	wire _w1997_ ;
	wire _w1996_ ;
	wire _w1995_ ;
	wire _w1994_ ;
	wire _w1993_ ;
	wire _w1992_ ;
	wire _w1991_ ;
	wire _w1990_ ;
	wire _w1989_ ;
	wire _w1988_ ;
	wire _w1987_ ;
	wire _w1986_ ;
	wire _w1985_ ;
	wire _w1984_ ;
	wire _w1983_ ;
	wire _w1982_ ;
	wire _w1981_ ;
	wire _w1980_ ;
	wire _w1979_ ;
	wire _w1978_ ;
	wire _w1977_ ;
	wire _w1976_ ;
	wire _w1975_ ;
	wire _w1974_ ;
	wire _w1973_ ;
	wire _w1972_ ;
	wire _w1971_ ;
	wire _w1970_ ;
	wire _w1969_ ;
	wire _w1968_ ;
	wire _w1967_ ;
	wire _w1966_ ;
	wire _w1965_ ;
	wire _w1964_ ;
	wire _w1963_ ;
	wire _w1962_ ;
	wire _w1961_ ;
	wire _w1960_ ;
	wire _w1959_ ;
	wire _w1958_ ;
	wire _w1957_ ;
	wire _w1956_ ;
	wire _w1955_ ;
	wire _w1954_ ;
	wire _w1953_ ;
	wire _w1952_ ;
	wire _w1951_ ;
	wire _w1950_ ;
	wire _w1949_ ;
	wire _w1948_ ;
	wire _w1947_ ;
	wire _w1946_ ;
	wire _w1945_ ;
	wire _w1944_ ;
	wire _w1943_ ;
	wire _w1942_ ;
	wire _w1941_ ;
	wire _w1940_ ;
	wire _w1939_ ;
	wire _w1938_ ;
	wire _w1937_ ;
	wire _w1936_ ;
	wire _w1935_ ;
	wire _w1934_ ;
	wire _w1933_ ;
	wire _w1932_ ;
	wire _w1931_ ;
	wire _w1930_ ;
	wire _w1929_ ;
	wire _w1928_ ;
	wire _w1927_ ;
	wire _w1926_ ;
	wire _w1925_ ;
	wire _w1924_ ;
	wire _w1923_ ;
	wire _w1922_ ;
	wire _w1921_ ;
	wire _w1920_ ;
	wire _w1919_ ;
	wire _w1918_ ;
	wire _w1917_ ;
	wire _w1916_ ;
	wire _w1915_ ;
	wire _w1914_ ;
	wire _w1913_ ;
	wire _w1912_ ;
	wire _w1911_ ;
	wire _w1910_ ;
	wire _w1909_ ;
	wire _w1908_ ;
	wire _w1907_ ;
	wire _w1906_ ;
	wire _w1905_ ;
	wire _w1904_ ;
	wire _w1903_ ;
	wire _w1902_ ;
	wire _w1901_ ;
	wire _w1900_ ;
	wire _w1899_ ;
	wire _w1898_ ;
	wire _w1897_ ;
	wire _w1896_ ;
	wire _w1895_ ;
	wire _w1894_ ;
	wire _w1893_ ;
	wire _w1892_ ;
	wire _w1891_ ;
	wire _w1890_ ;
	wire _w1889_ ;
	wire _w1888_ ;
	wire _w1887_ ;
	wire _w1886_ ;
	wire _w1885_ ;
	wire _w1884_ ;
	wire _w1883_ ;
	wire _w1882_ ;
	wire _w1881_ ;
	wire _w1880_ ;
	wire _w1879_ ;
	wire _w1878_ ;
	wire _w1877_ ;
	wire _w1876_ ;
	wire _w1875_ ;
	wire _w1874_ ;
	wire _w1873_ ;
	wire _w1872_ ;
	wire _w1871_ ;
	wire _w1870_ ;
	wire _w1869_ ;
	wire _w1868_ ;
	wire _w1867_ ;
	wire _w1866_ ;
	wire _w1865_ ;
	wire _w1864_ ;
	wire _w1863_ ;
	wire _w1862_ ;
	wire _w1861_ ;
	wire _w1860_ ;
	wire _w1859_ ;
	wire _w1858_ ;
	wire _w1857_ ;
	wire _w1856_ ;
	wire _w1855_ ;
	wire _w1854_ ;
	wire _w1853_ ;
	wire _w1852_ ;
	wire _w1851_ ;
	wire _w1850_ ;
	wire _w1849_ ;
	wire _w1848_ ;
	wire _w1847_ ;
	wire _w1846_ ;
	wire _w1845_ ;
	wire _w1844_ ;
	wire _w1843_ ;
	wire _w1842_ ;
	wire _w1841_ ;
	wire _w1840_ ;
	wire _w1839_ ;
	wire _w1838_ ;
	wire _w1837_ ;
	wire _w1836_ ;
	wire _w1835_ ;
	wire _w1834_ ;
	wire _w1833_ ;
	wire _w1832_ ;
	wire _w1831_ ;
	wire _w1830_ ;
	wire _w1829_ ;
	wire _w1828_ ;
	wire _w1827_ ;
	wire _w1826_ ;
	wire _w1825_ ;
	wire _w1824_ ;
	wire _w1823_ ;
	wire _w1822_ ;
	wire _w1821_ ;
	wire _w1820_ ;
	wire _w1819_ ;
	wire _w1818_ ;
	wire _w1817_ ;
	wire _w1816_ ;
	wire _w1815_ ;
	wire _w1814_ ;
	wire _w1813_ ;
	wire _w1812_ ;
	wire _w1811_ ;
	wire _w1810_ ;
	wire _w1809_ ;
	wire _w1808_ ;
	wire _w1807_ ;
	wire _w1806_ ;
	wire _w1805_ ;
	wire _w1804_ ;
	wire _w1803_ ;
	wire _w1802_ ;
	wire _w1801_ ;
	wire _w1800_ ;
	wire _w1799_ ;
	wire _w1798_ ;
	wire _w1797_ ;
	wire _w1796_ ;
	wire _w1795_ ;
	wire _w1794_ ;
	wire _w1793_ ;
	wire _w1792_ ;
	wire _w1791_ ;
	wire _w1790_ ;
	wire _w1789_ ;
	wire _w1788_ ;
	wire _w1787_ ;
	wire _w1786_ ;
	wire _w1785_ ;
	wire _w1784_ ;
	wire _w1783_ ;
	wire _w1782_ ;
	wire _w1781_ ;
	wire _w1780_ ;
	wire _w1779_ ;
	wire _w1778_ ;
	wire _w1777_ ;
	wire _w1776_ ;
	wire _w1775_ ;
	wire _w1774_ ;
	wire _w1773_ ;
	wire _w1772_ ;
	wire _w1771_ ;
	wire _w1770_ ;
	wire _w1769_ ;
	wire _w1768_ ;
	wire _w1767_ ;
	wire _w1766_ ;
	wire _w1765_ ;
	wire _w1764_ ;
	wire _w1763_ ;
	wire _w1762_ ;
	wire _w1761_ ;
	wire _w1760_ ;
	wire _w1759_ ;
	wire _w1758_ ;
	wire _w1757_ ;
	wire _w1756_ ;
	wire _w1755_ ;
	wire _w1754_ ;
	wire _w1753_ ;
	wire _w1752_ ;
	wire _w1751_ ;
	wire _w1750_ ;
	wire _w1749_ ;
	wire _w1748_ ;
	wire _w1747_ ;
	wire _w1746_ ;
	wire _w1745_ ;
	wire _w1744_ ;
	wire _w1743_ ;
	wire _w1742_ ;
	wire _w1741_ ;
	wire _w1740_ ;
	wire _w1739_ ;
	wire _w1738_ ;
	wire _w1737_ ;
	wire _w1736_ ;
	wire _w1735_ ;
	wire _w1734_ ;
	wire _w1733_ ;
	wire _w1732_ ;
	wire _w1731_ ;
	wire _w1730_ ;
	wire _w1729_ ;
	wire _w1728_ ;
	wire _w1727_ ;
	wire _w1726_ ;
	wire _w1725_ ;
	wire _w1724_ ;
	wire _w1723_ ;
	wire _w1722_ ;
	wire _w1721_ ;
	wire _w1720_ ;
	wire _w1719_ ;
	wire _w1718_ ;
	wire _w1717_ ;
	wire _w1716_ ;
	wire _w1715_ ;
	wire _w1714_ ;
	wire _w1713_ ;
	wire _w1712_ ;
	wire _w1711_ ;
	wire _w1710_ ;
	wire _w1709_ ;
	wire _w1708_ ;
	wire _w1707_ ;
	wire _w1706_ ;
	wire _w1705_ ;
	wire _w1704_ ;
	wire _w1703_ ;
	wire _w1702_ ;
	wire _w1701_ ;
	wire _w1700_ ;
	wire _w1699_ ;
	wire _w1698_ ;
	wire _w1697_ ;
	wire _w1696_ ;
	wire _w1695_ ;
	wire _w1694_ ;
	wire _w1693_ ;
	wire _w1692_ ;
	wire _w1691_ ;
	wire _w1690_ ;
	wire _w1689_ ;
	wire _w1688_ ;
	wire _w1687_ ;
	wire _w1686_ ;
	wire _w1685_ ;
	wire _w1684_ ;
	wire _w1683_ ;
	wire _w1682_ ;
	wire _w1681_ ;
	wire _w1680_ ;
	wire _w1679_ ;
	wire _w1678_ ;
	wire _w1677_ ;
	wire _w1676_ ;
	wire _w1675_ ;
	wire _w1674_ ;
	wire _w1673_ ;
	wire _w1672_ ;
	wire _w1671_ ;
	wire _w1670_ ;
	wire _w1669_ ;
	wire _w1668_ ;
	wire _w1667_ ;
	wire _w1666_ ;
	wire _w1665_ ;
	wire _w1664_ ;
	wire _w1663_ ;
	wire _w1662_ ;
	wire _w1661_ ;
	wire _w1660_ ;
	wire _w1659_ ;
	wire _w1658_ ;
	wire _w1657_ ;
	wire _w1656_ ;
	wire _w1655_ ;
	wire _w1654_ ;
	wire _w1653_ ;
	wire _w1652_ ;
	wire _w1651_ ;
	wire _w1650_ ;
	wire _w1649_ ;
	wire _w1648_ ;
	wire _w1647_ ;
	wire _w1646_ ;
	wire _w1645_ ;
	wire _w1644_ ;
	wire _w1643_ ;
	wire _w1642_ ;
	wire _w1641_ ;
	wire _w1640_ ;
	wire _w1639_ ;
	wire _w1638_ ;
	wire _w1637_ ;
	wire _w1636_ ;
	wire _w1635_ ;
	wire _w1634_ ;
	wire _w1633_ ;
	wire _w1632_ ;
	wire _w1631_ ;
	wire _w1630_ ;
	wire _w1629_ ;
	wire _w1628_ ;
	wire _w1627_ ;
	wire _w1626_ ;
	wire _w1625_ ;
	wire _w1624_ ;
	wire _w1623_ ;
	wire _w1622_ ;
	wire _w1621_ ;
	wire _w1620_ ;
	wire _w1619_ ;
	wire _w1618_ ;
	wire _w1617_ ;
	wire _w1616_ ;
	wire _w1615_ ;
	wire _w1614_ ;
	wire _w1613_ ;
	wire _w1612_ ;
	wire _w1611_ ;
	wire _w1610_ ;
	wire _w1609_ ;
	wire _w1608_ ;
	wire _w1607_ ;
	wire _w1606_ ;
	wire _w1605_ ;
	wire _w1604_ ;
	wire _w1603_ ;
	wire _w1602_ ;
	wire _w1601_ ;
	wire _w1600_ ;
	wire _w1599_ ;
	wire _w1598_ ;
	wire _w1597_ ;
	wire _w1596_ ;
	wire _w1595_ ;
	wire _w1594_ ;
	wire _w1593_ ;
	wire _w1592_ ;
	wire _w1591_ ;
	wire _w1590_ ;
	wire _w1589_ ;
	wire _w1588_ ;
	wire _w1587_ ;
	wire _w1586_ ;
	wire _w1585_ ;
	wire _w1584_ ;
	wire _w1583_ ;
	wire _w1582_ ;
	wire _w1581_ ;
	wire _w1580_ ;
	wire _w1579_ ;
	wire _w1578_ ;
	wire _w1577_ ;
	wire _w1576_ ;
	wire _w1575_ ;
	wire _w1574_ ;
	wire _w1573_ ;
	wire _w1572_ ;
	wire _w1571_ ;
	wire _w1570_ ;
	wire _w1569_ ;
	wire _w1568_ ;
	wire _w1567_ ;
	wire _w1566_ ;
	wire _w1565_ ;
	wire _w1564_ ;
	wire _w1563_ ;
	wire _w1562_ ;
	wire _w1561_ ;
	wire _w1560_ ;
	wire _w1559_ ;
	wire _w1558_ ;
	wire _w1557_ ;
	wire _w1556_ ;
	wire _w1555_ ;
	wire _w1554_ ;
	wire _w1553_ ;
	wire _w1552_ ;
	wire _w1551_ ;
	wire _w1550_ ;
	wire _w1549_ ;
	wire _w1548_ ;
	wire _w1547_ ;
	wire _w1546_ ;
	wire _w1545_ ;
	wire _w1544_ ;
	wire _w1543_ ;
	wire _w1542_ ;
	wire _w1541_ ;
	wire _w1540_ ;
	wire _w1539_ ;
	wire _w1538_ ;
	wire _w1537_ ;
	wire _w1536_ ;
	wire _w1535_ ;
	wire _w1534_ ;
	wire _w1533_ ;
	wire _w1532_ ;
	wire _w1531_ ;
	wire _w1530_ ;
	wire _w1529_ ;
	wire _w1528_ ;
	wire _w1527_ ;
	wire _w1526_ ;
	wire _w1525_ ;
	wire _w1524_ ;
	wire _w1523_ ;
	wire _w1522_ ;
	wire _w1521_ ;
	wire _w1520_ ;
	wire _w1519_ ;
	wire _w1518_ ;
	wire _w1517_ ;
	wire _w1516_ ;
	wire _w1515_ ;
	wire _w1514_ ;
	wire _w1513_ ;
	wire _w1512_ ;
	wire _w1511_ ;
	wire _w1510_ ;
	wire _w1509_ ;
	wire _w1508_ ;
	wire _w1507_ ;
	wire _w1506_ ;
	wire _w1505_ ;
	wire _w1504_ ;
	wire _w1503_ ;
	wire _w1502_ ;
	wire _w1501_ ;
	wire _w1500_ ;
	wire _w1499_ ;
	wire _w1498_ ;
	wire _w1497_ ;
	wire _w1496_ ;
	wire _w1495_ ;
	wire _w1494_ ;
	wire _w1493_ ;
	wire _w1492_ ;
	wire _w1491_ ;
	wire _w1490_ ;
	wire _w1489_ ;
	wire _w1488_ ;
	wire _w1487_ ;
	wire _w1486_ ;
	wire _w1485_ ;
	wire _w1484_ ;
	wire _w1483_ ;
	wire _w1482_ ;
	wire _w1481_ ;
	wire _w1480_ ;
	wire _w1479_ ;
	wire _w1478_ ;
	wire _w1477_ ;
	wire _w1476_ ;
	wire _w1475_ ;
	wire _w1474_ ;
	wire _w1473_ ;
	wire _w1472_ ;
	wire _w1471_ ;
	wire _w1470_ ;
	wire _w1469_ ;
	wire _w1468_ ;
	wire _w1467_ ;
	wire _w1466_ ;
	wire _w1465_ ;
	wire _w1464_ ;
	wire _w1463_ ;
	wire _w1462_ ;
	wire _w1461_ ;
	wire _w1460_ ;
	wire _w1459_ ;
	wire _w1458_ ;
	wire _w1457_ ;
	wire _w1456_ ;
	wire _w1455_ ;
	wire _w1454_ ;
	wire _w1453_ ;
	wire _w1452_ ;
	wire _w1451_ ;
	wire _w1450_ ;
	wire _w1449_ ;
	wire _w1448_ ;
	wire _w1447_ ;
	wire _w1446_ ;
	wire _w1445_ ;
	wire _w1444_ ;
	wire _w1443_ ;
	wire _w1442_ ;
	wire _w1441_ ;
	wire _w1440_ ;
	wire _w1439_ ;
	wire _w1438_ ;
	wire _w1437_ ;
	wire _w1436_ ;
	wire _w1435_ ;
	wire _w1434_ ;
	wire _w1433_ ;
	wire _w1432_ ;
	wire _w1431_ ;
	wire _w1430_ ;
	wire _w1429_ ;
	wire _w1428_ ;
	wire _w1427_ ;
	wire _w1426_ ;
	wire _w1425_ ;
	wire _w1424_ ;
	wire _w1423_ ;
	wire _w1422_ ;
	wire _w1421_ ;
	wire _w1420_ ;
	wire _w1419_ ;
	wire _w1418_ ;
	wire _w1417_ ;
	wire _w1416_ ;
	wire _w1415_ ;
	wire _w1414_ ;
	wire _w1413_ ;
	wire _w1412_ ;
	wire _w1411_ ;
	wire _w1410_ ;
	wire _w1409_ ;
	wire _w1408_ ;
	wire _w1407_ ;
	wire _w1406_ ;
	wire _w1405_ ;
	wire _w1404_ ;
	wire _w1403_ ;
	wire _w1402_ ;
	wire _w1401_ ;
	wire _w1400_ ;
	wire _w1399_ ;
	wire _w1398_ ;
	wire _w1397_ ;
	wire _w1396_ ;
	wire _w1395_ ;
	wire _w1394_ ;
	wire _w1393_ ;
	wire _w1392_ ;
	wire _w1391_ ;
	wire _w1390_ ;
	wire _w1389_ ;
	wire _w1388_ ;
	wire _w1387_ ;
	wire _w1386_ ;
	wire _w1385_ ;
	wire _w1384_ ;
	wire _w1383_ ;
	wire _w1382_ ;
	wire _w1381_ ;
	wire _w1380_ ;
	wire _w1379_ ;
	wire _w1378_ ;
	wire _w1377_ ;
	wire _w1376_ ;
	wire _w1375_ ;
	wire _w1374_ ;
	wire _w1373_ ;
	wire _w1372_ ;
	wire _w1371_ ;
	wire _w1370_ ;
	wire _w1369_ ;
	wire _w1368_ ;
	wire _w1367_ ;
	wire _w1366_ ;
	wire _w1365_ ;
	wire _w1364_ ;
	wire _w1363_ ;
	wire _w1362_ ;
	wire _w1361_ ;
	wire _w1360_ ;
	wire _w1359_ ;
	wire _w1358_ ;
	wire _w1357_ ;
	wire _w1356_ ;
	wire _w1355_ ;
	wire _w1354_ ;
	wire _w1353_ ;
	wire _w1352_ ;
	wire _w1351_ ;
	wire _w782_ ;
	wire _w781_ ;
	wire _w780_ ;
	wire _w779_ ;
	wire _w778_ ;
	wire _w777_ ;
	wire _w776_ ;
	wire _w775_ ;
	wire _w774_ ;
	wire _w773_ ;
	wire _w772_ ;
	wire _w771_ ;
	wire _w770_ ;
	wire _w769_ ;
	wire _w768_ ;
	wire _w767_ ;
	wire _w766_ ;
	wire _w765_ ;
	wire _w764_ ;
	wire _w763_ ;
	wire _w762_ ;
	wire _w761_ ;
	wire _w760_ ;
	wire _w759_ ;
	wire _w758_ ;
	wire _w757_ ;
	wire _w756_ ;
	wire _w755_ ;
	wire _w754_ ;
	wire _w753_ ;
	wire _w752_ ;
	wire _w751_ ;
	wire _w750_ ;
	wire _w749_ ;
	wire _w748_ ;
	wire _w747_ ;
	wire _w746_ ;
	wire _w745_ ;
	wire _w744_ ;
	wire _w743_ ;
	wire _w742_ ;
	wire _w741_ ;
	wire _w740_ ;
	wire _w739_ ;
	wire _w738_ ;
	wire _w737_ ;
	wire _w736_ ;
	wire _w735_ ;
	wire _w734_ ;
	wire _w733_ ;
	wire _w732_ ;
	wire _w731_ ;
	wire _w730_ ;
	wire _w729_ ;
	wire _w728_ ;
	wire _w727_ ;
	wire _w726_ ;
	wire _w725_ ;
	wire _w724_ ;
	wire _w723_ ;
	wire _w722_ ;
	wire _w721_ ;
	wire _w720_ ;
	wire _w719_ ;
	wire _w718_ ;
	wire _w717_ ;
	wire _w716_ ;
	wire _w715_ ;
	wire _w714_ ;
	wire _w713_ ;
	wire _w712_ ;
	wire _w711_ ;
	wire _w710_ ;
	wire _w709_ ;
	wire _w708_ ;
	wire _w707_ ;
	wire _w706_ ;
	wire _w705_ ;
	wire _w704_ ;
	wire _w703_ ;
	wire _w702_ ;
	wire _w701_ ;
	wire _w700_ ;
	wire _w699_ ;
	wire _w698_ ;
	wire _w697_ ;
	wire _w696_ ;
	wire _w695_ ;
	wire _w694_ ;
	wire _w693_ ;
	wire _w692_ ;
	wire _w691_ ;
	wire _w690_ ;
	wire _w689_ ;
	wire _w688_ ;
	wire _w687_ ;
	wire _w686_ ;
	wire _w685_ ;
	wire _w684_ ;
	wire _w683_ ;
	wire _w682_ ;
	wire _w681_ ;
	wire _w680_ ;
	wire _w679_ ;
	wire _w678_ ;
	wire _w677_ ;
	wire _w676_ ;
	wire _w675_ ;
	wire _w674_ ;
	wire _w673_ ;
	wire _w672_ ;
	wire _w671_ ;
	wire _w670_ ;
	wire _w669_ ;
	wire _w668_ ;
	wire _w667_ ;
	wire _w666_ ;
	wire _w665_ ;
	wire _w664_ ;
	wire _w663_ ;
	wire _w662_ ;
	wire _w661_ ;
	wire _w660_ ;
	wire _w659_ ;
	wire _w658_ ;
	wire _w657_ ;
	wire _w656_ ;
	wire _w655_ ;
	wire _w654_ ;
	wire _w653_ ;
	wire _w652_ ;
	wire _w651_ ;
	wire _w650_ ;
	wire _w649_ ;
	wire _w648_ ;
	wire _w647_ ;
	wire _w646_ ;
	wire _w645_ ;
	wire _w644_ ;
	wire _w643_ ;
	wire _w642_ ;
	wire _w641_ ;
	wire _w640_ ;
	wire _w639_ ;
	wire _w638_ ;
	wire _w637_ ;
	wire _w636_ ;
	wire _w635_ ;
	wire _w634_ ;
	wire _w633_ ;
	wire _w632_ ;
	wire _w631_ ;
	wire _w630_ ;
	wire _w629_ ;
	wire _w628_ ;
	wire _w627_ ;
	wire _w626_ ;
	wire _w625_ ;
	wire _w624_ ;
	wire _w623_ ;
	wire _w622_ ;
	wire _w621_ ;
	wire _w620_ ;
	wire _w619_ ;
	wire _w618_ ;
	wire _w617_ ;
	wire _w616_ ;
	wire _w615_ ;
	wire _w614_ ;
	wire _w613_ ;
	wire _w612_ ;
	wire _w611_ ;
	wire _w610_ ;
	wire _w609_ ;
	wire _w608_ ;
	wire _w607_ ;
	wire _w606_ ;
	wire _w605_ ;
	wire _w604_ ;
	wire _w603_ ;
	wire _w602_ ;
	wire _w601_ ;
	wire _w600_ ;
	wire _w599_ ;
	wire _w598_ ;
	wire _w597_ ;
	wire _w596_ ;
	wire _w595_ ;
	wire _w594_ ;
	wire _w593_ ;
	wire _w592_ ;
	wire _w591_ ;
	wire _w590_ ;
	wire _w589_ ;
	wire _w588_ ;
	wire _w587_ ;
	wire _w586_ ;
	wire _w585_ ;
	wire _w584_ ;
	wire _w583_ ;
	wire _w582_ ;
	wire _w581_ ;
	wire _w580_ ;
	wire _w579_ ;
	wire _w578_ ;
	wire _w577_ ;
	wire _w576_ ;
	wire _w575_ ;
	wire _w574_ ;
	wire _w573_ ;
	wire _w572_ ;
	wire _w571_ ;
	wire _w570_ ;
	wire _w569_ ;
	wire _w568_ ;
	wire _w567_ ;
	wire _w566_ ;
	wire _w565_ ;
	wire _w564_ ;
	wire _w563_ ;
	wire _w562_ ;
	wire _w561_ ;
	wire _w560_ ;
	wire _w559_ ;
	wire _w558_ ;
	wire _w557_ ;
	wire _w556_ ;
	wire _w555_ ;
	wire _w554_ ;
	wire _w553_ ;
	wire _w552_ ;
	wire _w551_ ;
	wire _w550_ ;
	wire _w549_ ;
	wire _w548_ ;
	wire _w547_ ;
	wire _w546_ ;
	wire _w545_ ;
	wire _w544_ ;
	wire _w543_ ;
	wire _w542_ ;
	wire _w541_ ;
	wire _w540_ ;
	wire _w539_ ;
	wire _w538_ ;
	wire _w537_ ;
	wire _w536_ ;
	wire _w535_ ;
	wire _w534_ ;
	wire _w533_ ;
	wire _w532_ ;
	wire _w531_ ;
	wire _w530_ ;
	wire _w529_ ;
	wire _w528_ ;
	wire _w527_ ;
	wire _w526_ ;
	wire _w525_ ;
	wire _w524_ ;
	wire _w523_ ;
	wire _w522_ ;
	wire _w521_ ;
	wire _w520_ ;
	wire _w519_ ;
	wire _w518_ ;
	wire _w517_ ;
	wire _w516_ ;
	wire _w515_ ;
	wire _w514_ ;
	wire _w513_ ;
	wire _w512_ ;
	wire _w511_ ;
	wire _w510_ ;
	wire _w509_ ;
	wire _w508_ ;
	wire _w507_ ;
	wire _w506_ ;
	wire _w505_ ;
	wire _w504_ ;
	wire _w503_ ;
	wire _w502_ ;
	wire _w501_ ;
	wire _w500_ ;
	wire _w499_ ;
	wire _w368_ ;
	wire _w367_ ;
	wire _w366_ ;
	wire _w365_ ;
	wire _w364_ ;
	wire _w363_ ;
	wire _w362_ ;
	wire _w361_ ;
	wire _w360_ ;
	wire _w359_ ;
	wire _w358_ ;
	wire _w357_ ;
	wire _w356_ ;
	wire _w355_ ;
	wire _w354_ ;
	wire _w353_ ;
	wire _w352_ ;
	wire _w351_ ;
	wire _w350_ ;
	wire _w349_ ;
	wire _w348_ ;
	wire _w347_ ;
	wire _w346_ ;
	wire _w345_ ;
	wire _w344_ ;
	wire _w343_ ;
	wire _w342_ ;
	wire _w341_ ;
	wire _w340_ ;
	wire _w339_ ;
	wire _w338_ ;
	wire _w337_ ;
	wire _w336_ ;
	wire _w335_ ;
	wire _w334_ ;
	wire _w333_ ;
	wire _w332_ ;
	wire _w331_ ;
	wire _w330_ ;
	wire _w329_ ;
	wire _w328_ ;
	wire _w327_ ;
	wire _w326_ ;
	wire _w325_ ;
	wire _w324_ ;
	wire _w323_ ;
	wire _w322_ ;
	wire _w321_ ;
	wire _w320_ ;
	wire _w319_ ;
	wire _w318_ ;
	wire _w317_ ;
	wire _w316_ ;
	wire _w315_ ;
	wire _w314_ ;
	wire _w313_ ;
	wire _w312_ ;
	wire _w311_ ;
	wire _w310_ ;
	wire _w309_ ;
	wire _w308_ ;
	wire _w307_ ;
	wire _w306_ ;
	wire _w305_ ;
	wire _w304_ ;
	wire _w303_ ;
	wire _w302_ ;
	wire _w301_ ;
	wire _w270_ ;
	wire _w269_ ;
	wire _w268_ ;
	wire _w267_ ;
	wire _w266_ ;
	wire _w265_ ;
	wire _w264_ ;
	wire _w263_ ;
	wire _w262_ ;
	wire _w261_ ;
	wire _w260_ ;
	wire _w259_ ;
	wire _w258_ ;
	wire _w257_ ;
	wire _w256_ ;
	wire _w255_ ;
	wire _w242_ ;
	wire _w243_ ;
	wire _w244_ ;
	wire _w245_ ;
	wire _w246_ ;
	wire _w247_ ;
	wire _w248_ ;
	wire _w249_ ;
	wire _w250_ ;
	wire _w251_ ;
	wire _w252_ ;
	wire _w253_ ;
	wire _w254_ ;
	wire _w271_ ;
	wire _w272_ ;
	wire _w273_ ;
	wire _w274_ ;
	wire _w275_ ;
	wire _w276_ ;
	wire _w277_ ;
	wire _w278_ ;
	wire _w279_ ;
	wire _w280_ ;
	wire _w281_ ;
	wire _w282_ ;
	wire _w283_ ;
	wire _w284_ ;
	wire _w285_ ;
	wire _w286_ ;
	wire _w287_ ;
	wire _w288_ ;
	wire _w289_ ;
	wire _w290_ ;
	wire _w291_ ;
	wire _w292_ ;
	wire _w293_ ;
	wire _w294_ ;
	wire _w295_ ;
	wire _w296_ ;
	wire _w297_ ;
	wire _w298_ ;
	wire _w299_ ;
	wire _w300_ ;
	wire _w369_ ;
	wire _w370_ ;
	wire _w371_ ;
	wire _w372_ ;
	wire _w373_ ;
	wire _w374_ ;
	wire _w375_ ;
	wire _w376_ ;
	wire _w377_ ;
	wire _w378_ ;
	wire _w379_ ;
	wire _w380_ ;
	wire _w381_ ;
	wire _w382_ ;
	wire _w383_ ;
	wire _w384_ ;
	wire _w385_ ;
	wire _w386_ ;
	wire _w387_ ;
	wire _w388_ ;
	wire _w389_ ;
	wire _w390_ ;
	wire _w391_ ;
	wire _w392_ ;
	wire _w393_ ;
	wire _w394_ ;
	wire _w395_ ;
	wire _w396_ ;
	wire _w397_ ;
	wire _w398_ ;
	wire _w399_ ;
	wire _w400_ ;
	wire _w401_ ;
	wire _w402_ ;
	wire _w403_ ;
	wire _w404_ ;
	wire _w405_ ;
	wire _w406_ ;
	wire _w407_ ;
	wire _w408_ ;
	wire _w409_ ;
	wire _w410_ ;
	wire _w411_ ;
	wire _w412_ ;
	wire _w413_ ;
	wire _w414_ ;
	wire _w415_ ;
	wire _w416_ ;
	wire _w417_ ;
	wire _w418_ ;
	wire _w419_ ;
	wire _w420_ ;
	wire _w421_ ;
	wire _w422_ ;
	wire _w423_ ;
	wire _w424_ ;
	wire _w425_ ;
	wire _w426_ ;
	wire _w427_ ;
	wire _w428_ ;
	wire _w429_ ;
	wire _w430_ ;
	wire _w431_ ;
	wire _w432_ ;
	wire _w433_ ;
	wire _w434_ ;
	wire _w435_ ;
	wire _w436_ ;
	wire _w437_ ;
	wire _w438_ ;
	wire _w439_ ;
	wire _w440_ ;
	wire _w441_ ;
	wire _w442_ ;
	wire _w443_ ;
	wire _w444_ ;
	wire _w445_ ;
	wire _w446_ ;
	wire _w447_ ;
	wire _w448_ ;
	wire _w449_ ;
	wire _w450_ ;
	wire _w451_ ;
	wire _w452_ ;
	wire _w453_ ;
	wire _w454_ ;
	wire _w455_ ;
	wire _w456_ ;
	wire _w457_ ;
	wire _w458_ ;
	wire _w459_ ;
	wire _w460_ ;
	wire _w461_ ;
	wire _w462_ ;
	wire _w463_ ;
	wire _w464_ ;
	wire _w465_ ;
	wire _w466_ ;
	wire _w467_ ;
	wire _w468_ ;
	wire _w469_ ;
	wire _w470_ ;
	wire _w471_ ;
	wire _w472_ ;
	wire _w473_ ;
	wire _w474_ ;
	wire _w475_ ;
	wire _w476_ ;
	wire _w477_ ;
	wire _w478_ ;
	wire _w479_ ;
	wire _w480_ ;
	wire _w481_ ;
	wire _w482_ ;
	wire _w483_ ;
	wire _w484_ ;
	wire _w485_ ;
	wire _w486_ ;
	wire _w487_ ;
	wire _w488_ ;
	wire _w489_ ;
	wire _w490_ ;
	wire _w491_ ;
	wire _w492_ ;
	wire _w493_ ;
	wire _w494_ ;
	wire _w495_ ;
	wire _w496_ ;
	wire _w497_ ;
	wire _w498_ ;
	wire _w783_ ;
	wire _w784_ ;
	wire _w785_ ;
	wire _w786_ ;
	wire _w787_ ;
	wire _w788_ ;
	wire _w789_ ;
	wire _w790_ ;
	wire _w791_ ;
	wire _w792_ ;
	wire _w793_ ;
	wire _w794_ ;
	wire _w795_ ;
	wire _w796_ ;
	wire _w797_ ;
	wire _w798_ ;
	wire _w799_ ;
	wire _w800_ ;
	wire _w801_ ;
	wire _w802_ ;
	wire _w803_ ;
	wire _w804_ ;
	wire _w805_ ;
	wire _w806_ ;
	wire _w807_ ;
	wire _w808_ ;
	wire _w809_ ;
	wire _w810_ ;
	wire _w811_ ;
	wire _w812_ ;
	wire _w813_ ;
	wire _w814_ ;
	wire _w815_ ;
	wire _w816_ ;
	wire _w817_ ;
	wire _w818_ ;
	wire _w819_ ;
	wire _w820_ ;
	wire _w821_ ;
	wire _w822_ ;
	wire _w823_ ;
	wire _w824_ ;
	wire _w825_ ;
	wire _w826_ ;
	wire _w827_ ;
	wire _w828_ ;
	wire _w829_ ;
	wire _w830_ ;
	wire _w831_ ;
	wire _w832_ ;
	wire _w833_ ;
	wire _w834_ ;
	wire _w835_ ;
	wire _w836_ ;
	wire _w837_ ;
	wire _w838_ ;
	wire _w839_ ;
	wire _w840_ ;
	wire _w841_ ;
	wire _w842_ ;
	wire _w843_ ;
	wire _w844_ ;
	wire _w845_ ;
	wire _w846_ ;
	wire _w847_ ;
	wire _w848_ ;
	wire _w849_ ;
	wire _w850_ ;
	wire _w851_ ;
	wire _w852_ ;
	wire _w853_ ;
	wire _w854_ ;
	wire _w855_ ;
	wire _w856_ ;
	wire _w857_ ;
	wire _w858_ ;
	wire _w859_ ;
	wire _w860_ ;
	wire _w861_ ;
	wire _w862_ ;
	wire _w863_ ;
	wire _w864_ ;
	wire _w865_ ;
	wire _w866_ ;
	wire _w867_ ;
	wire _w868_ ;
	wire _w869_ ;
	wire _w870_ ;
	wire _w871_ ;
	wire _w872_ ;
	wire _w873_ ;
	wire _w874_ ;
	wire _w875_ ;
	wire _w876_ ;
	wire _w877_ ;
	wire _w878_ ;
	wire _w879_ ;
	wire _w880_ ;
	wire _w881_ ;
	wire _w882_ ;
	wire _w883_ ;
	wire _w884_ ;
	wire _w885_ ;
	wire _w886_ ;
	wire _w887_ ;
	wire _w888_ ;
	wire _w889_ ;
	wire _w890_ ;
	wire _w891_ ;
	wire _w892_ ;
	wire _w893_ ;
	wire _w894_ ;
	wire _w895_ ;
	wire _w896_ ;
	wire _w897_ ;
	wire _w898_ ;
	wire _w899_ ;
	wire _w900_ ;
	wire _w901_ ;
	wire _w902_ ;
	wire _w903_ ;
	wire _w904_ ;
	wire _w905_ ;
	wire _w906_ ;
	wire _w907_ ;
	wire _w908_ ;
	wire _w909_ ;
	wire _w910_ ;
	wire _w911_ ;
	wire _w912_ ;
	wire _w913_ ;
	wire _w914_ ;
	wire _w915_ ;
	wire _w916_ ;
	wire _w917_ ;
	wire _w918_ ;
	wire _w919_ ;
	wire _w920_ ;
	wire _w921_ ;
	wire _w922_ ;
	wire _w923_ ;
	wire _w924_ ;
	wire _w925_ ;
	wire _w926_ ;
	wire _w927_ ;
	wire _w928_ ;
	wire _w929_ ;
	wire _w930_ ;
	wire _w931_ ;
	wire _w932_ ;
	wire _w933_ ;
	wire _w934_ ;
	wire _w935_ ;
	wire _w936_ ;
	wire _w937_ ;
	wire _w938_ ;
	wire _w939_ ;
	wire _w940_ ;
	wire _w941_ ;
	wire _w942_ ;
	wire _w943_ ;
	wire _w944_ ;
	wire _w945_ ;
	wire _w946_ ;
	wire _w947_ ;
	wire _w948_ ;
	wire _w949_ ;
	wire _w950_ ;
	wire _w951_ ;
	wire _w952_ ;
	wire _w953_ ;
	wire _w954_ ;
	wire _w955_ ;
	wire _w956_ ;
	wire _w957_ ;
	wire _w958_ ;
	wire _w959_ ;
	wire _w960_ ;
	wire _w961_ ;
	wire _w962_ ;
	wire _w963_ ;
	wire _w964_ ;
	wire _w965_ ;
	wire _w966_ ;
	wire _w967_ ;
	wire _w968_ ;
	wire _w969_ ;
	wire _w970_ ;
	wire _w971_ ;
	wire _w972_ ;
	wire _w973_ ;
	wire _w974_ ;
	wire _w975_ ;
	wire _w976_ ;
	wire _w977_ ;
	wire _w978_ ;
	wire _w979_ ;
	wire _w980_ ;
	wire _w981_ ;
	wire _w982_ ;
	wire _w983_ ;
	wire _w984_ ;
	wire _w985_ ;
	wire _w986_ ;
	wire _w987_ ;
	wire _w988_ ;
	wire _w989_ ;
	wire _w990_ ;
	wire _w991_ ;
	wire _w992_ ;
	wire _w993_ ;
	wire _w994_ ;
	wire _w995_ ;
	wire _w996_ ;
	wire _w997_ ;
	wire _w998_ ;
	wire _w999_ ;
	wire _w1000_ ;
	wire _w1001_ ;
	wire _w1002_ ;
	wire _w1003_ ;
	wire _w1004_ ;
	wire _w1005_ ;
	wire _w1006_ ;
	wire _w1007_ ;
	wire _w1008_ ;
	wire _w1009_ ;
	wire _w1010_ ;
	wire _w1011_ ;
	wire _w1012_ ;
	wire _w1013_ ;
	wire _w1014_ ;
	wire _w1015_ ;
	wire _w1016_ ;
	wire _w1017_ ;
	wire _w1018_ ;
	wire _w1019_ ;
	wire _w1020_ ;
	wire _w1021_ ;
	wire _w1022_ ;
	wire _w1023_ ;
	wire _w1024_ ;
	wire _w1025_ ;
	wire _w1026_ ;
	wire _w1027_ ;
	wire _w1028_ ;
	wire _w1029_ ;
	wire _w1030_ ;
	wire _w1031_ ;
	wire _w1032_ ;
	wire _w1033_ ;
	wire _w1034_ ;
	wire _w1035_ ;
	wire _w1036_ ;
	wire _w1037_ ;
	wire _w1038_ ;
	wire _w1039_ ;
	wire _w1040_ ;
	wire _w1041_ ;
	wire _w1042_ ;
	wire _w1043_ ;
	wire _w1044_ ;
	wire _w1045_ ;
	wire _w1046_ ;
	wire _w1047_ ;
	wire _w1048_ ;
	wire _w1049_ ;
	wire _w1050_ ;
	wire _w1051_ ;
	wire _w1052_ ;
	wire _w1053_ ;
	wire _w1054_ ;
	wire _w1055_ ;
	wire _w1056_ ;
	wire _w1057_ ;
	wire _w1058_ ;
	wire _w1059_ ;
	wire _w1060_ ;
	wire _w1061_ ;
	wire _w1062_ ;
	wire _w1063_ ;
	wire _w1064_ ;
	wire _w1065_ ;
	wire _w1066_ ;
	wire _w1067_ ;
	wire _w1068_ ;
	wire _w1069_ ;
	wire _w1070_ ;
	wire _w1071_ ;
	wire _w1072_ ;
	wire _w1073_ ;
	wire _w1074_ ;
	wire _w1075_ ;
	wire _w1076_ ;
	wire _w1077_ ;
	wire _w1078_ ;
	wire _w1079_ ;
	wire _w1080_ ;
	wire _w1081_ ;
	wire _w1082_ ;
	wire _w1083_ ;
	wire _w1084_ ;
	wire _w1085_ ;
	wire _w1086_ ;
	wire _w1087_ ;
	wire _w1088_ ;
	wire _w1089_ ;
	wire _w1090_ ;
	wire _w1091_ ;
	wire _w1092_ ;
	wire _w1093_ ;
	wire _w1094_ ;
	wire _w1095_ ;
	wire _w1096_ ;
	wire _w1097_ ;
	wire _w1098_ ;
	wire _w1099_ ;
	wire _w1100_ ;
	wire _w1101_ ;
	wire _w1102_ ;
	wire _w1103_ ;
	wire _w1104_ ;
	wire _w1105_ ;
	wire _w1106_ ;
	wire _w1107_ ;
	wire _w1108_ ;
	wire _w1109_ ;
	wire _w1110_ ;
	wire _w1111_ ;
	wire _w1112_ ;
	wire _w1113_ ;
	wire _w1114_ ;
	wire _w1115_ ;
	wire _w1116_ ;
	wire _w1117_ ;
	wire _w1118_ ;
	wire _w1119_ ;
	wire _w1120_ ;
	wire _w1121_ ;
	wire _w1122_ ;
	wire _w1123_ ;
	wire _w1124_ ;
	wire _w1125_ ;
	wire _w1126_ ;
	wire _w1127_ ;
	wire _w1128_ ;
	wire _w1129_ ;
	wire _w1130_ ;
	wire _w1131_ ;
	wire _w1132_ ;
	wire _w1133_ ;
	wire _w1134_ ;
	wire _w1135_ ;
	wire _w1136_ ;
	wire _w1137_ ;
	wire _w1138_ ;
	wire _w1139_ ;
	wire _w1140_ ;
	wire _w1141_ ;
	wire _w1142_ ;
	wire _w1143_ ;
	wire _w1144_ ;
	wire _w1145_ ;
	wire _w1146_ ;
	wire _w1147_ ;
	wire _w1148_ ;
	wire _w1149_ ;
	wire _w1150_ ;
	wire _w1151_ ;
	wire _w1152_ ;
	wire _w1153_ ;
	wire _w1154_ ;
	wire _w1155_ ;
	wire _w1156_ ;
	wire _w1157_ ;
	wire _w1158_ ;
	wire _w1159_ ;
	wire _w1160_ ;
	wire _w1161_ ;
	wire _w1162_ ;
	wire _w1163_ ;
	wire _w1164_ ;
	wire _w1165_ ;
	wire _w1166_ ;
	wire _w1167_ ;
	wire _w1168_ ;
	wire _w1169_ ;
	wire _w1170_ ;
	wire _w1171_ ;
	wire _w1172_ ;
	wire _w1173_ ;
	wire _w1174_ ;
	wire _w1175_ ;
	wire _w1176_ ;
	wire _w1177_ ;
	wire _w1178_ ;
	wire _w1179_ ;
	wire _w1180_ ;
	wire _w1181_ ;
	wire _w1182_ ;
	wire _w1183_ ;
	wire _w1184_ ;
	wire _w1185_ ;
	wire _w1186_ ;
	wire _w1187_ ;
	wire _w1188_ ;
	wire _w1189_ ;
	wire _w1190_ ;
	wire _w1191_ ;
	wire _w1192_ ;
	wire _w1193_ ;
	wire _w1194_ ;
	wire _w1195_ ;
	wire _w1196_ ;
	wire _w1197_ ;
	wire _w1198_ ;
	wire _w1199_ ;
	wire _w1200_ ;
	wire _w1201_ ;
	wire _w1202_ ;
	wire _w1203_ ;
	wire _w1204_ ;
	wire _w1205_ ;
	wire _w1206_ ;
	wire _w1207_ ;
	wire _w1208_ ;
	wire _w1209_ ;
	wire _w1210_ ;
	wire _w1211_ ;
	wire _w1212_ ;
	wire _w1213_ ;
	wire _w1214_ ;
	wire _w1215_ ;
	wire _w1216_ ;
	wire _w1217_ ;
	wire _w1218_ ;
	wire _w1219_ ;
	wire _w1220_ ;
	wire _w1221_ ;
	wire _w1222_ ;
	wire _w1223_ ;
	wire _w1224_ ;
	wire _w1225_ ;
	wire _w1226_ ;
	wire _w1227_ ;
	wire _w1228_ ;
	wire _w1229_ ;
	wire _w1230_ ;
	wire _w1231_ ;
	wire _w1232_ ;
	wire _w1233_ ;
	wire _w1234_ ;
	wire _w1235_ ;
	wire _w1236_ ;
	wire _w1237_ ;
	wire _w1238_ ;
	wire _w1239_ ;
	wire _w1240_ ;
	wire _w1241_ ;
	wire _w1242_ ;
	wire _w1243_ ;
	wire _w1244_ ;
	wire _w1245_ ;
	wire _w1246_ ;
	wire _w1247_ ;
	wire _w1248_ ;
	wire _w1249_ ;
	wire _w1250_ ;
	wire _w1251_ ;
	wire _w1252_ ;
	wire _w1253_ ;
	wire _w1254_ ;
	wire _w1255_ ;
	wire _w1256_ ;
	wire _w1257_ ;
	wire _w1258_ ;
	wire _w1259_ ;
	wire _w1260_ ;
	wire _w1261_ ;
	wire _w1262_ ;
	wire _w1263_ ;
	wire _w1264_ ;
	wire _w1265_ ;
	wire _w1266_ ;
	wire _w1267_ ;
	wire _w1268_ ;
	wire _w1269_ ;
	wire _w1270_ ;
	wire _w1271_ ;
	wire _w1272_ ;
	wire _w1273_ ;
	wire _w1274_ ;
	wire _w1275_ ;
	wire _w1276_ ;
	wire _w1277_ ;
	wire _w1278_ ;
	wire _w1279_ ;
	wire _w1280_ ;
	wire _w1281_ ;
	wire _w1282_ ;
	wire _w1283_ ;
	wire _w1284_ ;
	wire _w1285_ ;
	wire _w1286_ ;
	wire _w1287_ ;
	wire _w1288_ ;
	wire _w1289_ ;
	wire _w1290_ ;
	wire _w1291_ ;
	wire _w1292_ ;
	wire _w1293_ ;
	wire _w1294_ ;
	wire _w1295_ ;
	wire _w1296_ ;
	wire _w1297_ ;
	wire _w1298_ ;
	wire _w1299_ ;
	wire _w1300_ ;
	wire _w1301_ ;
	wire _w1302_ ;
	wire _w1303_ ;
	wire _w1304_ ;
	wire _w1305_ ;
	wire _w1306_ ;
	wire _w1307_ ;
	wire _w1308_ ;
	wire _w1309_ ;
	wire _w1310_ ;
	wire _w1311_ ;
	wire _w1312_ ;
	wire _w1313_ ;
	wire _w1314_ ;
	wire _w1315_ ;
	wire _w1316_ ;
	wire _w1317_ ;
	wire _w1318_ ;
	wire _w1319_ ;
	wire _w1320_ ;
	wire _w1321_ ;
	wire _w1322_ ;
	wire _w1323_ ;
	wire _w1324_ ;
	wire _w1325_ ;
	wire _w1326_ ;
	wire _w1327_ ;
	wire _w1328_ ;
	wire _w1329_ ;
	wire _w1330_ ;
	wire _w1331_ ;
	wire _w1332_ ;
	wire _w1333_ ;
	wire _w1334_ ;
	wire _w1335_ ;
	wire _w1336_ ;
	wire _w1337_ ;
	wire _w1338_ ;
	wire _w1339_ ;
	wire _w1340_ ;
	wire _w1341_ ;
	wire _w1342_ ;
	wire _w1343_ ;
	wire _w1344_ ;
	wire _w1345_ ;
	wire _w1346_ ;
	wire _w1347_ ;
	wire _w1348_ ;
	wire _w1349_ ;
	wire _w1350_ ;
	LUT2 #(
		.INIT('h9)
	) name0 (
		\ctrl_reg[4]/NET0131 ,
		\shift_cnt_reg[4]/NET0131 ,
		_w242_
	);
	LUT2 #(
		.INIT('h2)
	) name1 (
		\ctrl_reg[3]/NET0131 ,
		\shift_cnt_reg[3]/NET0131 ,
		_w243_
	);
	LUT2 #(
		.INIT('h4)
	) name2 (
		\ctrl_reg[3]/NET0131 ,
		\shift_cnt_reg[3]/NET0131 ,
		_w244_
	);
	LUT4 #(
		.INIT('h7310)
	) name3 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[1]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_cnt_reg[1]/NET0131 ,
		_w245_
	);
	LUT4 #(
		.INIT('h002b)
	) name4 (
		\ctrl_reg[2]/NET0131 ,
		\shift_cnt_reg[2]/NET0131 ,
		_w245_,
		_w244_,
		_w246_
	);
	LUT4 #(
		.INIT('h0a28)
	) name5 (
		\ctrl_reg[11]/NET0131 ,
		_w243_,
		_w242_,
		_w246_,
		_w247_
	);
	LUT4 #(
		.INIT('h0001)
	) name6 (
		\shift_cnt_reg[0]/NET0131 ,
		\shift_cnt_reg[1]/NET0131 ,
		\shift_cnt_reg[2]/NET0131 ,
		\shift_cnt_reg[3]/NET0131 ,
		_w248_
	);
	LUT3 #(
		.INIT('h14)
	) name7 (
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[4]/NET0131 ,
		_w248_,
		_w249_
	);
	LUT2 #(
		.INIT('h1)
	) name8 (
		_w247_,
		_w249_,
		_w250_
	);
	LUT2 #(
		.INIT('h9)
	) name9 (
		\ctrl_reg[2]/NET0131 ,
		\shift_cnt_reg[2]/NET0131 ,
		_w251_
	);
	LUT4 #(
		.INIT('h5401)
	) name10 (
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_cnt_reg[1]/NET0131 ,
		\shift_cnt_reg[2]/NET0131 ,
		_w252_
	);
	LUT4 #(
		.INIT('h007d)
	) name11 (
		\ctrl_reg[11]/NET0131 ,
		_w251_,
		_w245_,
		_w252_,
		_w253_
	);
	LUT2 #(
		.INIT('h9)
	) name12 (
		\ctrl_reg[3]/NET0131 ,
		\shift_cnt_reg[3]/NET0131 ,
		_w254_
	);
	LUT4 #(
		.INIT('h2bd4)
	) name13 (
		\ctrl_reg[2]/NET0131 ,
		\shift_cnt_reg[2]/NET0131 ,
		_w245_,
		_w254_,
		_w255_
	);
	LUT4 #(
		.INIT('h01fe)
	) name14 (
		\shift_cnt_reg[0]/NET0131 ,
		\shift_cnt_reg[1]/NET0131 ,
		\shift_cnt_reg[2]/NET0131 ,
		\shift_cnt_reg[3]/NET0131 ,
		_w256_
	);
	LUT2 #(
		.INIT('h1)
	) name15 (
		\ctrl_reg[11]/NET0131 ,
		_w256_,
		_w257_
	);
	LUT3 #(
		.INIT('h0d)
	) name16 (
		\ctrl_reg[11]/NET0131 ,
		_w255_,
		_w257_,
		_w258_
	);
	LUT4 #(
		.INIT('hc480)
	) name17 (
		\ctrl_reg[11]/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w259_
	);
	LUT4 #(
		.INIT('h9c63)
	) name18 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[1]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_cnt_reg[1]/NET0131 ,
		_w260_
	);
	LUT3 #(
		.INIT('h41)
	) name19 (
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_cnt_reg[1]/NET0131 ,
		_w261_
	);
	LUT3 #(
		.INIT('h0d)
	) name20 (
		\ctrl_reg[11]/NET0131 ,
		_w260_,
		_w261_,
		_w262_
	);
	LUT4 #(
		.INIT('h004b)
	) name21 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[51]/NET0131 ,
		_w263_
	);
	LUT4 #(
		.INIT('h00b4)
	) name22 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[50]/NET0131 ,
		_w264_
	);
	LUT2 #(
		.INIT('h1)
	) name23 (
		_w263_,
		_w264_,
		_w265_
	);
	LUT4 #(
		.INIT('h004b)
	) name24 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[49]/NET0131 ,
		_w266_
	);
	LUT4 #(
		.INIT('h00b4)
	) name25 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[48]/NET0131 ,
		_w267_
	);
	LUT2 #(
		.INIT('h1)
	) name26 (
		_w266_,
		_w267_,
		_w268_
	);
	LUT3 #(
		.INIT('h1b)
	) name27 (
		_w262_,
		_w265_,
		_w268_,
		_w269_
	);
	LUT4 #(
		.INIT('hfc54)
	) name28 (
		_w259_,
		_w247_,
		_w249_,
		_w269_,
		_w270_
	);
	LUT4 #(
		.INIT('h004b)
	) name29 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[59]/NET0131 ,
		_w271_
	);
	LUT4 #(
		.INIT('h00b4)
	) name30 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[58]/NET0131 ,
		_w272_
	);
	LUT2 #(
		.INIT('h1)
	) name31 (
		_w271_,
		_w272_,
		_w273_
	);
	LUT4 #(
		.INIT('h004b)
	) name32 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[57]/NET0131 ,
		_w274_
	);
	LUT4 #(
		.INIT('h00b4)
	) name33 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[56]/NET0131 ,
		_w275_
	);
	LUT2 #(
		.INIT('h1)
	) name34 (
		_w274_,
		_w275_,
		_w276_
	);
	LUT4 #(
		.INIT('h082a)
	) name35 (
		_w253_,
		_w262_,
		_w276_,
		_w273_,
		_w277_
	);
	LUT4 #(
		.INIT('h004b)
	) name36 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[61]/NET0131 ,
		_w278_
	);
	LUT4 #(
		.INIT('h00b4)
	) name37 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[60]/NET0131 ,
		_w279_
	);
	LUT2 #(
		.INIT('h1)
	) name38 (
		_w278_,
		_w279_,
		_w280_
	);
	LUT4 #(
		.INIT('h004b)
	) name39 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[63]/NET0131 ,
		_w281_
	);
	LUT4 #(
		.INIT('h00b4)
	) name40 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[62]/NET0131 ,
		_w282_
	);
	LUT2 #(
		.INIT('h1)
	) name41 (
		_w281_,
		_w282_,
		_w283_
	);
	LUT4 #(
		.INIT('h0145)
	) name42 (
		_w253_,
		_w262_,
		_w283_,
		_w280_,
		_w284_
	);
	LUT3 #(
		.INIT('h01)
	) name43 (
		_w258_,
		_w284_,
		_w277_,
		_w285_
	);
	LUT4 #(
		.INIT('h3120)
	) name44 (
		\ctrl_reg[11]/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w286_
	);
	LUT4 #(
		.INIT('h004b)
	) name45 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[55]/NET0131 ,
		_w287_
	);
	LUT4 #(
		.INIT('h00b4)
	) name46 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[54]/NET0131 ,
		_w288_
	);
	LUT2 #(
		.INIT('h1)
	) name47 (
		_w287_,
		_w288_,
		_w289_
	);
	LUT4 #(
		.INIT('h004b)
	) name48 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[53]/NET0131 ,
		_w290_
	);
	LUT4 #(
		.INIT('h00b4)
	) name49 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[52]/NET0131 ,
		_w291_
	);
	LUT2 #(
		.INIT('h1)
	) name50 (
		_w290_,
		_w291_,
		_w292_
	);
	LUT3 #(
		.INIT('h1b)
	) name51 (
		_w262_,
		_w289_,
		_w292_,
		_w293_
	);
	LUT2 #(
		.INIT('h2)
	) name52 (
		_w286_,
		_w293_,
		_w294_
	);
	LUT3 #(
		.INIT('h10)
	) name53 (
		_w285_,
		_w294_,
		_w270_,
		_w295_
	);
	LUT4 #(
		.INIT('h004b)
	) name54 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[35]/NET0131 ,
		_w296_
	);
	LUT4 #(
		.INIT('h00b4)
	) name55 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[34]/NET0131 ,
		_w297_
	);
	LUT2 #(
		.INIT('h1)
	) name56 (
		_w296_,
		_w297_,
		_w298_
	);
	LUT4 #(
		.INIT('h004b)
	) name57 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[33]/NET0131 ,
		_w299_
	);
	LUT4 #(
		.INIT('h00b4)
	) name58 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[32]/NET0131 ,
		_w300_
	);
	LUT2 #(
		.INIT('h1)
	) name59 (
		_w299_,
		_w300_,
		_w301_
	);
	LUT3 #(
		.INIT('h1b)
	) name60 (
		_w262_,
		_w298_,
		_w301_,
		_w302_
	);
	LUT4 #(
		.INIT('h004b)
	) name61 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[39]/NET0131 ,
		_w303_
	);
	LUT4 #(
		.INIT('h00b4)
	) name62 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[38]/NET0131 ,
		_w304_
	);
	LUT2 #(
		.INIT('h1)
	) name63 (
		_w303_,
		_w304_,
		_w305_
	);
	LUT4 #(
		.INIT('h004b)
	) name64 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[37]/NET0131 ,
		_w306_
	);
	LUT4 #(
		.INIT('h00b4)
	) name65 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[36]/NET0131 ,
		_w307_
	);
	LUT2 #(
		.INIT('h1)
	) name66 (
		_w306_,
		_w307_,
		_w308_
	);
	LUT3 #(
		.INIT('h1b)
	) name67 (
		_w262_,
		_w305_,
		_w308_,
		_w309_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name68 (
		_w253_,
		_w258_,
		_w302_,
		_w309_,
		_w310_
	);
	LUT4 #(
		.INIT('h004b)
	) name69 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[43]/NET0131 ,
		_w311_
	);
	LUT4 #(
		.INIT('h00b4)
	) name70 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[42]/NET0131 ,
		_w312_
	);
	LUT2 #(
		.INIT('h1)
	) name71 (
		_w311_,
		_w312_,
		_w313_
	);
	LUT4 #(
		.INIT('h004b)
	) name72 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[41]/NET0131 ,
		_w314_
	);
	LUT4 #(
		.INIT('h00b4)
	) name73 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[40]/NET0131 ,
		_w315_
	);
	LUT2 #(
		.INIT('h1)
	) name74 (
		_w314_,
		_w315_,
		_w316_
	);
	LUT4 #(
		.INIT('h082a)
	) name75 (
		_w253_,
		_w262_,
		_w316_,
		_w313_,
		_w317_
	);
	LUT4 #(
		.INIT('h004b)
	) name76 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[45]/NET0131 ,
		_w318_
	);
	LUT4 #(
		.INIT('h00b4)
	) name77 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[44]/NET0131 ,
		_w319_
	);
	LUT2 #(
		.INIT('h1)
	) name78 (
		_w318_,
		_w319_,
		_w320_
	);
	LUT4 #(
		.INIT('h004b)
	) name79 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[47]/NET0131 ,
		_w321_
	);
	LUT4 #(
		.INIT('h00b4)
	) name80 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[46]/NET0131 ,
		_w322_
	);
	LUT2 #(
		.INIT('h1)
	) name81 (
		_w321_,
		_w322_,
		_w323_
	);
	LUT4 #(
		.INIT('h0145)
	) name82 (
		_w253_,
		_w262_,
		_w323_,
		_w320_,
		_w324_
	);
	LUT3 #(
		.INIT('h01)
	) name83 (
		_w258_,
		_w324_,
		_w317_,
		_w325_
	);
	LUT2 #(
		.INIT('h9)
	) name84 (
		\ctrl_reg[5]/NET0131 ,
		\shift_cnt_reg[5]/NET0131 ,
		_w326_
	);
	LUT4 #(
		.INIT('h444d)
	) name85 (
		\ctrl_reg[4]/NET0131 ,
		\shift_cnt_reg[4]/NET0131 ,
		_w243_,
		_w246_,
		_w327_
	);
	LUT4 #(
		.INIT('h4150)
	) name86 (
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[4]/NET0131 ,
		\shift_cnt_reg[5]/NET0131 ,
		_w248_,
		_w328_
	);
	LUT4 #(
		.INIT('h007d)
	) name87 (
		\ctrl_reg[11]/NET0131 ,
		_w326_,
		_w327_,
		_w328_,
		_w329_
	);
	LUT4 #(
		.INIT('h00bf)
	) name88 (
		_w325_,
		_w250_,
		_w310_,
		_w329_,
		_w330_
	);
	LUT2 #(
		.INIT('h4)
	) name89 (
		_w295_,
		_w330_,
		_w331_
	);
	LUT4 #(
		.INIT('h004b)
	) name90 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[19]/NET0131 ,
		_w332_
	);
	LUT4 #(
		.INIT('h00b4)
	) name91 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[18]/NET0131 ,
		_w333_
	);
	LUT2 #(
		.INIT('h1)
	) name92 (
		_w332_,
		_w333_,
		_w334_
	);
	LUT2 #(
		.INIT('h8)
	) name93 (
		_w259_,
		_w334_,
		_w335_
	);
	LUT4 #(
		.INIT('h004b)
	) name94 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[23]/NET0131 ,
		_w336_
	);
	LUT4 #(
		.INIT('h00b4)
	) name95 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[22]/NET0131 ,
		_w337_
	);
	LUT2 #(
		.INIT('h1)
	) name96 (
		_w336_,
		_w337_,
		_w338_
	);
	LUT3 #(
		.INIT('h15)
	) name97 (
		_w262_,
		_w286_,
		_w338_,
		_w339_
	);
	LUT4 #(
		.INIT('h004b)
	) name98 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[17]/NET0131 ,
		_w340_
	);
	LUT4 #(
		.INIT('h00b4)
	) name99 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[16]/NET0131 ,
		_w341_
	);
	LUT2 #(
		.INIT('h1)
	) name100 (
		_w340_,
		_w341_,
		_w342_
	);
	LUT2 #(
		.INIT('h8)
	) name101 (
		_w259_,
		_w342_,
		_w343_
	);
	LUT4 #(
		.INIT('h004b)
	) name102 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[21]/NET0131 ,
		_w344_
	);
	LUT4 #(
		.INIT('h00b4)
	) name103 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[20]/NET0131 ,
		_w345_
	);
	LUT2 #(
		.INIT('h1)
	) name104 (
		_w344_,
		_w345_,
		_w346_
	);
	LUT3 #(
		.INIT('h2a)
	) name105 (
		_w262_,
		_w286_,
		_w346_,
		_w347_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name106 (
		_w335_,
		_w339_,
		_w343_,
		_w347_,
		_w348_
	);
	LUT4 #(
		.INIT('h004b)
	) name107 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[27]/NET0131 ,
		_w349_
	);
	LUT4 #(
		.INIT('h00b4)
	) name108 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[26]/NET0131 ,
		_w350_
	);
	LUT2 #(
		.INIT('h1)
	) name109 (
		_w349_,
		_w350_,
		_w351_
	);
	LUT4 #(
		.INIT('h004b)
	) name110 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[25]/NET0131 ,
		_w352_
	);
	LUT4 #(
		.INIT('h00b4)
	) name111 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[24]/NET0131 ,
		_w353_
	);
	LUT2 #(
		.INIT('h1)
	) name112 (
		_w352_,
		_w353_,
		_w354_
	);
	LUT4 #(
		.INIT('h082a)
	) name113 (
		_w253_,
		_w262_,
		_w354_,
		_w351_,
		_w355_
	);
	LUT4 #(
		.INIT('h004b)
	) name114 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[29]/NET0131 ,
		_w356_
	);
	LUT4 #(
		.INIT('h00b4)
	) name115 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[28]/NET0131 ,
		_w357_
	);
	LUT2 #(
		.INIT('h1)
	) name116 (
		_w356_,
		_w357_,
		_w358_
	);
	LUT4 #(
		.INIT('h004b)
	) name117 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[31]/NET0131 ,
		_w359_
	);
	LUT4 #(
		.INIT('h00b4)
	) name118 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[30]/NET0131 ,
		_w360_
	);
	LUT2 #(
		.INIT('h1)
	) name119 (
		_w359_,
		_w360_,
		_w361_
	);
	LUT4 #(
		.INIT('h0145)
	) name120 (
		_w253_,
		_w262_,
		_w361_,
		_w358_,
		_w362_
	);
	LUT3 #(
		.INIT('h01)
	) name121 (
		_w258_,
		_w362_,
		_w355_,
		_w363_
	);
	LUT2 #(
		.INIT('h1)
	) name122 (
		_w250_,
		_w363_,
		_w364_
	);
	LUT4 #(
		.INIT('h004b)
	) name123 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[3]/NET0131 ,
		_w365_
	);
	LUT4 #(
		.INIT('h00b4)
	) name124 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[2]/NET0131 ,
		_w366_
	);
	LUT2 #(
		.INIT('h1)
	) name125 (
		_w365_,
		_w366_,
		_w367_
	);
	LUT4 #(
		.INIT('h004b)
	) name126 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[1]/NET0131 ,
		_w368_
	);
	LUT4 #(
		.INIT('h00b4)
	) name127 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[0]/NET0131 ,
		_w369_
	);
	LUT2 #(
		.INIT('h1)
	) name128 (
		_w368_,
		_w369_,
		_w370_
	);
	LUT3 #(
		.INIT('h1b)
	) name129 (
		_w262_,
		_w367_,
		_w370_,
		_w371_
	);
	LUT4 #(
		.INIT('h0301)
	) name130 (
		_w259_,
		_w247_,
		_w249_,
		_w371_,
		_w372_
	);
	LUT4 #(
		.INIT('h004b)
	) name131 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[7]/NET0131 ,
		_w373_
	);
	LUT4 #(
		.INIT('h00b4)
	) name132 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[6]/NET0131 ,
		_w374_
	);
	LUT2 #(
		.INIT('h1)
	) name133 (
		_w373_,
		_w374_,
		_w375_
	);
	LUT4 #(
		.INIT('h004b)
	) name134 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[5]/NET0131 ,
		_w376_
	);
	LUT4 #(
		.INIT('h00b4)
	) name135 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[4]/NET0131 ,
		_w377_
	);
	LUT2 #(
		.INIT('h1)
	) name136 (
		_w376_,
		_w377_,
		_w378_
	);
	LUT3 #(
		.INIT('h1b)
	) name137 (
		_w262_,
		_w375_,
		_w378_,
		_w379_
	);
	LUT2 #(
		.INIT('h2)
	) name138 (
		_w286_,
		_w379_,
		_w380_
	);
	LUT4 #(
		.INIT('h004b)
	) name139 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[11]/NET0131 ,
		_w381_
	);
	LUT4 #(
		.INIT('h00b4)
	) name140 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[10]/NET0131 ,
		_w382_
	);
	LUT2 #(
		.INIT('h1)
	) name141 (
		_w381_,
		_w382_,
		_w383_
	);
	LUT4 #(
		.INIT('h004b)
	) name142 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[9]/NET0131 ,
		_w384_
	);
	LUT4 #(
		.INIT('h00b4)
	) name143 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[8]/NET0131 ,
		_w385_
	);
	LUT2 #(
		.INIT('h1)
	) name144 (
		_w384_,
		_w385_,
		_w386_
	);
	LUT4 #(
		.INIT('h082a)
	) name145 (
		_w253_,
		_w262_,
		_w386_,
		_w383_,
		_w387_
	);
	LUT4 #(
		.INIT('h004b)
	) name146 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[13]/NET0131 ,
		_w388_
	);
	LUT4 #(
		.INIT('h00b4)
	) name147 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[12]/NET0131 ,
		_w389_
	);
	LUT2 #(
		.INIT('h1)
	) name148 (
		_w388_,
		_w389_,
		_w390_
	);
	LUT4 #(
		.INIT('h004b)
	) name149 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[15]/NET0131 ,
		_w391_
	);
	LUT4 #(
		.INIT('h00b4)
	) name150 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[14]/NET0131 ,
		_w392_
	);
	LUT2 #(
		.INIT('h1)
	) name151 (
		_w391_,
		_w392_,
		_w393_
	);
	LUT4 #(
		.INIT('h0145)
	) name152 (
		_w253_,
		_w262_,
		_w393_,
		_w390_,
		_w394_
	);
	LUT3 #(
		.INIT('h01)
	) name153 (
		_w258_,
		_w394_,
		_w387_,
		_w395_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name154 (
		_w329_,
		_w380_,
		_w395_,
		_w372_,
		_w396_
	);
	LUT3 #(
		.INIT('hb0)
	) name155 (
		_w348_,
		_w364_,
		_w396_,
		_w397_
	);
	LUT4 #(
		.INIT('h0100)
	) name156 (
		\shift_cnt_reg[4]/NET0131 ,
		\shift_cnt_reg[5]/NET0131 ,
		\shift_cnt_reg[6]/NET0131 ,
		_w248_,
		_w398_
	);
	LUT4 #(
		.INIT('h1e0f)
	) name157 (
		\shift_cnt_reg[4]/NET0131 ,
		\shift_cnt_reg[5]/NET0131 ,
		\shift_cnt_reg[6]/NET0131 ,
		_w248_,
		_w399_
	);
	LUT2 #(
		.INIT('h1)
	) name158 (
		\ctrl_reg[11]/NET0131 ,
		_w399_,
		_w400_
	);
	LUT2 #(
		.INIT('h9)
	) name159 (
		\ctrl_reg[6]/NET0131 ,
		\shift_cnt_reg[6]/NET0131 ,
		_w401_
	);
	LUT4 #(
		.INIT('h2bd4)
	) name160 (
		\ctrl_reg[5]/NET0131 ,
		\shift_cnt_reg[5]/NET0131 ,
		_w327_,
		_w401_,
		_w402_
	);
	LUT3 #(
		.INIT('h31)
	) name161 (
		\ctrl_reg[11]/NET0131 ,
		_w400_,
		_w402_,
		_w403_
	);
	LUT3 #(
		.INIT('he0)
	) name162 (
		_w331_,
		_w397_,
		_w403_,
		_w404_
	);
	LUT4 #(
		.INIT('h004b)
	) name163 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[67]/NET0131 ,
		_w405_
	);
	LUT4 #(
		.INIT('h00b4)
	) name164 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[66]/NET0131 ,
		_w406_
	);
	LUT2 #(
		.INIT('h1)
	) name165 (
		_w405_,
		_w406_,
		_w407_
	);
	LUT4 #(
		.INIT('h004b)
	) name166 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[65]/NET0131 ,
		_w408_
	);
	LUT4 #(
		.INIT('h00b4)
	) name167 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[64]/NET0131 ,
		_w409_
	);
	LUT2 #(
		.INIT('h1)
	) name168 (
		_w408_,
		_w409_,
		_w410_
	);
	LUT3 #(
		.INIT('h1b)
	) name169 (
		_w262_,
		_w407_,
		_w410_,
		_w411_
	);
	LUT4 #(
		.INIT('h0301)
	) name170 (
		_w259_,
		_w247_,
		_w249_,
		_w411_,
		_w412_
	);
	LUT4 #(
		.INIT('h004b)
	) name171 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[71]/NET0131 ,
		_w413_
	);
	LUT4 #(
		.INIT('h00b4)
	) name172 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[70]/NET0131 ,
		_w414_
	);
	LUT2 #(
		.INIT('h1)
	) name173 (
		_w413_,
		_w414_,
		_w415_
	);
	LUT4 #(
		.INIT('h004b)
	) name174 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[69]/NET0131 ,
		_w416_
	);
	LUT4 #(
		.INIT('h00b4)
	) name175 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[68]/NET0131 ,
		_w417_
	);
	LUT2 #(
		.INIT('h1)
	) name176 (
		_w416_,
		_w417_,
		_w418_
	);
	LUT3 #(
		.INIT('h1b)
	) name177 (
		_w262_,
		_w415_,
		_w418_,
		_w419_
	);
	LUT2 #(
		.INIT('h2)
	) name178 (
		_w286_,
		_w419_,
		_w420_
	);
	LUT4 #(
		.INIT('h004b)
	) name179 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[73]/NET0131 ,
		_w421_
	);
	LUT4 #(
		.INIT('h00b4)
	) name180 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[72]/NET0131 ,
		_w422_
	);
	LUT2 #(
		.INIT('h1)
	) name181 (
		_w421_,
		_w422_,
		_w423_
	);
	LUT4 #(
		.INIT('h004b)
	) name182 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[75]/NET0131 ,
		_w424_
	);
	LUT4 #(
		.INIT('h00b4)
	) name183 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[74]/NET0131 ,
		_w425_
	);
	LUT2 #(
		.INIT('h1)
	) name184 (
		_w424_,
		_w425_,
		_w426_
	);
	LUT4 #(
		.INIT('h028a)
	) name185 (
		_w253_,
		_w262_,
		_w426_,
		_w423_,
		_w427_
	);
	LUT4 #(
		.INIT('h004b)
	) name186 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[79]/NET0131 ,
		_w428_
	);
	LUT4 #(
		.INIT('h00b4)
	) name187 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[78]/NET0131 ,
		_w429_
	);
	LUT2 #(
		.INIT('h1)
	) name188 (
		_w428_,
		_w429_,
		_w430_
	);
	LUT4 #(
		.INIT('h004b)
	) name189 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[77]/NET0131 ,
		_w431_
	);
	LUT4 #(
		.INIT('h00b4)
	) name190 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[76]/NET0131 ,
		_w432_
	);
	LUT2 #(
		.INIT('h1)
	) name191 (
		_w431_,
		_w432_,
		_w433_
	);
	LUT4 #(
		.INIT('h0415)
	) name192 (
		_w253_,
		_w262_,
		_w433_,
		_w430_,
		_w434_
	);
	LUT3 #(
		.INIT('h01)
	) name193 (
		_w258_,
		_w434_,
		_w427_,
		_w435_
	);
	LUT3 #(
		.INIT('h10)
	) name194 (
		_w420_,
		_w435_,
		_w412_,
		_w436_
	);
	LUT4 #(
		.INIT('h004b)
	) name195 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[83]/NET0131 ,
		_w437_
	);
	LUT4 #(
		.INIT('h00b4)
	) name196 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[82]/NET0131 ,
		_w438_
	);
	LUT2 #(
		.INIT('h1)
	) name197 (
		_w437_,
		_w438_,
		_w439_
	);
	LUT4 #(
		.INIT('h004b)
	) name198 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[81]/NET0131 ,
		_w440_
	);
	LUT4 #(
		.INIT('h00b4)
	) name199 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[80]/NET0131 ,
		_w441_
	);
	LUT2 #(
		.INIT('h1)
	) name200 (
		_w440_,
		_w441_,
		_w442_
	);
	LUT3 #(
		.INIT('h1b)
	) name201 (
		_w262_,
		_w439_,
		_w442_,
		_w443_
	);
	LUT4 #(
		.INIT('hfc54)
	) name202 (
		_w259_,
		_w247_,
		_w249_,
		_w443_,
		_w444_
	);
	LUT4 #(
		.INIT('h004b)
	) name203 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[87]/NET0131 ,
		_w445_
	);
	LUT4 #(
		.INIT('h00b4)
	) name204 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[86]/NET0131 ,
		_w446_
	);
	LUT2 #(
		.INIT('h1)
	) name205 (
		_w445_,
		_w446_,
		_w447_
	);
	LUT4 #(
		.INIT('h004b)
	) name206 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[85]/NET0131 ,
		_w448_
	);
	LUT4 #(
		.INIT('h00b4)
	) name207 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[84]/NET0131 ,
		_w449_
	);
	LUT2 #(
		.INIT('h1)
	) name208 (
		_w448_,
		_w449_,
		_w450_
	);
	LUT3 #(
		.INIT('h1b)
	) name209 (
		_w262_,
		_w447_,
		_w450_,
		_w451_
	);
	LUT2 #(
		.INIT('h2)
	) name210 (
		_w286_,
		_w451_,
		_w452_
	);
	LUT4 #(
		.INIT('h004b)
	) name211 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[91]/NET0131 ,
		_w453_
	);
	LUT4 #(
		.INIT('h00b4)
	) name212 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[90]/NET0131 ,
		_w454_
	);
	LUT2 #(
		.INIT('h1)
	) name213 (
		_w453_,
		_w454_,
		_w455_
	);
	LUT4 #(
		.INIT('h004b)
	) name214 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[89]/NET0131 ,
		_w456_
	);
	LUT4 #(
		.INIT('h00b4)
	) name215 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[88]/NET0131 ,
		_w457_
	);
	LUT2 #(
		.INIT('h1)
	) name216 (
		_w456_,
		_w457_,
		_w458_
	);
	LUT4 #(
		.INIT('h082a)
	) name217 (
		_w253_,
		_w262_,
		_w458_,
		_w455_,
		_w459_
	);
	LUT4 #(
		.INIT('h004b)
	) name218 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[93]/NET0131 ,
		_w460_
	);
	LUT4 #(
		.INIT('h00b4)
	) name219 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[92]/NET0131 ,
		_w461_
	);
	LUT2 #(
		.INIT('h1)
	) name220 (
		_w460_,
		_w461_,
		_w462_
	);
	LUT4 #(
		.INIT('h004b)
	) name221 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[95]/NET0131 ,
		_w463_
	);
	LUT4 #(
		.INIT('h00b4)
	) name222 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[94]/NET0131 ,
		_w464_
	);
	LUT2 #(
		.INIT('h1)
	) name223 (
		_w463_,
		_w464_,
		_w465_
	);
	LUT4 #(
		.INIT('h0145)
	) name224 (
		_w253_,
		_w262_,
		_w465_,
		_w462_,
		_w466_
	);
	LUT3 #(
		.INIT('h01)
	) name225 (
		_w258_,
		_w466_,
		_w459_,
		_w467_
	);
	LUT3 #(
		.INIT('h10)
	) name226 (
		_w452_,
		_w467_,
		_w444_,
		_w468_
	);
	LUT3 #(
		.INIT('ha8)
	) name227 (
		_w329_,
		_w436_,
		_w468_,
		_w469_
	);
	LUT4 #(
		.INIT('h004b)
	) name228 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[103]/NET0131 ,
		_w470_
	);
	LUT4 #(
		.INIT('h00b4)
	) name229 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[102]/NET0131 ,
		_w471_
	);
	LUT2 #(
		.INIT('h1)
	) name230 (
		_w470_,
		_w471_,
		_w472_
	);
	LUT4 #(
		.INIT('h004b)
	) name231 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[101]/NET0131 ,
		_w473_
	);
	LUT4 #(
		.INIT('h00b4)
	) name232 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[100]/NET0131 ,
		_w474_
	);
	LUT2 #(
		.INIT('h1)
	) name233 (
		_w473_,
		_w474_,
		_w475_
	);
	LUT3 #(
		.INIT('h1b)
	) name234 (
		_w262_,
		_w472_,
		_w475_,
		_w476_
	);
	LUT4 #(
		.INIT('h0301)
	) name235 (
		_w286_,
		_w247_,
		_w249_,
		_w476_,
		_w477_
	);
	LUT4 #(
		.INIT('h004b)
	) name236 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[99]/NET0131 ,
		_w478_
	);
	LUT4 #(
		.INIT('h00b4)
	) name237 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[98]/NET0131 ,
		_w479_
	);
	LUT2 #(
		.INIT('h1)
	) name238 (
		_w478_,
		_w479_,
		_w480_
	);
	LUT4 #(
		.INIT('h004b)
	) name239 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[97]/NET0131 ,
		_w481_
	);
	LUT4 #(
		.INIT('h00b4)
	) name240 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[96]/NET0131 ,
		_w482_
	);
	LUT2 #(
		.INIT('h1)
	) name241 (
		_w481_,
		_w482_,
		_w483_
	);
	LUT3 #(
		.INIT('h1b)
	) name242 (
		_w262_,
		_w480_,
		_w483_,
		_w484_
	);
	LUT2 #(
		.INIT('h2)
	) name243 (
		_w259_,
		_w484_,
		_w485_
	);
	LUT4 #(
		.INIT('h004b)
	) name244 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[107]/NET0131 ,
		_w486_
	);
	LUT4 #(
		.INIT('h00b4)
	) name245 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[106]/NET0131 ,
		_w487_
	);
	LUT2 #(
		.INIT('h1)
	) name246 (
		_w486_,
		_w487_,
		_w488_
	);
	LUT4 #(
		.INIT('h004b)
	) name247 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[105]/NET0131 ,
		_w489_
	);
	LUT4 #(
		.INIT('h00b4)
	) name248 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[104]/NET0131 ,
		_w490_
	);
	LUT2 #(
		.INIT('h1)
	) name249 (
		_w489_,
		_w490_,
		_w491_
	);
	LUT4 #(
		.INIT('h082a)
	) name250 (
		_w253_,
		_w262_,
		_w491_,
		_w488_,
		_w492_
	);
	LUT4 #(
		.INIT('h004b)
	) name251 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[109]/NET0131 ,
		_w493_
	);
	LUT4 #(
		.INIT('h00b4)
	) name252 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[108]/NET0131 ,
		_w494_
	);
	LUT2 #(
		.INIT('h1)
	) name253 (
		_w493_,
		_w494_,
		_w495_
	);
	LUT4 #(
		.INIT('h004b)
	) name254 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[111]/NET0131 ,
		_w496_
	);
	LUT4 #(
		.INIT('h00b4)
	) name255 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[110]/NET0131 ,
		_w497_
	);
	LUT2 #(
		.INIT('h1)
	) name256 (
		_w496_,
		_w497_,
		_w498_
	);
	LUT4 #(
		.INIT('h0145)
	) name257 (
		_w253_,
		_w262_,
		_w498_,
		_w495_,
		_w499_
	);
	LUT3 #(
		.INIT('h01)
	) name258 (
		_w258_,
		_w499_,
		_w492_,
		_w500_
	);
	LUT3 #(
		.INIT('h10)
	) name259 (
		_w485_,
		_w500_,
		_w477_,
		_w501_
	);
	LUT4 #(
		.INIT('h004b)
	) name260 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[119]/NET0131 ,
		_w502_
	);
	LUT4 #(
		.INIT('h00b4)
	) name261 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[118]/NET0131 ,
		_w503_
	);
	LUT2 #(
		.INIT('h1)
	) name262 (
		_w502_,
		_w503_,
		_w504_
	);
	LUT4 #(
		.INIT('h004b)
	) name263 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[117]/NET0131 ,
		_w505_
	);
	LUT4 #(
		.INIT('h00b4)
	) name264 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[116]/NET0131 ,
		_w506_
	);
	LUT2 #(
		.INIT('h1)
	) name265 (
		_w505_,
		_w506_,
		_w507_
	);
	LUT3 #(
		.INIT('h1b)
	) name266 (
		_w262_,
		_w504_,
		_w507_,
		_w508_
	);
	LUT4 #(
		.INIT('hfc54)
	) name267 (
		_w286_,
		_w247_,
		_w249_,
		_w508_,
		_w509_
	);
	LUT4 #(
		.INIT('h004b)
	) name268 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[115]/NET0131 ,
		_w510_
	);
	LUT4 #(
		.INIT('h00b4)
	) name269 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[114]/NET0131 ,
		_w511_
	);
	LUT2 #(
		.INIT('h1)
	) name270 (
		_w510_,
		_w511_,
		_w512_
	);
	LUT4 #(
		.INIT('h004b)
	) name271 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[113]/NET0131 ,
		_w513_
	);
	LUT4 #(
		.INIT('h00b4)
	) name272 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[112]/NET0131 ,
		_w514_
	);
	LUT2 #(
		.INIT('h1)
	) name273 (
		_w513_,
		_w514_,
		_w515_
	);
	LUT3 #(
		.INIT('h1b)
	) name274 (
		_w262_,
		_w512_,
		_w515_,
		_w516_
	);
	LUT2 #(
		.INIT('h2)
	) name275 (
		_w259_,
		_w516_,
		_w517_
	);
	LUT4 #(
		.INIT('h004b)
	) name276 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[123]/NET0131 ,
		_w518_
	);
	LUT4 #(
		.INIT('h00b4)
	) name277 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[122]/NET0131 ,
		_w519_
	);
	LUT2 #(
		.INIT('h1)
	) name278 (
		_w518_,
		_w519_,
		_w520_
	);
	LUT4 #(
		.INIT('h004b)
	) name279 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[121]/NET0131 ,
		_w521_
	);
	LUT4 #(
		.INIT('h00b4)
	) name280 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[120]/NET0131 ,
		_w522_
	);
	LUT2 #(
		.INIT('h1)
	) name281 (
		_w521_,
		_w522_,
		_w523_
	);
	LUT4 #(
		.INIT('h082a)
	) name282 (
		_w253_,
		_w262_,
		_w523_,
		_w520_,
		_w524_
	);
	LUT4 #(
		.INIT('h004b)
	) name283 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[125]/NET0131 ,
		_w525_
	);
	LUT4 #(
		.INIT('h00b4)
	) name284 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[124]/NET0131 ,
		_w526_
	);
	LUT2 #(
		.INIT('h1)
	) name285 (
		_w525_,
		_w526_,
		_w527_
	);
	LUT4 #(
		.INIT('h004b)
	) name286 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[127]/NET0131 ,
		_w528_
	);
	LUT4 #(
		.INIT('h00b4)
	) name287 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_data_reg[126]/NET0131 ,
		_w529_
	);
	LUT2 #(
		.INIT('h1)
	) name288 (
		_w528_,
		_w529_,
		_w530_
	);
	LUT4 #(
		.INIT('h0145)
	) name289 (
		_w253_,
		_w262_,
		_w530_,
		_w527_,
		_w531_
	);
	LUT3 #(
		.INIT('h01)
	) name290 (
		_w258_,
		_w531_,
		_w524_,
		_w532_
	);
	LUT3 #(
		.INIT('h10)
	) name291 (
		_w517_,
		_w532_,
		_w509_,
		_w533_
	);
	LUT4 #(
		.INIT('h2223)
	) name292 (
		_w329_,
		_w403_,
		_w501_,
		_w533_,
		_w534_
	);
	LUT2 #(
		.INIT('h4)
	) name293 (
		_w469_,
		_w534_,
		_w535_
	);
	LUT2 #(
		.INIT('h4)
	) name294 (
		\shift_cnt_reg[7]/NET0131 ,
		_w398_,
		_w536_
	);
	LUT3 #(
		.INIT('hac)
	) name295 (
		\clgen_neg_edge_reg/NET0131 ,
		\clgen_pos_edge_reg/NET0131 ,
		\ctrl_reg[10]/NET0131 ,
		_w537_
	);
	LUT4 #(
		.INIT('h40cc)
	) name296 (
		\shift_cnt_reg[7]/NET0131 ,
		\shift_tip_reg/NET0131 ,
		_w398_,
		_w537_,
		_w538_
	);
	LUT4 #(
		.INIT('haafc)
	) name297 (
		mosi_pad_o_pad,
		_w404_,
		_w535_,
		_w538_,
		_w539_
	);
	LUT2 #(
		.INIT('h1)
	) name298 (
		\clgen_cnt_reg[7]/NET0131 ,
		\clgen_cnt_reg[8]/NET0131 ,
		_w540_
	);
	LUT3 #(
		.INIT('h01)
	) name299 (
		\clgen_cnt_reg[7]/NET0131 ,
		\clgen_cnt_reg[8]/NET0131 ,
		\clgen_cnt_reg[9]/NET0131 ,
		_w541_
	);
	LUT2 #(
		.INIT('h1)
	) name300 (
		\clgen_cnt_reg[10]/NET0131 ,
		\clgen_cnt_reg[11]/NET0131 ,
		_w542_
	);
	LUT3 #(
		.INIT('h01)
	) name301 (
		\clgen_cnt_reg[4]/NET0131 ,
		\clgen_cnt_reg[5]/NET0131 ,
		\clgen_cnt_reg[6]/NET0131 ,
		_w543_
	);
	LUT3 #(
		.INIT('h80)
	) name302 (
		_w541_,
		_w542_,
		_w543_,
		_w544_
	);
	LUT2 #(
		.INIT('h1)
	) name303 (
		\clgen_cnt_reg[13]/NET0131 ,
		\clgen_cnt_reg[14]/NET0131 ,
		_w545_
	);
	LUT4 #(
		.INIT('h0001)
	) name304 (
		\clgen_cnt_reg[12]/NET0131 ,
		\clgen_cnt_reg[15]/NET0131 ,
		\clgen_cnt_reg[2]/NET0131 ,
		\clgen_cnt_reg[3]/NET0131 ,
		_w546_
	);
	LUT2 #(
		.INIT('h1)
	) name305 (
		\clgen_cnt_reg[0]/NET0131 ,
		\clgen_cnt_reg[1]/NET0131 ,
		_w547_
	);
	LUT3 #(
		.INIT('h80)
	) name306 (
		_w545_,
		_w546_,
		_w547_,
		_w548_
	);
	LUT3 #(
		.INIT('h2a)
	) name307 (
		\shift_tip_reg/NET0131 ,
		_w544_,
		_w548_,
		_w549_
	);
	LUT4 #(
		.INIT('h0001)
	) name308 (
		\clgen_cnt_reg[0]/NET0131 ,
		\clgen_cnt_reg[1]/NET0131 ,
		\clgen_cnt_reg[2]/NET0131 ,
		\clgen_cnt_reg[3]/NET0131 ,
		_w550_
	);
	LUT4 #(
		.INIT('h0100)
	) name309 (
		\clgen_cnt_reg[4]/NET0131 ,
		\clgen_cnt_reg[5]/NET0131 ,
		\clgen_cnt_reg[6]/NET0131 ,
		_w550_,
		_w551_
	);
	LUT4 #(
		.INIT('h1000)
	) name310 (
		\clgen_cnt_reg[10]/NET0131 ,
		\clgen_cnt_reg[11]/NET0131 ,
		_w541_,
		_w551_,
		_w552_
	);
	LUT4 #(
		.INIT('h6333)
	) name311 (
		\clgen_cnt_reg[12]/NET0131 ,
		\clgen_cnt_reg[15]/NET0131 ,
		_w545_,
		_w552_,
		_w553_
	);
	LUT3 #(
		.INIT('h2e)
	) name312 (
		\divider_reg[15]/NET0131 ,
		_w549_,
		_w553_,
		_w554_
	);
	LUT4 #(
		.INIT('h6333)
	) name313 (
		\clgen_cnt_reg[10]/NET0131 ,
		\clgen_cnt_reg[11]/NET0131 ,
		_w541_,
		_w551_,
		_w555_
	);
	LUT3 #(
		.INIT('h2e)
	) name314 (
		\divider_reg[11]/NET0131 ,
		_w549_,
		_w555_,
		_w556_
	);
	LUT4 #(
		.INIT('h60c0)
	) name315 (
		\clgen_pos_edge_reg/NET0131 ,
		\shift_cnt_reg[4]/NET0131 ,
		\shift_tip_reg/NET0131 ,
		_w248_,
		_w557_
	);
	LUT2 #(
		.INIT('h2)
	) name316 (
		\ctrl_reg[4]/NET0131 ,
		\shift_tip_reg/NET0131 ,
		_w558_
	);
	LUT2 #(
		.INIT('he)
	) name317 (
		_w557_,
		_w558_,
		_w559_
	);
	LUT2 #(
		.INIT('h9)
	) name318 (
		\clgen_cnt_reg[7]/NET0131 ,
		_w551_,
		_w560_
	);
	LUT3 #(
		.INIT('h2e)
	) name319 (
		\divider_reg[7]/NET0131 ,
		_w549_,
		_w560_,
		_w561_
	);
	LUT4 #(
		.INIT('h5cac)
	) name320 (
		\clgen_cnt_reg[12]/NET0131 ,
		\divider_reg[12]/NET0131 ,
		_w549_,
		_w552_,
		_w562_
	);
	LUT4 #(
		.INIT('hd0f0)
	) name321 (
		\clgen_pos_edge_reg/NET0131 ,
		\shift_cnt_reg[7]/NET0131 ,
		\shift_tip_reg/NET0131 ,
		_w398_,
		_w563_
	);
	LUT4 #(
		.INIT('h9030)
	) name322 (
		\clgen_pos_edge_reg/NET0131 ,
		\shift_cnt_reg[7]/NET0131 ,
		\shift_tip_reg/NET0131 ,
		_w398_,
		_w564_
	);
	LUT3 #(
		.INIT('h01)
	) name323 (
		\ctrl_reg[4]/NET0131 ,
		\ctrl_reg[5]/NET0131 ,
		\ctrl_reg[6]/NET0131 ,
		_w565_
	);
	LUT4 #(
		.INIT('h0001)
	) name324 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[1]/NET0131 ,
		\ctrl_reg[2]/NET0131 ,
		\ctrl_reg[3]/NET0131 ,
		_w566_
	);
	LUT3 #(
		.INIT('h15)
	) name325 (
		\shift_tip_reg/NET0131 ,
		_w565_,
		_w566_,
		_w567_
	);
	LUT2 #(
		.INIT('h1)
	) name326 (
		_w564_,
		_w567_,
		_w568_
	);
	LUT3 #(
		.INIT('h63)
	) name327 (
		\clgen_cnt_reg[7]/NET0131 ,
		\clgen_cnt_reg[8]/NET0131 ,
		_w551_,
		_w569_
	);
	LUT3 #(
		.INIT('h2e)
	) name328 (
		\divider_reg[8]/NET0131 ,
		_w549_,
		_w569_,
		_w570_
	);
	LUT4 #(
		.INIT('h40e0)
	) name329 (
		\clgen_pos_edge_reg/NET0131 ,
		\shift_cnt_reg[3]/NET0131 ,
		\shift_tip_reg/NET0131 ,
		_w256_,
		_w571_
	);
	LUT2 #(
		.INIT('h2)
	) name330 (
		\ctrl_reg[3]/NET0131 ,
		\shift_tip_reg/NET0131 ,
		_w572_
	);
	LUT2 #(
		.INIT('he)
	) name331 (
		_w571_,
		_w572_,
		_w573_
	);
	LUT2 #(
		.INIT('h9)
	) name332 (
		\clgen_cnt_reg[4]/NET0131 ,
		_w550_,
		_w574_
	);
	LUT4 #(
		.INIT('h002a)
	) name333 (
		\shift_tip_reg/NET0131 ,
		_w544_,
		_w548_,
		_w574_,
		_w575_
	);
	LUT4 #(
		.INIT('ha222)
	) name334 (
		\divider_reg[4]/NET0131 ,
		\shift_tip_reg/NET0131 ,
		_w544_,
		_w548_,
		_w576_
	);
	LUT2 #(
		.INIT('he)
	) name335 (
		_w575_,
		_w576_,
		_w577_
	);
	LUT4 #(
		.INIT('h1e0f)
	) name336 (
		\clgen_cnt_reg[12]/NET0131 ,
		\clgen_cnt_reg[13]/NET0131 ,
		\clgen_cnt_reg[14]/NET0131 ,
		_w552_,
		_w578_
	);
	LUT3 #(
		.INIT('h2e)
	) name337 (
		\divider_reg[14]/NET0131 ,
		_w549_,
		_w578_,
		_w579_
	);
	LUT4 #(
		.INIT('h40e0)
	) name338 (
		\clgen_pos_edge_reg/NET0131 ,
		\shift_cnt_reg[6]/NET0131 ,
		\shift_tip_reg/NET0131 ,
		_w399_,
		_w580_
	);
	LUT2 #(
		.INIT('h2)
	) name339 (
		\ctrl_reg[6]/NET0131 ,
		\shift_tip_reg/NET0131 ,
		_w581_
	);
	LUT2 #(
		.INIT('he)
	) name340 (
		_w580_,
		_w581_,
		_w582_
	);
	LUT2 #(
		.INIT('h8)
	) name341 (
		\wb_dat_i[8]_pad ,
		\wb_sel_i[1]_pad ,
		_w583_
	);
	LUT3 #(
		.INIT('h35)
	) name342 (
		\ctrl_reg[8]/NET0131 ,
		\wb_dat_i[8]_pad ,
		\wb_sel_i[1]_pad ,
		_w584_
	);
	LUT3 #(
		.INIT('h40)
	) name343 (
		\wb_adr_i[2]_pad ,
		wb_stb_i_pad,
		wb_we_i_pad,
		_w585_
	);
	LUT3 #(
		.INIT('h40)
	) name344 (
		\shift_tip_reg/NET0131 ,
		\wb_adr_i[4]_pad ,
		wb_cyc_i_pad,
		_w586_
	);
	LUT4 #(
		.INIT('h1000)
	) name345 (
		\shift_tip_reg/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		wb_cyc_i_pad,
		_w587_
	);
	LUT3 #(
		.INIT('h40)
	) name346 (
		_w584_,
		_w585_,
		_w587_,
		_w588_
	);
	LUT4 #(
		.INIT('h2000)
	) name347 (
		\clgen_pos_edge_reg/NET0131 ,
		\shift_cnt_reg[7]/NET0131 ,
		\shift_tip_reg/NET0131 ,
		_w398_,
		_w589_
	);
	LUT3 #(
		.INIT('h2a)
	) name348 (
		\ctrl_reg[8]/NET0131 ,
		_w585_,
		_w587_,
		_w590_
	);
	LUT3 #(
		.INIT('hba)
	) name349 (
		_w588_,
		_w589_,
		_w590_,
		_w591_
	);
	LUT4 #(
		.INIT('h01fe)
	) name350 (
		\clgen_cnt_reg[0]/NET0131 ,
		\clgen_cnt_reg[1]/NET0131 ,
		\clgen_cnt_reg[2]/NET0131 ,
		\clgen_cnt_reg[3]/NET0131 ,
		_w592_
	);
	LUT4 #(
		.INIT('h002a)
	) name351 (
		\shift_tip_reg/NET0131 ,
		_w544_,
		_w548_,
		_w592_,
		_w593_
	);
	LUT4 #(
		.INIT('ha222)
	) name352 (
		\divider_reg[3]/NET0131 ,
		\shift_tip_reg/NET0131 ,
		_w544_,
		_w548_,
		_w594_
	);
	LUT2 #(
		.INIT('he)
	) name353 (
		_w593_,
		_w594_,
		_w595_
	);
	LUT4 #(
		.INIT('h90c0)
	) name354 (
		\clgen_cnt_reg[12]/NET0131 ,
		\clgen_cnt_reg[13]/NET0131 ,
		_w549_,
		_w552_,
		_w596_
	);
	LUT4 #(
		.INIT('ha222)
	) name355 (
		\divider_reg[13]/NET0131 ,
		\shift_tip_reg/NET0131 ,
		_w544_,
		_w548_,
		_w597_
	);
	LUT2 #(
		.INIT('he)
	) name356 (
		_w596_,
		_w597_,
		_w598_
	);
	LUT3 #(
		.INIT('h95)
	) name357 (
		\clgen_cnt_reg[10]/NET0131 ,
		_w541_,
		_w551_,
		_w599_
	);
	LUT3 #(
		.INIT('h2e)
	) name358 (
		\divider_reg[10]/NET0131 ,
		_w549_,
		_w599_,
		_w600_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name359 (
		sclk_pad_o_pad,
		\shift_tip_reg/NET0131 ,
		_w544_,
		_w548_,
		_w601_
	);
	LUT2 #(
		.INIT('h4)
	) name360 (
		sclk_pad_o_pad,
		\shift_tip_reg/NET0131 ,
		_w602_
	);
	LUT3 #(
		.INIT('h80)
	) name361 (
		_w544_,
		_w548_,
		_w602_,
		_w603_
	);
	LUT3 #(
		.INIT('hdc)
	) name362 (
		_w536_,
		_w601_,
		_w603_,
		_w604_
	);
	LUT4 #(
		.INIT('hfd02)
	) name363 (
		\clgen_pos_edge_reg/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_cnt_reg[1]/NET0131 ,
		\shift_cnt_reg[2]/NET0131 ,
		_w605_
	);
	LUT3 #(
		.INIT('he2)
	) name364 (
		\ctrl_reg[2]/NET0131 ,
		\shift_tip_reg/NET0131 ,
		_w605_,
		_w606_
	);
	LUT2 #(
		.INIT('h2)
	) name365 (
		\clgen_cnt_reg[0]/NET0131 ,
		\clgen_cnt_reg[1]/NET0131 ,
		_w607_
	);
	LUT3 #(
		.INIT('h80)
	) name366 (
		_w545_,
		_w546_,
		_w607_,
		_w608_
	);
	LUT3 #(
		.INIT('h2a)
	) name367 (
		sclk_pad_o_pad,
		_w544_,
		_w608_,
		_w609_
	);
	LUT4 #(
		.INIT('h0001)
	) name368 (
		\divider_reg[13]/NET0131 ,
		\divider_reg[14]/NET0131 ,
		\divider_reg[15]/NET0131 ,
		\divider_reg[1]/NET0131 ,
		_w610_
	);
	LUT4 #(
		.INIT('h0001)
	) name369 (
		\divider_reg[0]/NET0131 ,
		\divider_reg[10]/NET0131 ,
		\divider_reg[11]/NET0131 ,
		\divider_reg[12]/NET0131 ,
		_w611_
	);
	LUT4 #(
		.INIT('h0001)
	) name370 (
		\divider_reg[6]/NET0131 ,
		\divider_reg[7]/NET0131 ,
		\divider_reg[8]/NET0131 ,
		\divider_reg[9]/NET0131 ,
		_w612_
	);
	LUT4 #(
		.INIT('h0001)
	) name371 (
		\divider_reg[2]/NET0131 ,
		\divider_reg[3]/NET0131 ,
		\divider_reg[4]/NET0131 ,
		\divider_reg[5]/NET0131 ,
		_w613_
	);
	LUT4 #(
		.INIT('h8000)
	) name372 (
		_w612_,
		_w613_,
		_w610_,
		_w611_,
		_w614_
	);
	LUT3 #(
		.INIT('hc8)
	) name373 (
		sclk_pad_o_pad,
		\shift_tip_reg/NET0131 ,
		_w614_,
		_w615_
	);
	LUT2 #(
		.INIT('h4)
	) name374 (
		_w609_,
		_w615_,
		_w616_
	);
	LUT4 #(
		.INIT('hd2f0)
	) name375 (
		\clgen_pos_edge_reg/NET0131 ,
		\shift_cnt_reg[4]/NET0131 ,
		\shift_cnt_reg[5]/NET0131 ,
		_w248_,
		_w617_
	);
	LUT3 #(
		.INIT('he2)
	) name376 (
		\ctrl_reg[5]/NET0131 ,
		\shift_tip_reg/NET0131 ,
		_w617_,
		_w618_
	);
	LUT2 #(
		.INIT('h2)
	) name377 (
		\ctrl_reg[8]/NET0131 ,
		\shift_tip_reg/NET0131 ,
		_w619_
	);
	LUT2 #(
		.INIT('he)
	) name378 (
		_w563_,
		_w619_,
		_w620_
	);
	LUT3 #(
		.INIT('h31)
	) name379 (
		\ctrl_reg[8]/NET0131 ,
		sclk_pad_o_pad,
		\shift_tip_reg/NET0131 ,
		_w621_
	);
	LUT2 #(
		.INIT('h2)
	) name380 (
		_w614_,
		_w621_,
		_w622_
	);
	LUT3 #(
		.INIT('h80)
	) name381 (
		_w544_,
		_w602_,
		_w608_,
		_w623_
	);
	LUT2 #(
		.INIT('he)
	) name382 (
		_w622_,
		_w623_,
		_w624_
	);
	LUT2 #(
		.INIT('h4)
	) name383 (
		wb_ack_o_pad,
		wb_int_o_pad,
		_w625_
	);
	LUT3 #(
		.INIT('hf8)
	) name384 (
		\ctrl_reg[12]/NET0131 ,
		_w589_,
		_w625_,
		_w626_
	);
	LUT4 #(
		.INIT('ha222)
	) name385 (
		\divider_reg[5]/NET0131 ,
		\shift_tip_reg/NET0131 ,
		_w544_,
		_w548_,
		_w627_
	);
	LUT3 #(
		.INIT('h63)
	) name386 (
		\clgen_cnt_reg[4]/NET0131 ,
		\clgen_cnt_reg[5]/NET0131 ,
		_w550_,
		_w628_
	);
	LUT4 #(
		.INIT('h002a)
	) name387 (
		\shift_tip_reg/NET0131 ,
		_w544_,
		_w548_,
		_w628_,
		_w629_
	);
	LUT2 #(
		.INIT('he)
	) name388 (
		_w627_,
		_w629_,
		_w630_
	);
	LUT4 #(
		.INIT('ha222)
	) name389 (
		\divider_reg[6]/NET0131 ,
		\shift_tip_reg/NET0131 ,
		_w544_,
		_w548_,
		_w631_
	);
	LUT4 #(
		.INIT('h1e0f)
	) name390 (
		\clgen_cnt_reg[4]/NET0131 ,
		\clgen_cnt_reg[5]/NET0131 ,
		\clgen_cnt_reg[6]/NET0131 ,
		_w550_,
		_w632_
	);
	LUT4 #(
		.INIT('h002a)
	) name391 (
		\shift_tip_reg/NET0131 ,
		_w544_,
		_w548_,
		_w632_,
		_w633_
	);
	LUT2 #(
		.INIT('he)
	) name392 (
		_w631_,
		_w633_,
		_w634_
	);
	LUT4 #(
		.INIT('ha222)
	) name393 (
		\divider_reg[0]/NET0131 ,
		\shift_tip_reg/NET0131 ,
		_w544_,
		_w548_,
		_w635_
	);
	LUT4 #(
		.INIT('h0444)
	) name394 (
		\clgen_cnt_reg[0]/NET0131 ,
		\shift_tip_reg/NET0131 ,
		_w544_,
		_w548_,
		_w636_
	);
	LUT2 #(
		.INIT('he)
	) name395 (
		_w635_,
		_w636_,
		_w637_
	);
	LUT3 #(
		.INIT('h95)
	) name396 (
		\clgen_cnt_reg[9]/NET0131 ,
		_w540_,
		_w551_,
		_w638_
	);
	LUT3 #(
		.INIT('h2e)
	) name397 (
		\divider_reg[9]/NET0131 ,
		_w549_,
		_w638_,
		_w639_
	);
	LUT3 #(
		.INIT('h1e)
	) name398 (
		\clgen_cnt_reg[0]/NET0131 ,
		\clgen_cnt_reg[1]/NET0131 ,
		\clgen_cnt_reg[2]/NET0131 ,
		_w640_
	);
	LUT4 #(
		.INIT('h002a)
	) name399 (
		\shift_tip_reg/NET0131 ,
		_w544_,
		_w548_,
		_w640_,
		_w641_
	);
	LUT4 #(
		.INIT('ha222)
	) name400 (
		\divider_reg[2]/NET0131 ,
		\shift_tip_reg/NET0131 ,
		_w544_,
		_w548_,
		_w642_
	);
	LUT2 #(
		.INIT('he)
	) name401 (
		_w641_,
		_w642_,
		_w643_
	);
	LUT4 #(
		.INIT('ha222)
	) name402 (
		\divider_reg[1]/NET0131 ,
		\shift_tip_reg/NET0131 ,
		_w544_,
		_w548_,
		_w644_
	);
	LUT2 #(
		.INIT('h9)
	) name403 (
		\clgen_cnt_reg[0]/NET0131 ,
		\clgen_cnt_reg[1]/NET0131 ,
		_w645_
	);
	LUT4 #(
		.INIT('h2a00)
	) name404 (
		\shift_tip_reg/NET0131 ,
		_w544_,
		_w548_,
		_w645_,
		_w646_
	);
	LUT2 #(
		.INIT('he)
	) name405 (
		_w644_,
		_w646_,
		_w647_
	);
	LUT4 #(
		.INIT('h2d00)
	) name406 (
		\clgen_pos_edge_reg/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_cnt_reg[1]/NET0131 ,
		\shift_tip_reg/NET0131 ,
		_w648_
	);
	LUT2 #(
		.INIT('h1)
	) name407 (
		\ctrl_reg[1]/NET0131 ,
		\shift_tip_reg/NET0131 ,
		_w649_
	);
	LUT2 #(
		.INIT('h1)
	) name408 (
		_w648_,
		_w649_,
		_w650_
	);
	LUT4 #(
		.INIT('h0008)
	) name409 (
		\shift_data_reg[35]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w651_
	);
	LUT4 #(
		.INIT('h0020)
	) name410 (
		\shift_data_reg[67]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w652_
	);
	LUT4 #(
		.INIT('h0002)
	) name411 (
		\shift_data_reg[3]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w653_
	);
	LUT3 #(
		.INIT('h01)
	) name412 (
		_w652_,
		_w653_,
		_w651_,
		_w654_
	);
	LUT4 #(
		.INIT('h0080)
	) name413 (
		\shift_data_reg[99]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w655_
	);
	LUT4 #(
		.INIT('h0200)
	) name414 (
		\ctrl_reg[3]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w656_
	);
	LUT4 #(
		.INIT('h2000)
	) name415 (
		\ss_reg[3]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w657_
	);
	LUT4 #(
		.INIT('h0800)
	) name416 (
		\divider_reg[3]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w658_
	);
	LUT4 #(
		.INIT('h0001)
	) name417 (
		_w655_,
		_w656_,
		_w657_,
		_w658_,
		_w659_
	);
	LUT2 #(
		.INIT('h7)
	) name418 (
		_w654_,
		_w659_,
		_w660_
	);
	LUT4 #(
		.INIT('h0008)
	) name419 (
		\shift_data_reg[39]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w661_
	);
	LUT4 #(
		.INIT('h0020)
	) name420 (
		\shift_data_reg[71]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w662_
	);
	LUT4 #(
		.INIT('h0002)
	) name421 (
		\shift_data_reg[7]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w663_
	);
	LUT3 #(
		.INIT('h01)
	) name422 (
		_w662_,
		_w663_,
		_w661_,
		_w664_
	);
	LUT4 #(
		.INIT('h0080)
	) name423 (
		\shift_data_reg[103]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w665_
	);
	LUT4 #(
		.INIT('h0200)
	) name424 (
		\ctrl_reg[7]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w666_
	);
	LUT4 #(
		.INIT('h2000)
	) name425 (
		\ss_reg[7]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w667_
	);
	LUT4 #(
		.INIT('h0800)
	) name426 (
		\divider_reg[7]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w668_
	);
	LUT4 #(
		.INIT('h0001)
	) name427 (
		_w665_,
		_w666_,
		_w667_,
		_w668_,
		_w669_
	);
	LUT2 #(
		.INIT('h7)
	) name428 (
		_w664_,
		_w669_,
		_w670_
	);
	LUT4 #(
		.INIT('h0008)
	) name429 (
		\shift_data_reg[40]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w671_
	);
	LUT4 #(
		.INIT('h0080)
	) name430 (
		\shift_data_reg[104]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w672_
	);
	LUT2 #(
		.INIT('h1)
	) name431 (
		_w671_,
		_w672_,
		_w673_
	);
	LUT4 #(
		.INIT('h0002)
	) name432 (
		\shift_data_reg[8]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w674_
	);
	LUT4 #(
		.INIT('h0800)
	) name433 (
		\divider_reg[8]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w675_
	);
	LUT4 #(
		.INIT('h0020)
	) name434 (
		\shift_data_reg[72]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w676_
	);
	LUT4 #(
		.INIT('h0200)
	) name435 (
		\ctrl_reg[8]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w677_
	);
	LUT4 #(
		.INIT('h0001)
	) name436 (
		_w674_,
		_w675_,
		_w676_,
		_w677_,
		_w678_
	);
	LUT2 #(
		.INIT('h7)
	) name437 (
		_w673_,
		_w678_,
		_w679_
	);
	LUT4 #(
		.INIT('h0008)
	) name438 (
		\shift_data_reg[41]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w680_
	);
	LUT4 #(
		.INIT('h0080)
	) name439 (
		\shift_data_reg[105]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w681_
	);
	LUT2 #(
		.INIT('h1)
	) name440 (
		_w680_,
		_w681_,
		_w682_
	);
	LUT4 #(
		.INIT('h0002)
	) name441 (
		\shift_data_reg[9]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w683_
	);
	LUT4 #(
		.INIT('h0800)
	) name442 (
		\divider_reg[9]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w684_
	);
	LUT4 #(
		.INIT('h0020)
	) name443 (
		\shift_data_reg[73]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w685_
	);
	LUT4 #(
		.INIT('h0200)
	) name444 (
		\ctrl_reg[9]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w686_
	);
	LUT4 #(
		.INIT('h0001)
	) name445 (
		_w683_,
		_w684_,
		_w685_,
		_w686_,
		_w687_
	);
	LUT2 #(
		.INIT('h7)
	) name446 (
		_w682_,
		_w687_,
		_w688_
	);
	LUT4 #(
		.INIT('h0008)
	) name447 (
		\shift_data_reg[42]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w689_
	);
	LUT4 #(
		.INIT('h0080)
	) name448 (
		\shift_data_reg[106]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w690_
	);
	LUT2 #(
		.INIT('h1)
	) name449 (
		_w689_,
		_w690_,
		_w691_
	);
	LUT4 #(
		.INIT('h0002)
	) name450 (
		\shift_data_reg[10]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w692_
	);
	LUT4 #(
		.INIT('h0800)
	) name451 (
		\divider_reg[10]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w693_
	);
	LUT4 #(
		.INIT('h0020)
	) name452 (
		\shift_data_reg[74]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w694_
	);
	LUT4 #(
		.INIT('h0200)
	) name453 (
		\ctrl_reg[10]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w695_
	);
	LUT4 #(
		.INIT('h0001)
	) name454 (
		_w692_,
		_w693_,
		_w694_,
		_w695_,
		_w696_
	);
	LUT2 #(
		.INIT('h7)
	) name455 (
		_w691_,
		_w696_,
		_w697_
	);
	LUT4 #(
		.INIT('h0008)
	) name456 (
		\shift_data_reg[43]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w698_
	);
	LUT4 #(
		.INIT('h0080)
	) name457 (
		\shift_data_reg[107]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w699_
	);
	LUT2 #(
		.INIT('h1)
	) name458 (
		_w698_,
		_w699_,
		_w700_
	);
	LUT4 #(
		.INIT('h0002)
	) name459 (
		\shift_data_reg[11]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w701_
	);
	LUT4 #(
		.INIT('h0800)
	) name460 (
		\divider_reg[11]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w702_
	);
	LUT4 #(
		.INIT('h0020)
	) name461 (
		\shift_data_reg[75]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w703_
	);
	LUT4 #(
		.INIT('h0200)
	) name462 (
		\ctrl_reg[11]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w704_
	);
	LUT4 #(
		.INIT('h0001)
	) name463 (
		_w701_,
		_w702_,
		_w703_,
		_w704_,
		_w705_
	);
	LUT2 #(
		.INIT('h7)
	) name464 (
		_w700_,
		_w705_,
		_w706_
	);
	LUT4 #(
		.INIT('h0008)
	) name465 (
		\shift_data_reg[44]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w707_
	);
	LUT4 #(
		.INIT('h0080)
	) name466 (
		\shift_data_reg[108]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w708_
	);
	LUT2 #(
		.INIT('h1)
	) name467 (
		_w707_,
		_w708_,
		_w709_
	);
	LUT4 #(
		.INIT('h0002)
	) name468 (
		\shift_data_reg[12]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w710_
	);
	LUT4 #(
		.INIT('h0800)
	) name469 (
		\divider_reg[12]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w711_
	);
	LUT4 #(
		.INIT('h0020)
	) name470 (
		\shift_data_reg[76]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w712_
	);
	LUT4 #(
		.INIT('h0200)
	) name471 (
		\ctrl_reg[12]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w713_
	);
	LUT4 #(
		.INIT('h0001)
	) name472 (
		_w710_,
		_w711_,
		_w712_,
		_w713_,
		_w714_
	);
	LUT2 #(
		.INIT('h7)
	) name473 (
		_w709_,
		_w714_,
		_w715_
	);
	LUT4 #(
		.INIT('h0008)
	) name474 (
		\shift_data_reg[45]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w716_
	);
	LUT4 #(
		.INIT('h0080)
	) name475 (
		\shift_data_reg[109]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w717_
	);
	LUT2 #(
		.INIT('h1)
	) name476 (
		_w716_,
		_w717_,
		_w718_
	);
	LUT4 #(
		.INIT('h0002)
	) name477 (
		\shift_data_reg[13]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w719_
	);
	LUT4 #(
		.INIT('h0800)
	) name478 (
		\divider_reg[13]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w720_
	);
	LUT4 #(
		.INIT('h0020)
	) name479 (
		\shift_data_reg[77]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w721_
	);
	LUT4 #(
		.INIT('h0200)
	) name480 (
		\ctrl_reg[13]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w722_
	);
	LUT4 #(
		.INIT('h0001)
	) name481 (
		_w719_,
		_w720_,
		_w721_,
		_w722_,
		_w723_
	);
	LUT2 #(
		.INIT('h7)
	) name482 (
		_w718_,
		_w723_,
		_w724_
	);
	LUT4 #(
		.INIT('h2000)
	) name483 (
		\ss_reg[2]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w725_
	);
	LUT4 #(
		.INIT('h0800)
	) name484 (
		\divider_reg[2]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w726_
	);
	LUT4 #(
		.INIT('h0080)
	) name485 (
		\shift_data_reg[98]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w727_
	);
	LUT3 #(
		.INIT('h01)
	) name486 (
		_w726_,
		_w727_,
		_w725_,
		_w728_
	);
	LUT4 #(
		.INIT('h0200)
	) name487 (
		\ctrl_reg[2]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w729_
	);
	LUT4 #(
		.INIT('h0002)
	) name488 (
		\shift_data_reg[2]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w730_
	);
	LUT4 #(
		.INIT('h0008)
	) name489 (
		\shift_data_reg[34]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w731_
	);
	LUT4 #(
		.INIT('h0020)
	) name490 (
		\shift_data_reg[66]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w732_
	);
	LUT4 #(
		.INIT('h0001)
	) name491 (
		_w729_,
		_w730_,
		_w731_,
		_w732_,
		_w733_
	);
	LUT2 #(
		.INIT('h7)
	) name492 (
		_w728_,
		_w733_,
		_w734_
	);
	LUT4 #(
		.INIT('h2000)
	) name493 (
		\ss_reg[5]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w735_
	);
	LUT4 #(
		.INIT('h0800)
	) name494 (
		\divider_reg[5]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w736_
	);
	LUT4 #(
		.INIT('h0080)
	) name495 (
		\shift_data_reg[101]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w737_
	);
	LUT3 #(
		.INIT('h01)
	) name496 (
		_w736_,
		_w737_,
		_w735_,
		_w738_
	);
	LUT4 #(
		.INIT('h0200)
	) name497 (
		\ctrl_reg[5]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w739_
	);
	LUT4 #(
		.INIT('h0002)
	) name498 (
		\shift_data_reg[5]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w740_
	);
	LUT4 #(
		.INIT('h0008)
	) name499 (
		\shift_data_reg[37]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w741_
	);
	LUT4 #(
		.INIT('h0020)
	) name500 (
		\shift_data_reg[69]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w742_
	);
	LUT4 #(
		.INIT('h0001)
	) name501 (
		_w739_,
		_w740_,
		_w741_,
		_w742_,
		_w743_
	);
	LUT2 #(
		.INIT('h7)
	) name502 (
		_w738_,
		_w743_,
		_w744_
	);
	LUT4 #(
		.INIT('h2000)
	) name503 (
		\ss_reg[6]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w745_
	);
	LUT4 #(
		.INIT('h0800)
	) name504 (
		\divider_reg[6]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w746_
	);
	LUT4 #(
		.INIT('h0080)
	) name505 (
		\shift_data_reg[102]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w747_
	);
	LUT3 #(
		.INIT('h01)
	) name506 (
		_w746_,
		_w747_,
		_w745_,
		_w748_
	);
	LUT4 #(
		.INIT('h0200)
	) name507 (
		\ctrl_reg[6]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w749_
	);
	LUT4 #(
		.INIT('h0002)
	) name508 (
		\shift_data_reg[6]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w750_
	);
	LUT4 #(
		.INIT('h0008)
	) name509 (
		\shift_data_reg[38]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w751_
	);
	LUT4 #(
		.INIT('h0020)
	) name510 (
		\shift_data_reg[70]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w752_
	);
	LUT4 #(
		.INIT('h0001)
	) name511 (
		_w749_,
		_w750_,
		_w751_,
		_w752_,
		_w753_
	);
	LUT2 #(
		.INIT('h7)
	) name512 (
		_w748_,
		_w753_,
		_w754_
	);
	LUT4 #(
		.INIT('h2000)
	) name513 (
		\ss_reg[4]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w755_
	);
	LUT4 #(
		.INIT('h0800)
	) name514 (
		\divider_reg[4]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w756_
	);
	LUT4 #(
		.INIT('h0080)
	) name515 (
		\shift_data_reg[100]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w757_
	);
	LUT3 #(
		.INIT('h01)
	) name516 (
		_w756_,
		_w757_,
		_w755_,
		_w758_
	);
	LUT4 #(
		.INIT('h0200)
	) name517 (
		\ctrl_reg[4]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w759_
	);
	LUT4 #(
		.INIT('h0002)
	) name518 (
		\shift_data_reg[4]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w760_
	);
	LUT4 #(
		.INIT('h0008)
	) name519 (
		\shift_data_reg[36]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w761_
	);
	LUT4 #(
		.INIT('h0020)
	) name520 (
		\shift_data_reg[68]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w762_
	);
	LUT4 #(
		.INIT('h0001)
	) name521 (
		_w759_,
		_w760_,
		_w761_,
		_w762_,
		_w763_
	);
	LUT2 #(
		.INIT('h7)
	) name522 (
		_w758_,
		_w763_,
		_w764_
	);
	LUT4 #(
		.INIT('h2000)
	) name523 (
		\ss_reg[0]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w765_
	);
	LUT4 #(
		.INIT('h0800)
	) name524 (
		\divider_reg[0]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w766_
	);
	LUT4 #(
		.INIT('h0080)
	) name525 (
		\shift_data_reg[96]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w767_
	);
	LUT3 #(
		.INIT('h01)
	) name526 (
		_w766_,
		_w767_,
		_w765_,
		_w768_
	);
	LUT4 #(
		.INIT('h0200)
	) name527 (
		\ctrl_reg[0]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w769_
	);
	LUT4 #(
		.INIT('h0002)
	) name528 (
		\shift_data_reg[0]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w770_
	);
	LUT4 #(
		.INIT('h0008)
	) name529 (
		\shift_data_reg[32]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w771_
	);
	LUT4 #(
		.INIT('h0020)
	) name530 (
		\shift_data_reg[64]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w772_
	);
	LUT4 #(
		.INIT('h0001)
	) name531 (
		_w769_,
		_w770_,
		_w771_,
		_w772_,
		_w773_
	);
	LUT2 #(
		.INIT('h7)
	) name532 (
		_w768_,
		_w773_,
		_w774_
	);
	LUT4 #(
		.INIT('h2000)
	) name533 (
		\ss_reg[1]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w775_
	);
	LUT4 #(
		.INIT('h0800)
	) name534 (
		\divider_reg[1]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w776_
	);
	LUT4 #(
		.INIT('h0080)
	) name535 (
		\shift_data_reg[97]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w777_
	);
	LUT3 #(
		.INIT('h01)
	) name536 (
		_w776_,
		_w777_,
		_w775_,
		_w778_
	);
	LUT4 #(
		.INIT('h0200)
	) name537 (
		\ctrl_reg[1]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w779_
	);
	LUT4 #(
		.INIT('h0002)
	) name538 (
		\shift_data_reg[1]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w780_
	);
	LUT4 #(
		.INIT('h0008)
	) name539 (
		\shift_data_reg[33]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w781_
	);
	LUT4 #(
		.INIT('h0020)
	) name540 (
		\shift_data_reg[65]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w782_
	);
	LUT4 #(
		.INIT('h0001)
	) name541 (
		_w779_,
		_w780_,
		_w781_,
		_w782_,
		_w783_
	);
	LUT2 #(
		.INIT('h7)
	) name542 (
		_w778_,
		_w783_,
		_w784_
	);
	LUT4 #(
		.INIT('h0020)
	) name543 (
		\shift_data_reg[78]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w785_
	);
	LUT4 #(
		.INIT('h0080)
	) name544 (
		\shift_data_reg[110]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w786_
	);
	LUT2 #(
		.INIT('h1)
	) name545 (
		_w785_,
		_w786_,
		_w787_
	);
	LUT4 #(
		.INIT('h0008)
	) name546 (
		\shift_data_reg[46]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w788_
	);
	LUT4 #(
		.INIT('h0002)
	) name547 (
		\shift_data_reg[14]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w789_
	);
	LUT4 #(
		.INIT('h0800)
	) name548 (
		\divider_reg[14]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w790_
	);
	LUT3 #(
		.INIT('h01)
	) name549 (
		_w789_,
		_w790_,
		_w788_,
		_w791_
	);
	LUT2 #(
		.INIT('h7)
	) name550 (
		_w787_,
		_w791_,
		_w792_
	);
	LUT4 #(
		.INIT('h0020)
	) name551 (
		\shift_data_reg[79]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w793_
	);
	LUT4 #(
		.INIT('h0080)
	) name552 (
		\shift_data_reg[111]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w794_
	);
	LUT2 #(
		.INIT('h1)
	) name553 (
		_w793_,
		_w794_,
		_w795_
	);
	LUT4 #(
		.INIT('h0008)
	) name554 (
		\shift_data_reg[47]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w796_
	);
	LUT4 #(
		.INIT('h0002)
	) name555 (
		\shift_data_reg[15]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w797_
	);
	LUT4 #(
		.INIT('h0800)
	) name556 (
		\divider_reg[15]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w798_
	);
	LUT3 #(
		.INIT('h01)
	) name557 (
		_w797_,
		_w798_,
		_w796_,
		_w799_
	);
	LUT2 #(
		.INIT('h7)
	) name558 (
		_w795_,
		_w799_,
		_w800_
	);
	LUT4 #(
		.INIT('h5acc)
	) name559 (
		\clgen_pos_edge_reg/NET0131 ,
		\ctrl_reg[0]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_tip_reg/NET0131 ,
		_w801_
	);
	LUT4 #(
		.INIT('h8000)
	) name560 (
		\wb_dat_i[0]_pad ,
		\wb_sel_i[0]_pad ,
		_w585_,
		_w587_,
		_w802_
	);
	LUT2 #(
		.INIT('he)
	) name561 (
		\ctrl_reg[0]/NET0131 ,
		_w802_,
		_w803_
	);
	LUT3 #(
		.INIT('h80)
	) name562 (
		\wb_adr_i[2]_pad ,
		wb_stb_i_pad,
		wb_we_i_pad,
		_w804_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name563 (
		\divider_reg[4]/NET0131 ,
		\wb_sel_i[0]_pad ,
		_w587_,
		_w804_,
		_w805_
	);
	LUT2 #(
		.INIT('h8)
	) name564 (
		\wb_dat_i[4]_pad ,
		\wb_sel_i[0]_pad ,
		_w806_
	);
	LUT3 #(
		.INIT('h80)
	) name565 (
		_w587_,
		_w804_,
		_w806_,
		_w807_
	);
	LUT2 #(
		.INIT('he)
	) name566 (
		_w805_,
		_w807_,
		_w808_
	);
	LUT4 #(
		.INIT('h4000)
	) name567 (
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		wb_stb_i_pad,
		wb_we_i_pad,
		_w809_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name568 (
		\ss_reg[4]/NET0131 ,
		\wb_sel_i[0]_pad ,
		_w586_,
		_w809_,
		_w810_
	);
	LUT3 #(
		.INIT('h80)
	) name569 (
		_w586_,
		_w806_,
		_w809_,
		_w811_
	);
	LUT2 #(
		.INIT('he)
	) name570 (
		_w810_,
		_w811_,
		_w812_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name571 (
		\divider_reg[10]/NET0131 ,
		\wb_sel_i[1]_pad ,
		_w587_,
		_w804_,
		_w813_
	);
	LUT2 #(
		.INIT('h8)
	) name572 (
		\wb_dat_i[10]_pad ,
		\wb_sel_i[1]_pad ,
		_w814_
	);
	LUT3 #(
		.INIT('h80)
	) name573 (
		_w587_,
		_w804_,
		_w814_,
		_w815_
	);
	LUT2 #(
		.INIT('he)
	) name574 (
		_w813_,
		_w815_,
		_w816_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name575 (
		\ctrl_reg[7]/NET0131 ,
		\wb_sel_i[0]_pad ,
		_w585_,
		_w587_,
		_w817_
	);
	LUT2 #(
		.INIT('h8)
	) name576 (
		\wb_dat_i[7]_pad ,
		\wb_sel_i[0]_pad ,
		_w818_
	);
	LUT3 #(
		.INIT('h80)
	) name577 (
		_w585_,
		_w587_,
		_w818_,
		_w819_
	);
	LUT2 #(
		.INIT('he)
	) name578 (
		_w817_,
		_w819_,
		_w820_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name579 (
		\divider_reg[13]/NET0131 ,
		\wb_sel_i[1]_pad ,
		_w587_,
		_w804_,
		_w821_
	);
	LUT2 #(
		.INIT('h8)
	) name580 (
		\wb_dat_i[13]_pad ,
		\wb_sel_i[1]_pad ,
		_w822_
	);
	LUT3 #(
		.INIT('h80)
	) name581 (
		_w587_,
		_w804_,
		_w822_,
		_w823_
	);
	LUT2 #(
		.INIT('he)
	) name582 (
		_w821_,
		_w823_,
		_w824_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name583 (
		\divider_reg[5]/NET0131 ,
		\wb_sel_i[0]_pad ,
		_w587_,
		_w804_,
		_w825_
	);
	LUT2 #(
		.INIT('h8)
	) name584 (
		\wb_dat_i[5]_pad ,
		\wb_sel_i[0]_pad ,
		_w826_
	);
	LUT3 #(
		.INIT('h80)
	) name585 (
		_w587_,
		_w804_,
		_w826_,
		_w827_
	);
	LUT2 #(
		.INIT('he)
	) name586 (
		_w825_,
		_w827_,
		_w828_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name587 (
		\ss_reg[7]/NET0131 ,
		\wb_sel_i[0]_pad ,
		_w586_,
		_w809_,
		_w829_
	);
	LUT3 #(
		.INIT('h80)
	) name588 (
		_w586_,
		_w809_,
		_w818_,
		_w830_
	);
	LUT2 #(
		.INIT('he)
	) name589 (
		_w829_,
		_w830_,
		_w831_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name590 (
		\divider_reg[2]/NET0131 ,
		\wb_sel_i[0]_pad ,
		_w587_,
		_w804_,
		_w832_
	);
	LUT2 #(
		.INIT('h8)
	) name591 (
		\wb_dat_i[2]_pad ,
		\wb_sel_i[0]_pad ,
		_w833_
	);
	LUT3 #(
		.INIT('h80)
	) name592 (
		_w587_,
		_w804_,
		_w833_,
		_w834_
	);
	LUT2 #(
		.INIT('he)
	) name593 (
		_w832_,
		_w834_,
		_w835_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name594 (
		\ctrl_reg[10]/NET0131 ,
		\wb_sel_i[1]_pad ,
		_w585_,
		_w587_,
		_w836_
	);
	LUT3 #(
		.INIT('h80)
	) name595 (
		_w585_,
		_w587_,
		_w814_,
		_w837_
	);
	LUT2 #(
		.INIT('he)
	) name596 (
		_w836_,
		_w837_,
		_w838_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name597 (
		\ctrl_reg[11]/NET0131 ,
		\wb_sel_i[1]_pad ,
		_w585_,
		_w587_,
		_w839_
	);
	LUT2 #(
		.INIT('h8)
	) name598 (
		\wb_dat_i[11]_pad ,
		\wb_sel_i[1]_pad ,
		_w840_
	);
	LUT3 #(
		.INIT('h80)
	) name599 (
		_w585_,
		_w587_,
		_w840_,
		_w841_
	);
	LUT2 #(
		.INIT('he)
	) name600 (
		_w839_,
		_w841_,
		_w842_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name601 (
		\divider_reg[14]/NET0131 ,
		\wb_sel_i[1]_pad ,
		_w587_,
		_w804_,
		_w843_
	);
	LUT2 #(
		.INIT('h8)
	) name602 (
		\wb_dat_i[14]_pad ,
		\wb_sel_i[1]_pad ,
		_w844_
	);
	LUT3 #(
		.INIT('h80)
	) name603 (
		_w587_,
		_w804_,
		_w844_,
		_w845_
	);
	LUT2 #(
		.INIT('he)
	) name604 (
		_w843_,
		_w845_,
		_w846_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name605 (
		\ss_reg[6]/NET0131 ,
		\wb_sel_i[0]_pad ,
		_w586_,
		_w809_,
		_w847_
	);
	LUT2 #(
		.INIT('h8)
	) name606 (
		\wb_dat_i[6]_pad ,
		\wb_sel_i[0]_pad ,
		_w848_
	);
	LUT3 #(
		.INIT('h80)
	) name607 (
		_w586_,
		_w809_,
		_w848_,
		_w849_
	);
	LUT2 #(
		.INIT('he)
	) name608 (
		_w847_,
		_w849_,
		_w850_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name609 (
		\ctrl_reg[13]/NET0131 ,
		\wb_sel_i[1]_pad ,
		_w585_,
		_w587_,
		_w851_
	);
	LUT3 #(
		.INIT('h80)
	) name610 (
		_w585_,
		_w587_,
		_w822_,
		_w852_
	);
	LUT2 #(
		.INIT('he)
	) name611 (
		_w851_,
		_w852_,
		_w853_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name612 (
		\ss_reg[5]/NET0131 ,
		\wb_sel_i[0]_pad ,
		_w586_,
		_w809_,
		_w854_
	);
	LUT3 #(
		.INIT('h80)
	) name613 (
		_w586_,
		_w809_,
		_w826_,
		_w855_
	);
	LUT2 #(
		.INIT('he)
	) name614 (
		_w854_,
		_w855_,
		_w856_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name615 (
		\ctrl_reg[1]/NET0131 ,
		\wb_sel_i[0]_pad ,
		_w585_,
		_w587_,
		_w857_
	);
	LUT2 #(
		.INIT('h8)
	) name616 (
		\wb_dat_i[1]_pad ,
		\wb_sel_i[0]_pad ,
		_w858_
	);
	LUT3 #(
		.INIT('h80)
	) name617 (
		_w585_,
		_w587_,
		_w858_,
		_w859_
	);
	LUT2 #(
		.INIT('he)
	) name618 (
		_w857_,
		_w859_,
		_w860_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name619 (
		\ctrl_reg[2]/NET0131 ,
		\wb_sel_i[0]_pad ,
		_w585_,
		_w587_,
		_w861_
	);
	LUT3 #(
		.INIT('h80)
	) name620 (
		_w585_,
		_w587_,
		_w833_,
		_w862_
	);
	LUT2 #(
		.INIT('he)
	) name621 (
		_w861_,
		_w862_,
		_w863_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name622 (
		\ss_reg[2]/NET0131 ,
		\wb_sel_i[0]_pad ,
		_w586_,
		_w809_,
		_w864_
	);
	LUT3 #(
		.INIT('h80)
	) name623 (
		_w586_,
		_w809_,
		_w833_,
		_w865_
	);
	LUT2 #(
		.INIT('he)
	) name624 (
		_w864_,
		_w865_,
		_w866_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name625 (
		\ctrl_reg[3]/NET0131 ,
		\wb_sel_i[0]_pad ,
		_w585_,
		_w587_,
		_w867_
	);
	LUT2 #(
		.INIT('h8)
	) name626 (
		\wb_dat_i[3]_pad ,
		\wb_sel_i[0]_pad ,
		_w868_
	);
	LUT3 #(
		.INIT('h80)
	) name627 (
		_w585_,
		_w587_,
		_w868_,
		_w869_
	);
	LUT2 #(
		.INIT('he)
	) name628 (
		_w867_,
		_w869_,
		_w870_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name629 (
		\ctrl_reg[4]/NET0131 ,
		\wb_sel_i[0]_pad ,
		_w585_,
		_w587_,
		_w871_
	);
	LUT3 #(
		.INIT('h80)
	) name630 (
		_w585_,
		_w587_,
		_w806_,
		_w872_
	);
	LUT2 #(
		.INIT('he)
	) name631 (
		_w871_,
		_w872_,
		_w873_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name632 (
		\ctrl_reg[5]/NET0131 ,
		\wb_sel_i[0]_pad ,
		_w585_,
		_w587_,
		_w874_
	);
	LUT3 #(
		.INIT('h80)
	) name633 (
		_w585_,
		_w587_,
		_w826_,
		_w875_
	);
	LUT2 #(
		.INIT('he)
	) name634 (
		_w874_,
		_w875_,
		_w876_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name635 (
		\ctrl_reg[12]/NET0131 ,
		\wb_sel_i[1]_pad ,
		_w585_,
		_w587_,
		_w877_
	);
	LUT2 #(
		.INIT('h8)
	) name636 (
		\wb_dat_i[12]_pad ,
		\wb_sel_i[1]_pad ,
		_w878_
	);
	LUT3 #(
		.INIT('h80)
	) name637 (
		_w585_,
		_w587_,
		_w878_,
		_w879_
	);
	LUT2 #(
		.INIT('he)
	) name638 (
		_w877_,
		_w879_,
		_w880_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name639 (
		\ctrl_reg[6]/NET0131 ,
		\wb_sel_i[0]_pad ,
		_w585_,
		_w587_,
		_w881_
	);
	LUT3 #(
		.INIT('h80)
	) name640 (
		_w585_,
		_w587_,
		_w848_,
		_w882_
	);
	LUT2 #(
		.INIT('he)
	) name641 (
		_w881_,
		_w882_,
		_w883_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name642 (
		\ctrl_reg[9]/NET0131 ,
		\wb_sel_i[1]_pad ,
		_w585_,
		_w587_,
		_w884_
	);
	LUT2 #(
		.INIT('h8)
	) name643 (
		\wb_dat_i[9]_pad ,
		\wb_sel_i[1]_pad ,
		_w885_
	);
	LUT3 #(
		.INIT('h80)
	) name644 (
		_w585_,
		_w587_,
		_w885_,
		_w886_
	);
	LUT2 #(
		.INIT('he)
	) name645 (
		_w884_,
		_w886_,
		_w887_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name646 (
		\divider_reg[0]/NET0131 ,
		\wb_sel_i[0]_pad ,
		_w587_,
		_w804_,
		_w888_
	);
	LUT2 #(
		.INIT('h8)
	) name647 (
		\wb_dat_i[0]_pad ,
		\wb_sel_i[0]_pad ,
		_w889_
	);
	LUT3 #(
		.INIT('h80)
	) name648 (
		_w587_,
		_w804_,
		_w889_,
		_w890_
	);
	LUT2 #(
		.INIT('he)
	) name649 (
		_w888_,
		_w890_,
		_w891_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name650 (
		\divider_reg[11]/NET0131 ,
		\wb_sel_i[1]_pad ,
		_w587_,
		_w804_,
		_w892_
	);
	LUT3 #(
		.INIT('h80)
	) name651 (
		_w587_,
		_w804_,
		_w840_,
		_w893_
	);
	LUT2 #(
		.INIT('he)
	) name652 (
		_w892_,
		_w893_,
		_w894_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name653 (
		\divider_reg[12]/NET0131 ,
		\wb_sel_i[1]_pad ,
		_w587_,
		_w804_,
		_w895_
	);
	LUT3 #(
		.INIT('h80)
	) name654 (
		_w587_,
		_w804_,
		_w878_,
		_w896_
	);
	LUT2 #(
		.INIT('he)
	) name655 (
		_w895_,
		_w896_,
		_w897_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name656 (
		\divider_reg[15]/NET0131 ,
		\wb_sel_i[1]_pad ,
		_w587_,
		_w804_,
		_w898_
	);
	LUT2 #(
		.INIT('h8)
	) name657 (
		\wb_dat_i[15]_pad ,
		\wb_sel_i[1]_pad ,
		_w899_
	);
	LUT3 #(
		.INIT('h80)
	) name658 (
		_w587_,
		_w804_,
		_w899_,
		_w900_
	);
	LUT2 #(
		.INIT('he)
	) name659 (
		_w898_,
		_w900_,
		_w901_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name660 (
		\divider_reg[8]/NET0131 ,
		\wb_sel_i[1]_pad ,
		_w587_,
		_w804_,
		_w902_
	);
	LUT3 #(
		.INIT('h80)
	) name661 (
		_w583_,
		_w587_,
		_w804_,
		_w903_
	);
	LUT2 #(
		.INIT('he)
	) name662 (
		_w902_,
		_w903_,
		_w904_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name663 (
		\divider_reg[1]/NET0131 ,
		\wb_sel_i[0]_pad ,
		_w587_,
		_w804_,
		_w905_
	);
	LUT3 #(
		.INIT('h80)
	) name664 (
		_w587_,
		_w804_,
		_w858_,
		_w906_
	);
	LUT2 #(
		.INIT('he)
	) name665 (
		_w905_,
		_w906_,
		_w907_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name666 (
		\divider_reg[6]/NET0131 ,
		\wb_sel_i[0]_pad ,
		_w587_,
		_w804_,
		_w908_
	);
	LUT3 #(
		.INIT('h80)
	) name667 (
		_w587_,
		_w804_,
		_w848_,
		_w909_
	);
	LUT2 #(
		.INIT('he)
	) name668 (
		_w908_,
		_w909_,
		_w910_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name669 (
		\divider_reg[3]/NET0131 ,
		\wb_sel_i[0]_pad ,
		_w587_,
		_w804_,
		_w911_
	);
	LUT3 #(
		.INIT('h80)
	) name670 (
		_w587_,
		_w804_,
		_w868_,
		_w912_
	);
	LUT2 #(
		.INIT('he)
	) name671 (
		_w911_,
		_w912_,
		_w913_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name672 (
		\ss_reg[0]/NET0131 ,
		\wb_sel_i[0]_pad ,
		_w586_,
		_w809_,
		_w914_
	);
	LUT3 #(
		.INIT('h80)
	) name673 (
		_w586_,
		_w809_,
		_w889_,
		_w915_
	);
	LUT2 #(
		.INIT('he)
	) name674 (
		_w914_,
		_w915_,
		_w916_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name675 (
		\ss_reg[1]/NET0131 ,
		\wb_sel_i[0]_pad ,
		_w586_,
		_w809_,
		_w917_
	);
	LUT3 #(
		.INIT('h80)
	) name676 (
		_w586_,
		_w809_,
		_w858_,
		_w918_
	);
	LUT2 #(
		.INIT('he)
	) name677 (
		_w917_,
		_w918_,
		_w919_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name678 (
		\ss_reg[3]/NET0131 ,
		\wb_sel_i[0]_pad ,
		_w586_,
		_w809_,
		_w920_
	);
	LUT3 #(
		.INIT('h80)
	) name679 (
		_w586_,
		_w809_,
		_w868_,
		_w921_
	);
	LUT2 #(
		.INIT('he)
	) name680 (
		_w920_,
		_w921_,
		_w922_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name681 (
		\divider_reg[7]/NET0131 ,
		\wb_sel_i[0]_pad ,
		_w587_,
		_w804_,
		_w923_
	);
	LUT3 #(
		.INIT('h80)
	) name682 (
		_w587_,
		_w804_,
		_w818_,
		_w924_
	);
	LUT2 #(
		.INIT('he)
	) name683 (
		_w923_,
		_w924_,
		_w925_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name684 (
		\divider_reg[9]/NET0131 ,
		\wb_sel_i[1]_pad ,
		_w587_,
		_w804_,
		_w926_
	);
	LUT3 #(
		.INIT('h80)
	) name685 (
		_w587_,
		_w804_,
		_w885_,
		_w927_
	);
	LUT2 #(
		.INIT('he)
	) name686 (
		_w926_,
		_w927_,
		_w928_
	);
	LUT4 #(
		.INIT('h0080)
	) name687 (
		\shift_data_reg[120]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w929_
	);
	LUT4 #(
		.INIT('h0008)
	) name688 (
		\shift_data_reg[56]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w930_
	);
	LUT4 #(
		.INIT('h0020)
	) name689 (
		\shift_data_reg[88]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w931_
	);
	LUT4 #(
		.INIT('h0002)
	) name690 (
		\shift_data_reg[24]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w932_
	);
	LUT4 #(
		.INIT('hfffe)
	) name691 (
		_w929_,
		_w930_,
		_w931_,
		_w932_,
		_w933_
	);
	LUT4 #(
		.INIT('h0080)
	) name692 (
		\shift_data_reg[122]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w934_
	);
	LUT4 #(
		.INIT('h0020)
	) name693 (
		\shift_data_reg[90]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w935_
	);
	LUT4 #(
		.INIT('h0002)
	) name694 (
		\shift_data_reg[26]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w936_
	);
	LUT4 #(
		.INIT('h0008)
	) name695 (
		\shift_data_reg[58]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w937_
	);
	LUT4 #(
		.INIT('hfffe)
	) name696 (
		_w934_,
		_w935_,
		_w936_,
		_w937_,
		_w938_
	);
	LUT4 #(
		.INIT('h0080)
	) name697 (
		\shift_data_reg[125]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w939_
	);
	LUT4 #(
		.INIT('h0008)
	) name698 (
		\shift_data_reg[61]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w940_
	);
	LUT4 #(
		.INIT('h0020)
	) name699 (
		\shift_data_reg[93]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w941_
	);
	LUT4 #(
		.INIT('h0002)
	) name700 (
		\shift_data_reg[29]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w942_
	);
	LUT4 #(
		.INIT('hfffe)
	) name701 (
		_w939_,
		_w940_,
		_w941_,
		_w942_,
		_w943_
	);
	LUT4 #(
		.INIT('h0080)
	) name702 (
		\shift_data_reg[126]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w944_
	);
	LUT4 #(
		.INIT('h0008)
	) name703 (
		\shift_data_reg[62]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w945_
	);
	LUT4 #(
		.INIT('h0020)
	) name704 (
		\shift_data_reg[94]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w946_
	);
	LUT4 #(
		.INIT('h0002)
	) name705 (
		\shift_data_reg[30]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w947_
	);
	LUT4 #(
		.INIT('hfffe)
	) name706 (
		_w944_,
		_w945_,
		_w946_,
		_w947_,
		_w948_
	);
	LUT4 #(
		.INIT('h0080)
	) name707 (
		\shift_data_reg[127]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w949_
	);
	LUT4 #(
		.INIT('h0008)
	) name708 (
		\shift_data_reg[63]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w950_
	);
	LUT4 #(
		.INIT('h0020)
	) name709 (
		\shift_data_reg[95]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w951_
	);
	LUT4 #(
		.INIT('h0002)
	) name710 (
		\shift_data_reg[31]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w952_
	);
	LUT4 #(
		.INIT('hfffe)
	) name711 (
		_w949_,
		_w950_,
		_w951_,
		_w952_,
		_w953_
	);
	LUT4 #(
		.INIT('h0080)
	) name712 (
		\shift_data_reg[121]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w954_
	);
	LUT4 #(
		.INIT('h0008)
	) name713 (
		\shift_data_reg[57]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w955_
	);
	LUT4 #(
		.INIT('h0020)
	) name714 (
		\shift_data_reg[89]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w956_
	);
	LUT4 #(
		.INIT('h0002)
	) name715 (
		\shift_data_reg[25]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w957_
	);
	LUT4 #(
		.INIT('hfffe)
	) name716 (
		_w954_,
		_w955_,
		_w956_,
		_w957_,
		_w958_
	);
	LUT4 #(
		.INIT('h0080)
	) name717 (
		\shift_data_reg[123]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w959_
	);
	LUT4 #(
		.INIT('h0008)
	) name718 (
		\shift_data_reg[59]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w960_
	);
	LUT4 #(
		.INIT('h0020)
	) name719 (
		\shift_data_reg[91]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w961_
	);
	LUT4 #(
		.INIT('h0002)
	) name720 (
		\shift_data_reg[27]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w962_
	);
	LUT4 #(
		.INIT('hfffe)
	) name721 (
		_w959_,
		_w960_,
		_w961_,
		_w962_,
		_w963_
	);
	LUT4 #(
		.INIT('h0080)
	) name722 (
		\shift_data_reg[124]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w964_
	);
	LUT4 #(
		.INIT('h0008)
	) name723 (
		\shift_data_reg[60]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w965_
	);
	LUT4 #(
		.INIT('h0020)
	) name724 (
		\shift_data_reg[92]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w966_
	);
	LUT4 #(
		.INIT('h0002)
	) name725 (
		\shift_data_reg[28]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w967_
	);
	LUT4 #(
		.INIT('hfffe)
	) name726 (
		_w964_,
		_w965_,
		_w966_,
		_w967_,
		_w968_
	);
	LUT4 #(
		.INIT('h0080)
	) name727 (
		\shift_data_reg[114]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w969_
	);
	LUT4 #(
		.INIT('h0008)
	) name728 (
		\shift_data_reg[50]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w970_
	);
	LUT4 #(
		.INIT('h0020)
	) name729 (
		\shift_data_reg[82]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w971_
	);
	LUT4 #(
		.INIT('h0002)
	) name730 (
		\shift_data_reg[18]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w972_
	);
	LUT4 #(
		.INIT('hfffe)
	) name731 (
		_w969_,
		_w970_,
		_w971_,
		_w972_,
		_w973_
	);
	LUT4 #(
		.INIT('h0080)
	) name732 (
		\shift_data_reg[116]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w974_
	);
	LUT4 #(
		.INIT('h0008)
	) name733 (
		\shift_data_reg[52]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w975_
	);
	LUT4 #(
		.INIT('h0020)
	) name734 (
		\shift_data_reg[84]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w976_
	);
	LUT4 #(
		.INIT('h0002)
	) name735 (
		\shift_data_reg[20]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w977_
	);
	LUT4 #(
		.INIT('hfffe)
	) name736 (
		_w974_,
		_w975_,
		_w976_,
		_w977_,
		_w978_
	);
	LUT4 #(
		.INIT('h0080)
	) name737 (
		\shift_data_reg[119]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w979_
	);
	LUT4 #(
		.INIT('h0008)
	) name738 (
		\shift_data_reg[55]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w980_
	);
	LUT4 #(
		.INIT('h0020)
	) name739 (
		\shift_data_reg[87]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w981_
	);
	LUT4 #(
		.INIT('h0002)
	) name740 (
		\shift_data_reg[23]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w982_
	);
	LUT4 #(
		.INIT('hfffe)
	) name741 (
		_w979_,
		_w980_,
		_w981_,
		_w982_,
		_w983_
	);
	LUT4 #(
		.INIT('h0002)
	) name742 (
		\shift_data_reg[16]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w984_
	);
	LUT4 #(
		.INIT('h0020)
	) name743 (
		\shift_data_reg[80]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w985_
	);
	LUT4 #(
		.INIT('h0008)
	) name744 (
		\shift_data_reg[48]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w986_
	);
	LUT4 #(
		.INIT('h0080)
	) name745 (
		\shift_data_reg[112]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w987_
	);
	LUT4 #(
		.INIT('hfffe)
	) name746 (
		_w984_,
		_w985_,
		_w986_,
		_w987_,
		_w988_
	);
	LUT4 #(
		.INIT('h0002)
	) name747 (
		\shift_data_reg[17]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w989_
	);
	LUT4 #(
		.INIT('h0020)
	) name748 (
		\shift_data_reg[81]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w990_
	);
	LUT4 #(
		.INIT('h0008)
	) name749 (
		\shift_data_reg[49]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w991_
	);
	LUT4 #(
		.INIT('h0080)
	) name750 (
		\shift_data_reg[113]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w992_
	);
	LUT4 #(
		.INIT('hfffe)
	) name751 (
		_w989_,
		_w990_,
		_w991_,
		_w992_,
		_w993_
	);
	LUT4 #(
		.INIT('h0002)
	) name752 (
		\shift_data_reg[19]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w994_
	);
	LUT4 #(
		.INIT('h0020)
	) name753 (
		\shift_data_reg[83]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w995_
	);
	LUT4 #(
		.INIT('h0008)
	) name754 (
		\shift_data_reg[51]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w996_
	);
	LUT4 #(
		.INIT('h0080)
	) name755 (
		\shift_data_reg[115]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w997_
	);
	LUT4 #(
		.INIT('hfffe)
	) name756 (
		_w994_,
		_w995_,
		_w996_,
		_w997_,
		_w998_
	);
	LUT4 #(
		.INIT('h0080)
	) name757 (
		\shift_data_reg[117]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w999_
	);
	LUT4 #(
		.INIT('h0008)
	) name758 (
		\shift_data_reg[53]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w1000_
	);
	LUT4 #(
		.INIT('h0020)
	) name759 (
		\shift_data_reg[85]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w1001_
	);
	LUT4 #(
		.INIT('h0002)
	) name760 (
		\shift_data_reg[21]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w1002_
	);
	LUT4 #(
		.INIT('hfffe)
	) name761 (
		_w999_,
		_w1000_,
		_w1001_,
		_w1002_,
		_w1003_
	);
	LUT4 #(
		.INIT('h0002)
	) name762 (
		\shift_data_reg[22]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w1004_
	);
	LUT4 #(
		.INIT('h0020)
	) name763 (
		\shift_data_reg[86]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w1005_
	);
	LUT4 #(
		.INIT('h0008)
	) name764 (
		\shift_data_reg[54]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w1006_
	);
	LUT4 #(
		.INIT('h0080)
	) name765 (
		\shift_data_reg[118]/NET0131 ,
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w1007_
	);
	LUT4 #(
		.INIT('hfffe)
	) name766 (
		_w1004_,
		_w1005_,
		_w1006_,
		_w1007_,
		_w1008_
	);
	LUT3 #(
		.INIT('h40)
	) name767 (
		wb_ack_o_pad,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w1009_
	);
	LUT4 #(
		.INIT('h5401)
	) name768 (
		\ctrl_reg[11]/NET0131 ,
		\ctrl_reg[9]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_cnt_reg[1]/NET0131 ,
		_w1010_
	);
	LUT3 #(
		.INIT('h14)
	) name769 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[9]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		_w1011_
	);
	LUT3 #(
		.INIT('h78)
	) name770 (
		\ctrl_reg[9]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_cnt_reg[1]/NET0131 ,
		_w1012_
	);
	LUT4 #(
		.INIT('h6a95)
	) name771 (
		\ctrl_reg[1]/NET0131 ,
		\ctrl_reg[9]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_cnt_reg[1]/NET0131 ,
		_w1013_
	);
	LUT4 #(
		.INIT('h1331)
	) name772 (
		\ctrl_reg[11]/NET0131 ,
		_w1010_,
		_w1011_,
		_w1013_,
		_w1014_
	);
	LUT4 #(
		.INIT('h4bb4)
	) name773 (
		\ctrl_reg[0]/NET0131 ,
		\ctrl_reg[11]/NET0131 ,
		\ctrl_reg[9]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		_w1015_
	);
	LUT2 #(
		.INIT('h1)
	) name774 (
		_w1014_,
		_w1015_,
		_w1016_
	);
	LUT3 #(
		.INIT('hd4)
	) name775 (
		\ctrl_reg[1]/NET0131 ,
		_w1011_,
		_w1012_,
		_w1017_
	);
	LUT4 #(
		.INIT('h8000)
	) name776 (
		\ctrl_reg[9]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_cnt_reg[1]/NET0131 ,
		\shift_cnt_reg[2]/NET0131 ,
		_w1018_
	);
	LUT4 #(
		.INIT('h7f80)
	) name777 (
		\ctrl_reg[9]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_cnt_reg[1]/NET0131 ,
		\shift_cnt_reg[2]/NET0131 ,
		_w1019_
	);
	LUT2 #(
		.INIT('h9)
	) name778 (
		\ctrl_reg[2]/NET0131 ,
		_w1019_,
		_w1020_
	);
	LUT4 #(
		.INIT('h5401)
	) name779 (
		\ctrl_reg[9]/NET0131 ,
		\shift_cnt_reg[0]/NET0131 ,
		\shift_cnt_reg[1]/NET0131 ,
		\shift_cnt_reg[2]/NET0131 ,
		_w1021_
	);
	LUT3 #(
		.INIT('h15)
	) name780 (
		\ctrl_reg[11]/NET0131 ,
		\ctrl_reg[9]/NET0131 ,
		\shift_cnt_reg[2]/NET0131 ,
		_w1022_
	);
	LUT2 #(
		.INIT('h4)
	) name781 (
		_w1021_,
		_w1022_,
		_w1023_
	);
	LUT4 #(
		.INIT('h00d7)
	) name782 (
		\ctrl_reg[11]/NET0131 ,
		_w1017_,
		_w1020_,
		_w1023_,
		_w1024_
	);
	LUT2 #(
		.INIT('h8)
	) name783 (
		_w1016_,
		_w1024_,
		_w1025_
	);
	LUT3 #(
		.INIT('h51)
	) name784 (
		\ctrl_reg[11]/NET0131 ,
		\ctrl_reg[9]/NET0131 ,
		\shift_cnt_reg[3]/NET0131 ,
		_w1026_
	);
	LUT3 #(
		.INIT('hb0)
	) name785 (
		\ctrl_reg[9]/NET0131 ,
		_w256_,
		_w1026_,
		_w1027_
	);
	LUT3 #(
		.INIT('hd4)
	) name786 (
		\ctrl_reg[2]/NET0131 ,
		_w1017_,
		_w1019_,
		_w1028_
	);
	LUT3 #(
		.INIT('h14)
	) name787 (
		\ctrl_reg[3]/NET0131 ,
		\shift_cnt_reg[3]/NET0131 ,
		_w1018_,
		_w1029_
	);
	LUT3 #(
		.INIT('h82)
	) name788 (
		\ctrl_reg[3]/NET0131 ,
		\shift_cnt_reg[3]/NET0131 ,
		_w1018_,
		_w1030_
	);
	LUT3 #(
		.INIT('h69)
	) name789 (
		\ctrl_reg[3]/NET0131 ,
		\shift_cnt_reg[3]/NET0131 ,
		_w1018_,
		_w1031_
	);
	LUT4 #(
		.INIT('h1331)
	) name790 (
		\ctrl_reg[11]/NET0131 ,
		_w1027_,
		_w1028_,
		_w1031_,
		_w1032_
	);
	LUT2 #(
		.INIT('h8)
	) name791 (
		_w1025_,
		_w1032_,
		_w1033_
	);
	LUT4 #(
		.INIT('h1450)
	) name792 (
		\ctrl_reg[4]/NET0131 ,
		\shift_cnt_reg[3]/NET0131 ,
		\shift_cnt_reg[4]/NET0131 ,
		_w1018_,
		_w1034_
	);
	LUT4 #(
		.INIT('h002b)
	) name793 (
		\ctrl_reg[2]/NET0131 ,
		_w1017_,
		_w1019_,
		_w1029_,
		_w1035_
	);
	LUT4 #(
		.INIT('h820a)
	) name794 (
		\ctrl_reg[4]/NET0131 ,
		\shift_cnt_reg[3]/NET0131 ,
		\shift_cnt_reg[4]/NET0131 ,
		_w1018_,
		_w1036_
	);
	LUT2 #(
		.INIT('h1)
	) name795 (
		_w1030_,
		_w1036_,
		_w1037_
	);
	LUT3 #(
		.INIT('h10)
	) name796 (
		_w1034_,
		_w1035_,
		_w1037_,
		_w1038_
	);
	LUT4 #(
		.INIT('h69a5)
	) name797 (
		\ctrl_reg[4]/NET0131 ,
		\shift_cnt_reg[3]/NET0131 ,
		\shift_cnt_reg[4]/NET0131 ,
		_w1018_,
		_w1039_
	);
	LUT4 #(
		.INIT('ha0a2)
	) name798 (
		\ctrl_reg[11]/NET0131 ,
		_w1030_,
		_w1039_,
		_w1035_,
		_w1040_
	);
	LUT4 #(
		.INIT('h1405)
	) name799 (
		\ctrl_reg[11]/NET0131 ,
		\ctrl_reg[9]/NET0131 ,
		\shift_cnt_reg[4]/NET0131 ,
		_w248_,
		_w1041_
	);
	LUT3 #(
		.INIT('h0b)
	) name800 (
		_w1038_,
		_w1040_,
		_w1041_,
		_w1042_
	);
	LUT4 #(
		.INIT('h8000)
	) name801 (
		\shift_cnt_reg[3]/NET0131 ,
		\shift_cnt_reg[4]/NET0131 ,
		\shift_cnt_reg[5]/NET0131 ,
		_w1018_,
		_w1043_
	);
	LUT4 #(
		.INIT('h78f0)
	) name802 (
		\shift_cnt_reg[3]/NET0131 ,
		\shift_cnt_reg[4]/NET0131 ,
		\shift_cnt_reg[5]/NET0131 ,
		_w1018_,
		_w1044_
	);
	LUT2 #(
		.INIT('h2)
	) name803 (
		\ctrl_reg[5]/NET0131 ,
		_w1044_,
		_w1045_
	);
	LUT3 #(
		.INIT('h45)
	) name804 (
		_w1034_,
		_w1035_,
		_w1037_,
		_w1046_
	);
	LUT2 #(
		.INIT('h4)
	) name805 (
		\ctrl_reg[5]/NET0131 ,
		_w1044_,
		_w1047_
	);
	LUT4 #(
		.INIT('h0045)
	) name806 (
		_w1034_,
		_w1035_,
		_w1037_,
		_w1047_,
		_w1048_
	);
	LUT4 #(
		.INIT('h2882)
	) name807 (
		\ctrl_reg[11]/NET0131 ,
		\ctrl_reg[5]/NET0131 ,
		_w1046_,
		_w1044_,
		_w1049_
	);
	LUT4 #(
		.INIT('h1405)
	) name808 (
		\ctrl_reg[9]/NET0131 ,
		\shift_cnt_reg[4]/NET0131 ,
		\shift_cnt_reg[5]/NET0131 ,
		_w248_,
		_w1050_
	);
	LUT3 #(
		.INIT('h51)
	) name809 (
		\ctrl_reg[11]/NET0131 ,
		\ctrl_reg[9]/NET0131 ,
		\shift_cnt_reg[5]/NET0131 ,
		_w1051_
	);
	LUT2 #(
		.INIT('h4)
	) name810 (
		_w1050_,
		_w1051_,
		_w1052_
	);
	LUT2 #(
		.INIT('h1)
	) name811 (
		_w1049_,
		_w1052_,
		_w1053_
	);
	LUT3 #(
		.INIT('ha8)
	) name812 (
		_w1042_,
		_w1049_,
		_w1052_,
		_w1054_
	);
	LUT2 #(
		.INIT('h1)
	) name813 (
		\shift_tip_reg/NET0131 ,
		\wb_adr_i[4]_pad ,
		_w1055_
	);
	LUT2 #(
		.INIT('h8)
	) name814 (
		\wb_adr_i[3]_pad ,
		wb_cyc_i_pad,
		_w1056_
	);
	LUT4 #(
		.INIT('h0400)
	) name815 (
		\shift_tip_reg/NET0131 ,
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		wb_cyc_i_pad,
		_w1057_
	);
	LUT2 #(
		.INIT('h8)
	) name816 (
		_w585_,
		_w1057_,
		_w1058_
	);
	LUT2 #(
		.INIT('h8)
	) name817 (
		_w804_,
		_w1057_,
		_w1059_
	);
	LUT3 #(
		.INIT('h1f)
	) name818 (
		_w585_,
		_w804_,
		_w1057_,
		_w1060_
	);
	LUT2 #(
		.INIT('h6)
	) name819 (
		_w401_,
		_w1043_,
		_w1061_
	);
	LUT4 #(
		.INIT('h02a8)
	) name820 (
		\ctrl_reg[11]/NET0131 ,
		_w1045_,
		_w1048_,
		_w1061_,
		_w1062_
	);
	LUT3 #(
		.INIT('h51)
	) name821 (
		\ctrl_reg[11]/NET0131 ,
		\ctrl_reg[9]/NET0131 ,
		\shift_cnt_reg[6]/NET0131 ,
		_w1063_
	);
	LUT3 #(
		.INIT('hb0)
	) name822 (
		\ctrl_reg[9]/NET0131 ,
		_w399_,
		_w1063_,
		_w1064_
	);
	LUT2 #(
		.INIT('h1)
	) name823 (
		_w1062_,
		_w1064_,
		_w1065_
	);
	LUT3 #(
		.INIT('h02)
	) name824 (
		_w1060_,
		_w1062_,
		_w1064_,
		_w1066_
	);
	LUT3 #(
		.INIT('h80)
	) name825 (
		_w1033_,
		_w1054_,
		_w1066_,
		_w1067_
	);
	LUT3 #(
		.INIT('hac)
	) name826 (
		\shift_data_reg[16]/NET0131 ,
		\shift_data_reg[17]/NET0131 ,
		_w1015_,
		_w1068_
	);
	LUT2 #(
		.INIT('h8)
	) name827 (
		_w1014_,
		_w1068_,
		_w1069_
	);
	LUT3 #(
		.INIT('hac)
	) name828 (
		\shift_data_reg[18]/NET0131 ,
		\shift_data_reg[19]/NET0131 ,
		_w1015_,
		_w1070_
	);
	LUT2 #(
		.INIT('h4)
	) name829 (
		_w1014_,
		_w1070_,
		_w1071_
	);
	LUT3 #(
		.INIT('h01)
	) name830 (
		_w1024_,
		_w1071_,
		_w1069_,
		_w1072_
	);
	LUT3 #(
		.INIT('hac)
	) name831 (
		\shift_data_reg[22]/NET0131 ,
		\shift_data_reg[23]/NET0131 ,
		_w1015_,
		_w1073_
	);
	LUT2 #(
		.INIT('h4)
	) name832 (
		_w1014_,
		_w1073_,
		_w1074_
	);
	LUT3 #(
		.INIT('hac)
	) name833 (
		\shift_data_reg[20]/NET0131 ,
		\shift_data_reg[21]/NET0131 ,
		_w1015_,
		_w1075_
	);
	LUT2 #(
		.INIT('h8)
	) name834 (
		_w1014_,
		_w1075_,
		_w1076_
	);
	LUT3 #(
		.INIT('h02)
	) name835 (
		_w1024_,
		_w1076_,
		_w1074_,
		_w1077_
	);
	LUT3 #(
		.INIT('h02)
	) name836 (
		_w1032_,
		_w1077_,
		_w1072_,
		_w1078_
	);
	LUT3 #(
		.INIT('hac)
	) name837 (
		\shift_data_reg[24]/NET0131 ,
		\shift_data_reg[25]/NET0131 ,
		_w1015_,
		_w1079_
	);
	LUT2 #(
		.INIT('h8)
	) name838 (
		_w1014_,
		_w1079_,
		_w1080_
	);
	LUT3 #(
		.INIT('hac)
	) name839 (
		\shift_data_reg[26]/NET0131 ,
		\shift_data_reg[27]/NET0131 ,
		_w1015_,
		_w1081_
	);
	LUT2 #(
		.INIT('h4)
	) name840 (
		_w1014_,
		_w1081_,
		_w1082_
	);
	LUT3 #(
		.INIT('h01)
	) name841 (
		_w1024_,
		_w1082_,
		_w1080_,
		_w1083_
	);
	LUT3 #(
		.INIT('hac)
	) name842 (
		\shift_data_reg[30]/NET0131 ,
		\shift_data_reg[31]/NET0131 ,
		_w1015_,
		_w1084_
	);
	LUT2 #(
		.INIT('h4)
	) name843 (
		_w1014_,
		_w1084_,
		_w1085_
	);
	LUT3 #(
		.INIT('hac)
	) name844 (
		\shift_data_reg[28]/NET0131 ,
		\shift_data_reg[29]/NET0131 ,
		_w1015_,
		_w1086_
	);
	LUT2 #(
		.INIT('h8)
	) name845 (
		_w1014_,
		_w1086_,
		_w1087_
	);
	LUT3 #(
		.INIT('h02)
	) name846 (
		_w1024_,
		_w1087_,
		_w1085_,
		_w1088_
	);
	LUT3 #(
		.INIT('h01)
	) name847 (
		_w1032_,
		_w1088_,
		_w1083_,
		_w1089_
	);
	LUT3 #(
		.INIT('ha8)
	) name848 (
		_w1042_,
		_w1078_,
		_w1089_,
		_w1090_
	);
	LUT3 #(
		.INIT('hac)
	) name849 (
		\shift_data_reg[8]/NET0131 ,
		\shift_data_reg[9]/NET0131 ,
		_w1015_,
		_w1091_
	);
	LUT2 #(
		.INIT('h8)
	) name850 (
		_w1014_,
		_w1091_,
		_w1092_
	);
	LUT3 #(
		.INIT('hac)
	) name851 (
		\shift_data_reg[10]/NET0131 ,
		\shift_data_reg[11]/NET0131 ,
		_w1015_,
		_w1093_
	);
	LUT2 #(
		.INIT('h4)
	) name852 (
		_w1014_,
		_w1093_,
		_w1094_
	);
	LUT3 #(
		.INIT('h01)
	) name853 (
		_w1024_,
		_w1094_,
		_w1092_,
		_w1095_
	);
	LUT3 #(
		.INIT('hac)
	) name854 (
		\shift_data_reg[14]/NET0131 ,
		\shift_data_reg[15]/NET0131 ,
		_w1015_,
		_w1096_
	);
	LUT2 #(
		.INIT('h4)
	) name855 (
		_w1014_,
		_w1096_,
		_w1097_
	);
	LUT3 #(
		.INIT('hac)
	) name856 (
		\shift_data_reg[12]/NET0131 ,
		\shift_data_reg[13]/NET0131 ,
		_w1015_,
		_w1098_
	);
	LUT2 #(
		.INIT('h8)
	) name857 (
		_w1014_,
		_w1098_,
		_w1099_
	);
	LUT3 #(
		.INIT('h02)
	) name858 (
		_w1024_,
		_w1099_,
		_w1097_,
		_w1100_
	);
	LUT3 #(
		.INIT('h01)
	) name859 (
		_w1032_,
		_w1100_,
		_w1095_,
		_w1101_
	);
	LUT3 #(
		.INIT('hac)
	) name860 (
		\shift_data_reg[0]/NET0131 ,
		\shift_data_reg[1]/NET0131 ,
		_w1015_,
		_w1102_
	);
	LUT2 #(
		.INIT('h8)
	) name861 (
		_w1014_,
		_w1102_,
		_w1103_
	);
	LUT3 #(
		.INIT('hac)
	) name862 (
		\shift_data_reg[2]/NET0131 ,
		\shift_data_reg[3]/NET0131 ,
		_w1015_,
		_w1104_
	);
	LUT2 #(
		.INIT('h4)
	) name863 (
		_w1014_,
		_w1104_,
		_w1105_
	);
	LUT3 #(
		.INIT('h01)
	) name864 (
		_w1024_,
		_w1105_,
		_w1103_,
		_w1106_
	);
	LUT3 #(
		.INIT('hac)
	) name865 (
		\shift_data_reg[6]/NET0131 ,
		\shift_data_reg[7]/NET0131 ,
		_w1015_,
		_w1107_
	);
	LUT2 #(
		.INIT('h4)
	) name866 (
		_w1014_,
		_w1107_,
		_w1108_
	);
	LUT3 #(
		.INIT('hac)
	) name867 (
		\shift_data_reg[4]/NET0131 ,
		\shift_data_reg[5]/NET0131 ,
		_w1015_,
		_w1109_
	);
	LUT2 #(
		.INIT('h8)
	) name868 (
		_w1014_,
		_w1109_,
		_w1110_
	);
	LUT3 #(
		.INIT('h02)
	) name869 (
		_w1024_,
		_w1110_,
		_w1108_,
		_w1111_
	);
	LUT3 #(
		.INIT('h02)
	) name870 (
		_w1032_,
		_w1111_,
		_w1106_,
		_w1112_
	);
	LUT3 #(
		.INIT('h54)
	) name871 (
		_w1042_,
		_w1101_,
		_w1112_,
		_w1113_
	);
	LUT3 #(
		.INIT('h02)
	) name872 (
		_w1053_,
		_w1113_,
		_w1090_,
		_w1114_
	);
	LUT3 #(
		.INIT('hac)
	) name873 (
		\shift_data_reg[56]/NET0131 ,
		\shift_data_reg[57]/NET0131 ,
		_w1015_,
		_w1115_
	);
	LUT2 #(
		.INIT('h8)
	) name874 (
		_w1014_,
		_w1115_,
		_w1116_
	);
	LUT3 #(
		.INIT('hac)
	) name875 (
		\shift_data_reg[58]/NET0131 ,
		\shift_data_reg[59]/NET0131 ,
		_w1015_,
		_w1117_
	);
	LUT2 #(
		.INIT('h4)
	) name876 (
		_w1014_,
		_w1117_,
		_w1118_
	);
	LUT3 #(
		.INIT('h01)
	) name877 (
		_w1024_,
		_w1118_,
		_w1116_,
		_w1119_
	);
	LUT3 #(
		.INIT('hac)
	) name878 (
		\shift_data_reg[62]/NET0131 ,
		\shift_data_reg[63]/NET0131 ,
		_w1015_,
		_w1120_
	);
	LUT2 #(
		.INIT('h4)
	) name879 (
		_w1014_,
		_w1120_,
		_w1121_
	);
	LUT3 #(
		.INIT('hac)
	) name880 (
		\shift_data_reg[60]/NET0131 ,
		\shift_data_reg[61]/NET0131 ,
		_w1015_,
		_w1122_
	);
	LUT2 #(
		.INIT('h8)
	) name881 (
		_w1014_,
		_w1122_,
		_w1123_
	);
	LUT3 #(
		.INIT('h02)
	) name882 (
		_w1024_,
		_w1123_,
		_w1121_,
		_w1124_
	);
	LUT3 #(
		.INIT('h01)
	) name883 (
		_w1032_,
		_w1124_,
		_w1119_,
		_w1125_
	);
	LUT3 #(
		.INIT('hac)
	) name884 (
		\shift_data_reg[52]/NET0131 ,
		\shift_data_reg[53]/NET0131 ,
		_w1015_,
		_w1126_
	);
	LUT2 #(
		.INIT('h8)
	) name885 (
		_w1014_,
		_w1126_,
		_w1127_
	);
	LUT3 #(
		.INIT('hac)
	) name886 (
		\shift_data_reg[54]/NET0131 ,
		\shift_data_reg[55]/NET0131 ,
		_w1015_,
		_w1128_
	);
	LUT2 #(
		.INIT('h4)
	) name887 (
		_w1014_,
		_w1128_,
		_w1129_
	);
	LUT3 #(
		.INIT('h02)
	) name888 (
		_w1024_,
		_w1129_,
		_w1127_,
		_w1130_
	);
	LUT3 #(
		.INIT('hac)
	) name889 (
		\shift_data_reg[50]/NET0131 ,
		\shift_data_reg[51]/NET0131 ,
		_w1015_,
		_w1131_
	);
	LUT2 #(
		.INIT('h4)
	) name890 (
		_w1014_,
		_w1131_,
		_w1132_
	);
	LUT3 #(
		.INIT('hac)
	) name891 (
		\shift_data_reg[48]/NET0131 ,
		\shift_data_reg[49]/NET0131 ,
		_w1015_,
		_w1133_
	);
	LUT2 #(
		.INIT('h8)
	) name892 (
		_w1014_,
		_w1133_,
		_w1134_
	);
	LUT3 #(
		.INIT('h01)
	) name893 (
		_w1024_,
		_w1134_,
		_w1132_,
		_w1135_
	);
	LUT3 #(
		.INIT('h02)
	) name894 (
		_w1032_,
		_w1135_,
		_w1130_,
		_w1136_
	);
	LUT3 #(
		.INIT('ha8)
	) name895 (
		_w1042_,
		_w1125_,
		_w1136_,
		_w1137_
	);
	LUT3 #(
		.INIT('hac)
	) name896 (
		\shift_data_reg[40]/NET0131 ,
		\shift_data_reg[41]/NET0131 ,
		_w1015_,
		_w1138_
	);
	LUT2 #(
		.INIT('h8)
	) name897 (
		_w1014_,
		_w1138_,
		_w1139_
	);
	LUT3 #(
		.INIT('hac)
	) name898 (
		\shift_data_reg[42]/NET0131 ,
		\shift_data_reg[43]/NET0131 ,
		_w1015_,
		_w1140_
	);
	LUT2 #(
		.INIT('h4)
	) name899 (
		_w1014_,
		_w1140_,
		_w1141_
	);
	LUT3 #(
		.INIT('h01)
	) name900 (
		_w1024_,
		_w1141_,
		_w1139_,
		_w1142_
	);
	LUT3 #(
		.INIT('hac)
	) name901 (
		\shift_data_reg[46]/NET0131 ,
		\shift_data_reg[47]/NET0131 ,
		_w1015_,
		_w1143_
	);
	LUT2 #(
		.INIT('h4)
	) name902 (
		_w1014_,
		_w1143_,
		_w1144_
	);
	LUT3 #(
		.INIT('hac)
	) name903 (
		\shift_data_reg[44]/NET0131 ,
		\shift_data_reg[45]/NET0131 ,
		_w1015_,
		_w1145_
	);
	LUT2 #(
		.INIT('h8)
	) name904 (
		_w1014_,
		_w1145_,
		_w1146_
	);
	LUT3 #(
		.INIT('h02)
	) name905 (
		_w1024_,
		_w1146_,
		_w1144_,
		_w1147_
	);
	LUT3 #(
		.INIT('h01)
	) name906 (
		_w1032_,
		_w1147_,
		_w1142_,
		_w1148_
	);
	LUT3 #(
		.INIT('hac)
	) name907 (
		\shift_data_reg[38]/NET0131 ,
		\shift_data_reg[39]/NET0131 ,
		_w1015_,
		_w1149_
	);
	LUT2 #(
		.INIT('h4)
	) name908 (
		_w1014_,
		_w1149_,
		_w1150_
	);
	LUT3 #(
		.INIT('hac)
	) name909 (
		\shift_data_reg[36]/NET0131 ,
		\shift_data_reg[37]/NET0131 ,
		_w1015_,
		_w1151_
	);
	LUT2 #(
		.INIT('h8)
	) name910 (
		_w1014_,
		_w1151_,
		_w1152_
	);
	LUT3 #(
		.INIT('h02)
	) name911 (
		_w1024_,
		_w1152_,
		_w1150_,
		_w1153_
	);
	LUT3 #(
		.INIT('hac)
	) name912 (
		\shift_data_reg[32]/NET0131 ,
		\shift_data_reg[33]/NET0131 ,
		_w1015_,
		_w1154_
	);
	LUT2 #(
		.INIT('h8)
	) name913 (
		_w1014_,
		_w1154_,
		_w1155_
	);
	LUT3 #(
		.INIT('hac)
	) name914 (
		\shift_data_reg[34]/NET0131 ,
		\shift_data_reg[35]/NET0131 ,
		_w1015_,
		_w1156_
	);
	LUT2 #(
		.INIT('h4)
	) name915 (
		_w1014_,
		_w1156_,
		_w1157_
	);
	LUT3 #(
		.INIT('h01)
	) name916 (
		_w1024_,
		_w1157_,
		_w1155_,
		_w1158_
	);
	LUT3 #(
		.INIT('h02)
	) name917 (
		_w1032_,
		_w1158_,
		_w1153_,
		_w1159_
	);
	LUT3 #(
		.INIT('h54)
	) name918 (
		_w1042_,
		_w1148_,
		_w1159_,
		_w1160_
	);
	LUT3 #(
		.INIT('hac)
	) name919 (
		\clgen_neg_edge_reg/NET0131 ,
		\clgen_pos_edge_reg/NET0131 ,
		\ctrl_reg[9]/NET0131 ,
		_w1161_
	);
	LUT4 #(
		.INIT('hef00)
	) name920 (
		sclk_pad_o_pad,
		\shift_cnt_reg[7]/NET0131 ,
		_w398_,
		_w1161_,
		_w1162_
	);
	LUT3 #(
		.INIT('h01)
	) name921 (
		_w1062_,
		_w1064_,
		_w1162_,
		_w1163_
	);
	LUT4 #(
		.INIT('hfe00)
	) name922 (
		_w1053_,
		_w1160_,
		_w1137_,
		_w1163_,
		_w1164_
	);
	LUT2 #(
		.INIT('h4)
	) name923 (
		_w1114_,
		_w1164_,
		_w1165_
	);
	LUT2 #(
		.INIT('h8)
	) name924 (
		miso_pad_i_pad,
		_w1162_,
		_w1166_
	);
	LUT3 #(
		.INIT('hac)
	) name925 (
		\shift_data_reg[80]/NET0131 ,
		\shift_data_reg[81]/NET0131 ,
		_w1015_,
		_w1167_
	);
	LUT2 #(
		.INIT('h8)
	) name926 (
		_w1014_,
		_w1167_,
		_w1168_
	);
	LUT3 #(
		.INIT('hac)
	) name927 (
		\shift_data_reg[82]/NET0131 ,
		\shift_data_reg[83]/NET0131 ,
		_w1015_,
		_w1169_
	);
	LUT2 #(
		.INIT('h4)
	) name928 (
		_w1014_,
		_w1169_,
		_w1170_
	);
	LUT3 #(
		.INIT('h01)
	) name929 (
		_w1024_,
		_w1170_,
		_w1168_,
		_w1171_
	);
	LUT3 #(
		.INIT('hac)
	) name930 (
		\shift_data_reg[86]/NET0131 ,
		\shift_data_reg[87]/NET0131 ,
		_w1015_,
		_w1172_
	);
	LUT2 #(
		.INIT('h4)
	) name931 (
		_w1014_,
		_w1172_,
		_w1173_
	);
	LUT3 #(
		.INIT('hac)
	) name932 (
		\shift_data_reg[84]/NET0131 ,
		\shift_data_reg[85]/NET0131 ,
		_w1015_,
		_w1174_
	);
	LUT2 #(
		.INIT('h8)
	) name933 (
		_w1014_,
		_w1174_,
		_w1175_
	);
	LUT3 #(
		.INIT('h02)
	) name934 (
		_w1024_,
		_w1175_,
		_w1173_,
		_w1176_
	);
	LUT3 #(
		.INIT('h02)
	) name935 (
		_w1032_,
		_w1176_,
		_w1171_,
		_w1177_
	);
	LUT3 #(
		.INIT('hac)
	) name936 (
		\shift_data_reg[88]/NET0131 ,
		\shift_data_reg[89]/NET0131 ,
		_w1015_,
		_w1178_
	);
	LUT2 #(
		.INIT('h8)
	) name937 (
		_w1014_,
		_w1178_,
		_w1179_
	);
	LUT3 #(
		.INIT('hac)
	) name938 (
		\shift_data_reg[90]/NET0131 ,
		\shift_data_reg[91]/NET0131 ,
		_w1015_,
		_w1180_
	);
	LUT2 #(
		.INIT('h4)
	) name939 (
		_w1014_,
		_w1180_,
		_w1181_
	);
	LUT3 #(
		.INIT('h01)
	) name940 (
		_w1024_,
		_w1181_,
		_w1179_,
		_w1182_
	);
	LUT3 #(
		.INIT('hac)
	) name941 (
		\shift_data_reg[94]/NET0131 ,
		\shift_data_reg[95]/NET0131 ,
		_w1015_,
		_w1183_
	);
	LUT2 #(
		.INIT('h4)
	) name942 (
		_w1014_,
		_w1183_,
		_w1184_
	);
	LUT3 #(
		.INIT('hac)
	) name943 (
		\shift_data_reg[92]/NET0131 ,
		\shift_data_reg[93]/NET0131 ,
		_w1015_,
		_w1185_
	);
	LUT2 #(
		.INIT('h8)
	) name944 (
		_w1014_,
		_w1185_,
		_w1186_
	);
	LUT3 #(
		.INIT('h02)
	) name945 (
		_w1024_,
		_w1186_,
		_w1184_,
		_w1187_
	);
	LUT3 #(
		.INIT('h01)
	) name946 (
		_w1032_,
		_w1187_,
		_w1182_,
		_w1188_
	);
	LUT3 #(
		.INIT('ha8)
	) name947 (
		_w1042_,
		_w1177_,
		_w1188_,
		_w1189_
	);
	LUT3 #(
		.INIT('hac)
	) name948 (
		\shift_data_reg[72]/NET0131 ,
		\shift_data_reg[73]/NET0131 ,
		_w1015_,
		_w1190_
	);
	LUT2 #(
		.INIT('h8)
	) name949 (
		_w1014_,
		_w1190_,
		_w1191_
	);
	LUT3 #(
		.INIT('hac)
	) name950 (
		\shift_data_reg[74]/NET0131 ,
		\shift_data_reg[75]/NET0131 ,
		_w1015_,
		_w1192_
	);
	LUT2 #(
		.INIT('h4)
	) name951 (
		_w1014_,
		_w1192_,
		_w1193_
	);
	LUT3 #(
		.INIT('h01)
	) name952 (
		_w1024_,
		_w1193_,
		_w1191_,
		_w1194_
	);
	LUT3 #(
		.INIT('hac)
	) name953 (
		\shift_data_reg[78]/NET0131 ,
		\shift_data_reg[79]/NET0131 ,
		_w1015_,
		_w1195_
	);
	LUT2 #(
		.INIT('h4)
	) name954 (
		_w1014_,
		_w1195_,
		_w1196_
	);
	LUT3 #(
		.INIT('hac)
	) name955 (
		\shift_data_reg[76]/NET0131 ,
		\shift_data_reg[77]/NET0131 ,
		_w1015_,
		_w1197_
	);
	LUT2 #(
		.INIT('h8)
	) name956 (
		_w1014_,
		_w1197_,
		_w1198_
	);
	LUT3 #(
		.INIT('h02)
	) name957 (
		_w1024_,
		_w1198_,
		_w1196_,
		_w1199_
	);
	LUT3 #(
		.INIT('h01)
	) name958 (
		_w1032_,
		_w1199_,
		_w1194_,
		_w1200_
	);
	LUT3 #(
		.INIT('hac)
	) name959 (
		\shift_data_reg[64]/NET0131 ,
		\shift_data_reg[65]/NET0131 ,
		_w1015_,
		_w1201_
	);
	LUT2 #(
		.INIT('h8)
	) name960 (
		_w1014_,
		_w1201_,
		_w1202_
	);
	LUT3 #(
		.INIT('hac)
	) name961 (
		\shift_data_reg[66]/NET0131 ,
		\shift_data_reg[67]/NET0131 ,
		_w1015_,
		_w1203_
	);
	LUT2 #(
		.INIT('h4)
	) name962 (
		_w1014_,
		_w1203_,
		_w1204_
	);
	LUT3 #(
		.INIT('h01)
	) name963 (
		_w1024_,
		_w1204_,
		_w1202_,
		_w1205_
	);
	LUT3 #(
		.INIT('hac)
	) name964 (
		\shift_data_reg[70]/NET0131 ,
		\shift_data_reg[71]/NET0131 ,
		_w1015_,
		_w1206_
	);
	LUT2 #(
		.INIT('h4)
	) name965 (
		_w1014_,
		_w1206_,
		_w1207_
	);
	LUT3 #(
		.INIT('hac)
	) name966 (
		\shift_data_reg[68]/NET0131 ,
		\shift_data_reg[69]/NET0131 ,
		_w1015_,
		_w1208_
	);
	LUT2 #(
		.INIT('h8)
	) name967 (
		_w1014_,
		_w1208_,
		_w1209_
	);
	LUT3 #(
		.INIT('h02)
	) name968 (
		_w1024_,
		_w1209_,
		_w1207_,
		_w1210_
	);
	LUT3 #(
		.INIT('h02)
	) name969 (
		_w1032_,
		_w1210_,
		_w1205_,
		_w1211_
	);
	LUT3 #(
		.INIT('h54)
	) name970 (
		_w1042_,
		_w1200_,
		_w1211_,
		_w1212_
	);
	LUT3 #(
		.INIT('h02)
	) name971 (
		_w1053_,
		_w1212_,
		_w1189_,
		_w1213_
	);
	LUT3 #(
		.INIT('hac)
	) name972 (
		\shift_data_reg[116]/NET0131 ,
		\shift_data_reg[117]/NET0131 ,
		_w1015_,
		_w1214_
	);
	LUT2 #(
		.INIT('h8)
	) name973 (
		_w1014_,
		_w1214_,
		_w1215_
	);
	LUT3 #(
		.INIT('hac)
	) name974 (
		\shift_data_reg[118]/NET0131 ,
		\shift_data_reg[119]/NET0131 ,
		_w1015_,
		_w1216_
	);
	LUT2 #(
		.INIT('h4)
	) name975 (
		_w1014_,
		_w1216_,
		_w1217_
	);
	LUT3 #(
		.INIT('h02)
	) name976 (
		_w1024_,
		_w1217_,
		_w1215_,
		_w1218_
	);
	LUT3 #(
		.INIT('hac)
	) name977 (
		\shift_data_reg[114]/NET0131 ,
		\shift_data_reg[115]/NET0131 ,
		_w1015_,
		_w1219_
	);
	LUT2 #(
		.INIT('h4)
	) name978 (
		_w1014_,
		_w1219_,
		_w1220_
	);
	LUT3 #(
		.INIT('hac)
	) name979 (
		\shift_data_reg[112]/NET0131 ,
		\shift_data_reg[113]/NET0131 ,
		_w1015_,
		_w1221_
	);
	LUT2 #(
		.INIT('h8)
	) name980 (
		_w1014_,
		_w1221_,
		_w1222_
	);
	LUT3 #(
		.INIT('h01)
	) name981 (
		_w1024_,
		_w1222_,
		_w1220_,
		_w1223_
	);
	LUT3 #(
		.INIT('h02)
	) name982 (
		_w1032_,
		_w1223_,
		_w1218_,
		_w1224_
	);
	LUT3 #(
		.INIT('hac)
	) name983 (
		\shift_data_reg[124]/NET0131 ,
		\shift_data_reg[125]/NET0131 ,
		_w1015_,
		_w1225_
	);
	LUT2 #(
		.INIT('h8)
	) name984 (
		_w1014_,
		_w1225_,
		_w1226_
	);
	LUT3 #(
		.INIT('hac)
	) name985 (
		\shift_data_reg[126]/NET0131 ,
		\shift_data_reg[127]/NET0131 ,
		_w1015_,
		_w1227_
	);
	LUT2 #(
		.INIT('h4)
	) name986 (
		_w1014_,
		_w1227_,
		_w1228_
	);
	LUT3 #(
		.INIT('h02)
	) name987 (
		_w1024_,
		_w1228_,
		_w1226_,
		_w1229_
	);
	LUT3 #(
		.INIT('hac)
	) name988 (
		\shift_data_reg[122]/NET0131 ,
		\shift_data_reg[123]/NET0131 ,
		_w1015_,
		_w1230_
	);
	LUT2 #(
		.INIT('h4)
	) name989 (
		_w1014_,
		_w1230_,
		_w1231_
	);
	LUT3 #(
		.INIT('hac)
	) name990 (
		\shift_data_reg[120]/NET0131 ,
		\shift_data_reg[121]/NET0131 ,
		_w1015_,
		_w1232_
	);
	LUT2 #(
		.INIT('h8)
	) name991 (
		_w1014_,
		_w1232_,
		_w1233_
	);
	LUT3 #(
		.INIT('h01)
	) name992 (
		_w1024_,
		_w1233_,
		_w1231_,
		_w1234_
	);
	LUT3 #(
		.INIT('h01)
	) name993 (
		_w1032_,
		_w1234_,
		_w1229_,
		_w1235_
	);
	LUT3 #(
		.INIT('h02)
	) name994 (
		_w1042_,
		_w1235_,
		_w1224_,
		_w1236_
	);
	LUT3 #(
		.INIT('hac)
	) name995 (
		\shift_data_reg[108]/NET0131 ,
		\shift_data_reg[109]/NET0131 ,
		_w1015_,
		_w1237_
	);
	LUT2 #(
		.INIT('h8)
	) name996 (
		_w1014_,
		_w1237_,
		_w1238_
	);
	LUT3 #(
		.INIT('hac)
	) name997 (
		\shift_data_reg[110]/NET0131 ,
		\shift_data_reg[111]/NET0131 ,
		_w1015_,
		_w1239_
	);
	LUT2 #(
		.INIT('h4)
	) name998 (
		_w1014_,
		_w1239_,
		_w1240_
	);
	LUT3 #(
		.INIT('h02)
	) name999 (
		_w1024_,
		_w1240_,
		_w1238_,
		_w1241_
	);
	LUT3 #(
		.INIT('hac)
	) name1000 (
		\shift_data_reg[106]/NET0131 ,
		\shift_data_reg[107]/NET0131 ,
		_w1015_,
		_w1242_
	);
	LUT2 #(
		.INIT('h4)
	) name1001 (
		_w1014_,
		_w1242_,
		_w1243_
	);
	LUT3 #(
		.INIT('hac)
	) name1002 (
		\shift_data_reg[104]/NET0131 ,
		\shift_data_reg[105]/NET0131 ,
		_w1015_,
		_w1244_
	);
	LUT2 #(
		.INIT('h8)
	) name1003 (
		_w1014_,
		_w1244_,
		_w1245_
	);
	LUT3 #(
		.INIT('h01)
	) name1004 (
		_w1024_,
		_w1245_,
		_w1243_,
		_w1246_
	);
	LUT3 #(
		.INIT('h01)
	) name1005 (
		_w1032_,
		_w1246_,
		_w1241_,
		_w1247_
	);
	LUT3 #(
		.INIT('hac)
	) name1006 (
		\shift_data_reg[100]/NET0131 ,
		\shift_data_reg[101]/NET0131 ,
		_w1015_,
		_w1248_
	);
	LUT2 #(
		.INIT('h8)
	) name1007 (
		_w1014_,
		_w1248_,
		_w1249_
	);
	LUT3 #(
		.INIT('hac)
	) name1008 (
		\shift_data_reg[102]/NET0131 ,
		\shift_data_reg[103]/NET0131 ,
		_w1015_,
		_w1250_
	);
	LUT2 #(
		.INIT('h4)
	) name1009 (
		_w1014_,
		_w1250_,
		_w1251_
	);
	LUT3 #(
		.INIT('h02)
	) name1010 (
		_w1024_,
		_w1251_,
		_w1249_,
		_w1252_
	);
	LUT3 #(
		.INIT('hac)
	) name1011 (
		\shift_data_reg[98]/NET0131 ,
		\shift_data_reg[99]/NET0131 ,
		_w1015_,
		_w1253_
	);
	LUT2 #(
		.INIT('h4)
	) name1012 (
		_w1014_,
		_w1253_,
		_w1254_
	);
	LUT3 #(
		.INIT('hac)
	) name1013 (
		\shift_data_reg[96]/NET0131 ,
		\shift_data_reg[97]/NET0131 ,
		_w1015_,
		_w1255_
	);
	LUT2 #(
		.INIT('h8)
	) name1014 (
		_w1014_,
		_w1255_,
		_w1256_
	);
	LUT3 #(
		.INIT('h01)
	) name1015 (
		_w1024_,
		_w1256_,
		_w1254_,
		_w1257_
	);
	LUT3 #(
		.INIT('h02)
	) name1016 (
		_w1032_,
		_w1257_,
		_w1252_,
		_w1258_
	);
	LUT3 #(
		.INIT('h01)
	) name1017 (
		_w1042_,
		_w1258_,
		_w1247_,
		_w1259_
	);
	LUT3 #(
		.INIT('h0e)
	) name1018 (
		_w1062_,
		_w1064_,
		_w1162_,
		_w1260_
	);
	LUT4 #(
		.INIT('hab00)
	) name1019 (
		_w1053_,
		_w1236_,
		_w1259_,
		_w1260_,
		_w1261_
	);
	LUT3 #(
		.INIT('h45)
	) name1020 (
		_w1166_,
		_w1213_,
		_w1261_,
		_w1262_
	);
	LUT4 #(
		.INIT('h4000)
	) name1021 (
		\wb_adr_i[3]_pad ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		wb_we_i_pad,
		_w1263_
	);
	LUT2 #(
		.INIT('h8)
	) name1022 (
		_w1055_,
		_w1263_,
		_w1264_
	);
	LUT4 #(
		.INIT('h1555)
	) name1023 (
		\shift_data_reg[55]/NET0131 ,
		_w1033_,
		_w1054_,
		_w1066_,
		_w1265_
	);
	LUT2 #(
		.INIT('h1)
	) name1024 (
		_w1264_,
		_w1265_,
		_w1266_
	);
	LUT4 #(
		.INIT('hdf00)
	) name1025 (
		_w1067_,
		_w1165_,
		_w1262_,
		_w1266_,
		_w1267_
	);
	LUT3 #(
		.INIT('h80)
	) name1026 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1268_
	);
	LUT2 #(
		.INIT('h8)
	) name1027 (
		\wb_dat_i[23]_pad ,
		\wb_sel_i[2]_pad ,
		_w1269_
	);
	LUT4 #(
		.INIT('h8000)
	) name1028 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1269_,
		_w1270_
	);
	LUT2 #(
		.INIT('h8)
	) name1029 (
		\wb_adr_i[2]_pad ,
		\wb_sel_i[2]_pad ,
		_w1271_
	);
	LUT4 #(
		.INIT('h0080)
	) name1030 (
		\shift_data_reg[55]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1271_,
		_w1272_
	);
	LUT2 #(
		.INIT('h1)
	) name1031 (
		_w1270_,
		_w1272_,
		_w1273_
	);
	LUT2 #(
		.INIT('hb)
	) name1032 (
		_w1267_,
		_w1273_,
		_w1274_
	);
	LUT3 #(
		.INIT('h80)
	) name1033 (
		_w804_,
		_w826_,
		_w1057_,
		_w1275_
	);
	LUT2 #(
		.INIT('h2)
	) name1034 (
		_w1014_,
		_w1015_,
		_w1276_
	);
	LUT2 #(
		.INIT('h8)
	) name1035 (
		_w1024_,
		_w1276_,
		_w1277_
	);
	LUT3 #(
		.INIT('h54)
	) name1036 (
		_w1042_,
		_w1049_,
		_w1052_,
		_w1278_
	);
	LUT3 #(
		.INIT('ha8)
	) name1037 (
		_w1032_,
		_w1062_,
		_w1064_,
		_w1279_
	);
	LUT3 #(
		.INIT('h80)
	) name1038 (
		_w1277_,
		_w1278_,
		_w1279_,
		_w1280_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1039 (
		_w1060_,
		_w1165_,
		_w1262_,
		_w1280_,
		_w1281_
	);
	LUT4 #(
		.INIT('h1555)
	) name1040 (
		_w1059_,
		_w1277_,
		_w1278_,
		_w1279_,
		_w1282_
	);
	LUT4 #(
		.INIT('h373f)
	) name1041 (
		_w585_,
		_w1055_,
		_w1263_,
		_w1056_,
		_w1283_
	);
	LUT3 #(
		.INIT('h40)
	) name1042 (
		\wb_sel_i[0]_pad ,
		_w804_,
		_w1057_,
		_w1284_
	);
	LUT2 #(
		.INIT('h2)
	) name1043 (
		_w1283_,
		_w1284_,
		_w1285_
	);
	LUT3 #(
		.INIT('h8a)
	) name1044 (
		\shift_data_reg[101]/NET0131 ,
		_w1282_,
		_w1285_,
		_w1286_
	);
	LUT4 #(
		.INIT('hff54)
	) name1045 (
		_w1264_,
		_w1275_,
		_w1281_,
		_w1286_,
		_w1287_
	);
	LUT4 #(
		.INIT('h1000)
	) name1046 (
		_w1032_,
		_w1065_,
		_w1277_,
		_w1278_,
		_w1288_
	);
	LUT2 #(
		.INIT('h4)
	) name1047 (
		_w1264_,
		_w1060_,
		_w1289_
	);
	LUT3 #(
		.INIT('hc8)
	) name1048 (
		\shift_data_reg[109]/NET0131 ,
		_w1289_,
		_w1288_,
		_w1290_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1049 (
		_w1165_,
		_w1262_,
		_w1288_,
		_w1290_,
		_w1291_
	);
	LUT2 #(
		.INIT('h2)
	) name1050 (
		\shift_data_reg[109]/NET0131 ,
		\wb_sel_i[1]_pad ,
		_w1292_
	);
	LUT4 #(
		.INIT('h00d5)
	) name1051 (
		_w822_,
		_w1055_,
		_w1263_,
		_w1292_,
		_w1293_
	);
	LUT4 #(
		.INIT('hf531)
	) name1052 (
		\shift_data_reg[109]/NET0131 ,
		_w1059_,
		_w1283_,
		_w1293_,
		_w1294_
	);
	LUT2 #(
		.INIT('hb)
	) name1053 (
		_w1291_,
		_w1294_,
		_w1295_
	);
	LUT2 #(
		.INIT('h4)
	) name1054 (
		_w1014_,
		_w1015_,
		_w1296_
	);
	LUT2 #(
		.INIT('h8)
	) name1055 (
		_w1024_,
		_w1296_,
		_w1297_
	);
	LUT4 #(
		.INIT('h1000)
	) name1056 (
		_w1032_,
		_w1065_,
		_w1278_,
		_w1297_,
		_w1298_
	);
	LUT3 #(
		.INIT('hc8)
	) name1057 (
		\shift_data_reg[110]/NET0131 ,
		_w1289_,
		_w1298_,
		_w1299_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1058 (
		_w1165_,
		_w1262_,
		_w1298_,
		_w1299_,
		_w1300_
	);
	LUT2 #(
		.INIT('h2)
	) name1059 (
		\shift_data_reg[110]/NET0131 ,
		\wb_sel_i[1]_pad ,
		_w1301_
	);
	LUT4 #(
		.INIT('h00d5)
	) name1060 (
		_w844_,
		_w1055_,
		_w1263_,
		_w1301_,
		_w1302_
	);
	LUT4 #(
		.INIT('hf531)
	) name1061 (
		\shift_data_reg[110]/NET0131 ,
		_w1059_,
		_w1283_,
		_w1302_,
		_w1303_
	);
	LUT2 #(
		.INIT('hb)
	) name1062 (
		_w1300_,
		_w1303_,
		_w1304_
	);
	LUT2 #(
		.INIT('h8)
	) name1063 (
		_w1014_,
		_w1015_,
		_w1305_
	);
	LUT2 #(
		.INIT('h4)
	) name1064 (
		_w1024_,
		_w1305_,
		_w1306_
	);
	LUT4 #(
		.INIT('h0008)
	) name1065 (
		_w1032_,
		_w1060_,
		_w1062_,
		_w1064_,
		_w1307_
	);
	LUT3 #(
		.INIT('h80)
	) name1066 (
		_w1278_,
		_w1306_,
		_w1307_,
		_w1308_
	);
	LUT4 #(
		.INIT('h1555)
	) name1067 (
		\shift_data_reg[32]/NET0131 ,
		_w1278_,
		_w1306_,
		_w1307_,
		_w1309_
	);
	LUT2 #(
		.INIT('h1)
	) name1068 (
		_w1264_,
		_w1309_,
		_w1310_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1069 (
		_w1165_,
		_w1262_,
		_w1308_,
		_w1310_,
		_w1311_
	);
	LUT4 #(
		.INIT('h8000)
	) name1070 (
		\wb_adr_i[2]_pad ,
		_w889_,
		_w1055_,
		_w1263_,
		_w1312_
	);
	LUT2 #(
		.INIT('h8)
	) name1071 (
		\wb_adr_i[2]_pad ,
		\wb_sel_i[0]_pad ,
		_w1313_
	);
	LUT4 #(
		.INIT('h0080)
	) name1072 (
		\shift_data_reg[32]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1313_,
		_w1314_
	);
	LUT2 #(
		.INIT('h1)
	) name1073 (
		_w1312_,
		_w1314_,
		_w1315_
	);
	LUT2 #(
		.INIT('hb)
	) name1074 (
		_w1311_,
		_w1315_,
		_w1316_
	);
	LUT3 #(
		.INIT('h80)
	) name1075 (
		_w1025_,
		_w1278_,
		_w1307_,
		_w1317_
	);
	LUT4 #(
		.INIT('h1555)
	) name1076 (
		\shift_data_reg[39]/NET0131 ,
		_w1025_,
		_w1278_,
		_w1307_,
		_w1318_
	);
	LUT2 #(
		.INIT('h1)
	) name1077 (
		_w1264_,
		_w1318_,
		_w1319_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1078 (
		_w1165_,
		_w1262_,
		_w1317_,
		_w1319_,
		_w1320_
	);
	LUT4 #(
		.INIT('h8000)
	) name1079 (
		\wb_adr_i[2]_pad ,
		_w818_,
		_w1055_,
		_w1263_,
		_w1321_
	);
	LUT4 #(
		.INIT('h0080)
	) name1080 (
		\shift_data_reg[39]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1313_,
		_w1322_
	);
	LUT2 #(
		.INIT('h1)
	) name1081 (
		_w1321_,
		_w1322_,
		_w1323_
	);
	LUT2 #(
		.INIT('hb)
	) name1082 (
		_w1320_,
		_w1323_,
		_w1324_
	);
	LUT4 #(
		.INIT('h0004)
	) name1083 (
		_w1032_,
		_w1060_,
		_w1062_,
		_w1064_,
		_w1325_
	);
	LUT3 #(
		.INIT('h80)
	) name1084 (
		_w1025_,
		_w1054_,
		_w1325_,
		_w1326_
	);
	LUT4 #(
		.INIT('h1555)
	) name1085 (
		\shift_data_reg[63]/NET0131 ,
		_w1025_,
		_w1054_,
		_w1325_,
		_w1327_
	);
	LUT2 #(
		.INIT('h1)
	) name1086 (
		_w1264_,
		_w1327_,
		_w1328_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1087 (
		_w1165_,
		_w1262_,
		_w1326_,
		_w1328_,
		_w1329_
	);
	LUT2 #(
		.INIT('h8)
	) name1088 (
		\wb_dat_i[31]_pad ,
		\wb_sel_i[3]_pad ,
		_w1330_
	);
	LUT4 #(
		.INIT('h8000)
	) name1089 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1330_,
		_w1331_
	);
	LUT2 #(
		.INIT('h8)
	) name1090 (
		\wb_adr_i[2]_pad ,
		\wb_sel_i[3]_pad ,
		_w1332_
	);
	LUT4 #(
		.INIT('h0080)
	) name1091 (
		\shift_data_reg[63]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1332_,
		_w1333_
	);
	LUT2 #(
		.INIT('h1)
	) name1092 (
		_w1331_,
		_w1333_,
		_w1334_
	);
	LUT2 #(
		.INIT('hb)
	) name1093 (
		_w1329_,
		_w1334_,
		_w1335_
	);
	LUT3 #(
		.INIT('h80)
	) name1094 (
		_w1054_,
		_w1306_,
		_w1325_,
		_w1336_
	);
	LUT4 #(
		.INIT('h1555)
	) name1095 (
		\shift_data_reg[56]/NET0131 ,
		_w1054_,
		_w1306_,
		_w1325_,
		_w1337_
	);
	LUT2 #(
		.INIT('h1)
	) name1096 (
		_w1264_,
		_w1337_,
		_w1338_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1097 (
		_w1165_,
		_w1262_,
		_w1336_,
		_w1338_,
		_w1339_
	);
	LUT2 #(
		.INIT('h8)
	) name1098 (
		\wb_dat_i[24]_pad ,
		\wb_sel_i[3]_pad ,
		_w1340_
	);
	LUT4 #(
		.INIT('h8000)
	) name1099 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1340_,
		_w1341_
	);
	LUT4 #(
		.INIT('h0080)
	) name1100 (
		\shift_data_reg[56]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1332_,
		_w1342_
	);
	LUT2 #(
		.INIT('h1)
	) name1101 (
		_w1341_,
		_w1342_,
		_w1343_
	);
	LUT2 #(
		.INIT('hb)
	) name1102 (
		_w1339_,
		_w1343_,
		_w1344_
	);
	LUT3 #(
		.INIT('h80)
	) name1103 (
		\shift_data_reg[89]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1345_
	);
	LUT3 #(
		.INIT('h40)
	) name1104 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1346_
	);
	LUT2 #(
		.INIT('h8)
	) name1105 (
		\wb_dat_i[25]_pad ,
		\wb_sel_i[3]_pad ,
		_w1347_
	);
	LUT3 #(
		.INIT('h35)
	) name1106 (
		\shift_data_reg[89]/NET0131 ,
		\wb_dat_i[25]_pad ,
		\wb_sel_i[3]_pad ,
		_w1348_
	);
	LUT3 #(
		.INIT('h08)
	) name1107 (
		_w585_,
		_w1057_,
		_w1348_,
		_w1349_
	);
	LUT3 #(
		.INIT('h54)
	) name1108 (
		_w1059_,
		_w1062_,
		_w1064_,
		_w1350_
	);
	LUT3 #(
		.INIT('h02)
	) name1109 (
		_w1042_,
		_w1049_,
		_w1052_,
		_w1351_
	);
	LUT2 #(
		.INIT('h4)
	) name1110 (
		_w1024_,
		_w1276_,
		_w1352_
	);
	LUT4 #(
		.INIT('h4000)
	) name1111 (
		_w1032_,
		_w1350_,
		_w1351_,
		_w1352_,
		_w1353_
	);
	LUT2 #(
		.INIT('h1)
	) name1112 (
		_w1268_,
		_w1058_,
		_w1354_
	);
	LUT3 #(
		.INIT('he0)
	) name1113 (
		\shift_data_reg[89]/NET0131 ,
		_w1353_,
		_w1354_,
		_w1355_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1114 (
		_w1165_,
		_w1262_,
		_w1353_,
		_w1355_,
		_w1356_
	);
	LUT4 #(
		.INIT('hbbba)
	) name1115 (
		_w1345_,
		_w1346_,
		_w1349_,
		_w1356_,
		_w1357_
	);
	LUT2 #(
		.INIT('h8)
	) name1116 (
		\wb_dat_i[28]_pad ,
		\wb_sel_i[3]_pad ,
		_w1358_
	);
	LUT3 #(
		.INIT('h35)
	) name1117 (
		\shift_data_reg[92]/NET0131 ,
		\wb_dat_i[28]_pad ,
		\wb_sel_i[3]_pad ,
		_w1359_
	);
	LUT3 #(
		.INIT('h08)
	) name1118 (
		_w585_,
		_w1057_,
		_w1359_,
		_w1360_
	);
	LUT2 #(
		.INIT('h8)
	) name1119 (
		_w1024_,
		_w1305_,
		_w1361_
	);
	LUT4 #(
		.INIT('h4000)
	) name1120 (
		_w1032_,
		_w1350_,
		_w1351_,
		_w1361_,
		_w1362_
	);
	LUT3 #(
		.INIT('hc8)
	) name1121 (
		\shift_data_reg[92]/NET0131 ,
		_w1354_,
		_w1362_,
		_w1363_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1122 (
		_w1165_,
		_w1262_,
		_w1362_,
		_w1363_,
		_w1364_
	);
	LUT3 #(
		.INIT('h80)
	) name1123 (
		\shift_data_reg[92]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1365_
	);
	LUT4 #(
		.INIT('hff54)
	) name1124 (
		_w1346_,
		_w1360_,
		_w1364_,
		_w1365_,
		_w1366_
	);
	LUT3 #(
		.INIT('h35)
	) name1125 (
		\shift_data_reg[64]/NET0131 ,
		\wb_dat_i[0]_pad ,
		\wb_sel_i[0]_pad ,
		_w1367_
	);
	LUT3 #(
		.INIT('h08)
	) name1126 (
		_w585_,
		_w1057_,
		_w1367_,
		_w1368_
	);
	LUT2 #(
		.INIT('h8)
	) name1127 (
		_w1032_,
		_w1306_,
		_w1369_
	);
	LUT3 #(
		.INIT('h01)
	) name1128 (
		_w1042_,
		_w1049_,
		_w1052_,
		_w1370_
	);
	LUT3 #(
		.INIT('h80)
	) name1129 (
		_w1350_,
		_w1369_,
		_w1370_,
		_w1371_
	);
	LUT4 #(
		.INIT('h1555)
	) name1130 (
		\shift_data_reg[64]/NET0131 ,
		_w1350_,
		_w1369_,
		_w1370_,
		_w1372_
	);
	LUT2 #(
		.INIT('h2)
	) name1131 (
		_w1354_,
		_w1372_,
		_w1373_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1132 (
		_w1165_,
		_w1262_,
		_w1371_,
		_w1373_,
		_w1374_
	);
	LUT3 #(
		.INIT('h80)
	) name1133 (
		\shift_data_reg[64]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1375_
	);
	LUT4 #(
		.INIT('hff54)
	) name1134 (
		_w1346_,
		_w1368_,
		_w1374_,
		_w1375_,
		_w1376_
	);
	LUT3 #(
		.INIT('h35)
	) name1135 (
		\shift_data_reg[65]/NET0131 ,
		\wb_dat_i[1]_pad ,
		\wb_sel_i[0]_pad ,
		_w1377_
	);
	LUT3 #(
		.INIT('h08)
	) name1136 (
		_w585_,
		_w1057_,
		_w1377_,
		_w1378_
	);
	LUT2 #(
		.INIT('h8)
	) name1137 (
		_w1032_,
		_w1352_,
		_w1379_
	);
	LUT3 #(
		.INIT('h80)
	) name1138 (
		_w1350_,
		_w1370_,
		_w1379_,
		_w1380_
	);
	LUT4 #(
		.INIT('h1555)
	) name1139 (
		\shift_data_reg[65]/NET0131 ,
		_w1350_,
		_w1370_,
		_w1379_,
		_w1381_
	);
	LUT2 #(
		.INIT('h2)
	) name1140 (
		_w1354_,
		_w1381_,
		_w1382_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1141 (
		_w1165_,
		_w1262_,
		_w1380_,
		_w1382_,
		_w1383_
	);
	LUT3 #(
		.INIT('h80)
	) name1142 (
		\shift_data_reg[65]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1384_
	);
	LUT4 #(
		.INIT('hff54)
	) name1143 (
		_w1346_,
		_w1378_,
		_w1383_,
		_w1384_,
		_w1385_
	);
	LUT3 #(
		.INIT('h35)
	) name1144 (
		\shift_data_reg[66]/NET0131 ,
		\wb_dat_i[2]_pad ,
		\wb_sel_i[0]_pad ,
		_w1386_
	);
	LUT3 #(
		.INIT('h08)
	) name1145 (
		_w585_,
		_w1057_,
		_w1386_,
		_w1387_
	);
	LUT2 #(
		.INIT('h4)
	) name1146 (
		_w1024_,
		_w1296_,
		_w1388_
	);
	LUT2 #(
		.INIT('h8)
	) name1147 (
		_w1032_,
		_w1388_,
		_w1389_
	);
	LUT3 #(
		.INIT('h80)
	) name1148 (
		_w1350_,
		_w1370_,
		_w1389_,
		_w1390_
	);
	LUT4 #(
		.INIT('h1555)
	) name1149 (
		\shift_data_reg[66]/NET0131 ,
		_w1350_,
		_w1370_,
		_w1389_,
		_w1391_
	);
	LUT2 #(
		.INIT('h2)
	) name1150 (
		_w1354_,
		_w1391_,
		_w1392_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1151 (
		_w1165_,
		_w1262_,
		_w1390_,
		_w1392_,
		_w1393_
	);
	LUT3 #(
		.INIT('h80)
	) name1152 (
		\shift_data_reg[66]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1394_
	);
	LUT4 #(
		.INIT('hff54)
	) name1153 (
		_w1346_,
		_w1387_,
		_w1393_,
		_w1394_,
		_w1395_
	);
	LUT3 #(
		.INIT('h35)
	) name1154 (
		\shift_data_reg[67]/NET0131 ,
		\wb_dat_i[3]_pad ,
		\wb_sel_i[0]_pad ,
		_w1396_
	);
	LUT3 #(
		.INIT('h08)
	) name1155 (
		_w585_,
		_w1057_,
		_w1396_,
		_w1397_
	);
	LUT2 #(
		.INIT('h2)
	) name1156 (
		_w1016_,
		_w1024_,
		_w1398_
	);
	LUT4 #(
		.INIT('h8000)
	) name1157 (
		_w1032_,
		_w1350_,
		_w1370_,
		_w1398_,
		_w1399_
	);
	LUT3 #(
		.INIT('hc8)
	) name1158 (
		\shift_data_reg[67]/NET0131 ,
		_w1354_,
		_w1399_,
		_w1400_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1159 (
		_w1165_,
		_w1262_,
		_w1399_,
		_w1400_,
		_w1401_
	);
	LUT3 #(
		.INIT('h80)
	) name1160 (
		\shift_data_reg[67]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1402_
	);
	LUT4 #(
		.INIT('hff54)
	) name1161 (
		_w1346_,
		_w1397_,
		_w1401_,
		_w1402_,
		_w1403_
	);
	LUT3 #(
		.INIT('h35)
	) name1162 (
		\shift_data_reg[68]/NET0131 ,
		\wb_dat_i[4]_pad ,
		\wb_sel_i[0]_pad ,
		_w1404_
	);
	LUT3 #(
		.INIT('h08)
	) name1163 (
		_w585_,
		_w1057_,
		_w1404_,
		_w1405_
	);
	LUT2 #(
		.INIT('h8)
	) name1164 (
		_w1032_,
		_w1361_,
		_w1406_
	);
	LUT3 #(
		.INIT('h80)
	) name1165 (
		_w1350_,
		_w1370_,
		_w1406_,
		_w1407_
	);
	LUT4 #(
		.INIT('h1555)
	) name1166 (
		\shift_data_reg[68]/NET0131 ,
		_w1350_,
		_w1370_,
		_w1406_,
		_w1408_
	);
	LUT2 #(
		.INIT('h2)
	) name1167 (
		_w1354_,
		_w1408_,
		_w1409_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1168 (
		_w1165_,
		_w1262_,
		_w1407_,
		_w1409_,
		_w1410_
	);
	LUT3 #(
		.INIT('h80)
	) name1169 (
		\shift_data_reg[68]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1411_
	);
	LUT4 #(
		.INIT('hff54)
	) name1170 (
		_w1346_,
		_w1405_,
		_w1410_,
		_w1411_,
		_w1412_
	);
	LUT3 #(
		.INIT('h35)
	) name1171 (
		\shift_data_reg[69]/NET0131 ,
		\wb_dat_i[5]_pad ,
		\wb_sel_i[0]_pad ,
		_w1413_
	);
	LUT3 #(
		.INIT('h08)
	) name1172 (
		_w585_,
		_w1057_,
		_w1413_,
		_w1414_
	);
	LUT4 #(
		.INIT('h8000)
	) name1173 (
		_w1032_,
		_w1277_,
		_w1350_,
		_w1370_,
		_w1415_
	);
	LUT3 #(
		.INIT('hc8)
	) name1174 (
		\shift_data_reg[69]/NET0131 ,
		_w1354_,
		_w1415_,
		_w1416_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1175 (
		_w1165_,
		_w1262_,
		_w1415_,
		_w1416_,
		_w1417_
	);
	LUT3 #(
		.INIT('h80)
	) name1176 (
		\shift_data_reg[69]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1418_
	);
	LUT4 #(
		.INIT('hff54)
	) name1177 (
		_w1346_,
		_w1414_,
		_w1417_,
		_w1418_,
		_w1419_
	);
	LUT3 #(
		.INIT('h80)
	) name1178 (
		\shift_data_reg[70]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1420_
	);
	LUT3 #(
		.INIT('h35)
	) name1179 (
		\shift_data_reg[70]/NET0131 ,
		\wb_dat_i[6]_pad ,
		\wb_sel_i[0]_pad ,
		_w1421_
	);
	LUT3 #(
		.INIT('h08)
	) name1180 (
		_w585_,
		_w1057_,
		_w1421_,
		_w1422_
	);
	LUT4 #(
		.INIT('h8000)
	) name1181 (
		_w1032_,
		_w1297_,
		_w1350_,
		_w1370_,
		_w1423_
	);
	LUT3 #(
		.INIT('hc8)
	) name1182 (
		\shift_data_reg[70]/NET0131 ,
		_w1354_,
		_w1423_,
		_w1424_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1183 (
		_w1165_,
		_w1262_,
		_w1423_,
		_w1424_,
		_w1425_
	);
	LUT4 #(
		.INIT('hdddc)
	) name1184 (
		_w1346_,
		_w1420_,
		_w1422_,
		_w1425_,
		_w1426_
	);
	LUT3 #(
		.INIT('h35)
	) name1185 (
		\shift_data_reg[71]/NET0131 ,
		\wb_dat_i[7]_pad ,
		\wb_sel_i[0]_pad ,
		_w1427_
	);
	LUT3 #(
		.INIT('h08)
	) name1186 (
		_w585_,
		_w1057_,
		_w1427_,
		_w1428_
	);
	LUT4 #(
		.INIT('h0002)
	) name1187 (
		_w1032_,
		_w1042_,
		_w1049_,
		_w1052_,
		_w1429_
	);
	LUT3 #(
		.INIT('h80)
	) name1188 (
		_w1025_,
		_w1350_,
		_w1429_,
		_w1430_
	);
	LUT4 #(
		.INIT('h1555)
	) name1189 (
		\shift_data_reg[71]/NET0131 ,
		_w1025_,
		_w1350_,
		_w1429_,
		_w1431_
	);
	LUT2 #(
		.INIT('h2)
	) name1190 (
		_w1354_,
		_w1431_,
		_w1432_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1191 (
		_w1165_,
		_w1262_,
		_w1430_,
		_w1432_,
		_w1433_
	);
	LUT3 #(
		.INIT('h80)
	) name1192 (
		\shift_data_reg[71]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1434_
	);
	LUT4 #(
		.INIT('hff54)
	) name1193 (
		_w1346_,
		_w1428_,
		_w1433_,
		_w1434_,
		_w1435_
	);
	LUT3 #(
		.INIT('h35)
	) name1194 (
		\shift_data_reg[72]/NET0131 ,
		\wb_dat_i[8]_pad ,
		\wb_sel_i[1]_pad ,
		_w1436_
	);
	LUT3 #(
		.INIT('h08)
	) name1195 (
		_w585_,
		_w1057_,
		_w1436_,
		_w1437_
	);
	LUT4 #(
		.INIT('h4000)
	) name1196 (
		_w1032_,
		_w1306_,
		_w1350_,
		_w1370_,
		_w1438_
	);
	LUT3 #(
		.INIT('hc8)
	) name1197 (
		\shift_data_reg[72]/NET0131 ,
		_w1354_,
		_w1438_,
		_w1439_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1198 (
		_w1165_,
		_w1262_,
		_w1438_,
		_w1439_,
		_w1440_
	);
	LUT3 #(
		.INIT('h80)
	) name1199 (
		\shift_data_reg[72]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1441_
	);
	LUT4 #(
		.INIT('hff54)
	) name1200 (
		_w1346_,
		_w1437_,
		_w1440_,
		_w1441_,
		_w1442_
	);
	LUT3 #(
		.INIT('h35)
	) name1201 (
		\shift_data_reg[74]/NET0131 ,
		\wb_dat_i[10]_pad ,
		\wb_sel_i[1]_pad ,
		_w1443_
	);
	LUT3 #(
		.INIT('h08)
	) name1202 (
		_w585_,
		_w1057_,
		_w1443_,
		_w1444_
	);
	LUT2 #(
		.INIT('h4)
	) name1203 (
		_w1032_,
		_w1388_,
		_w1445_
	);
	LUT3 #(
		.INIT('h80)
	) name1204 (
		_w1350_,
		_w1370_,
		_w1445_,
		_w1446_
	);
	LUT4 #(
		.INIT('h1555)
	) name1205 (
		\shift_data_reg[74]/NET0131 ,
		_w1350_,
		_w1370_,
		_w1445_,
		_w1447_
	);
	LUT2 #(
		.INIT('h2)
	) name1206 (
		_w1354_,
		_w1447_,
		_w1448_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1207 (
		_w1165_,
		_w1262_,
		_w1446_,
		_w1448_,
		_w1449_
	);
	LUT3 #(
		.INIT('h80)
	) name1208 (
		\shift_data_reg[74]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1450_
	);
	LUT4 #(
		.INIT('hff54)
	) name1209 (
		_w1346_,
		_w1444_,
		_w1449_,
		_w1450_,
		_w1451_
	);
	LUT3 #(
		.INIT('h35)
	) name1210 (
		\shift_data_reg[75]/NET0131 ,
		\wb_dat_i[11]_pad ,
		\wb_sel_i[1]_pad ,
		_w1452_
	);
	LUT3 #(
		.INIT('h08)
	) name1211 (
		_w585_,
		_w1057_,
		_w1452_,
		_w1453_
	);
	LUT4 #(
		.INIT('h4000)
	) name1212 (
		_w1032_,
		_w1350_,
		_w1370_,
		_w1398_,
		_w1454_
	);
	LUT3 #(
		.INIT('hc8)
	) name1213 (
		\shift_data_reg[75]/NET0131 ,
		_w1354_,
		_w1454_,
		_w1455_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1214 (
		_w1165_,
		_w1262_,
		_w1454_,
		_w1455_,
		_w1456_
	);
	LUT3 #(
		.INIT('h80)
	) name1215 (
		\shift_data_reg[75]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1457_
	);
	LUT4 #(
		.INIT('hff54)
	) name1216 (
		_w1346_,
		_w1453_,
		_w1456_,
		_w1457_,
		_w1458_
	);
	LUT3 #(
		.INIT('h35)
	) name1217 (
		\shift_data_reg[73]/NET0131 ,
		\wb_dat_i[9]_pad ,
		\wb_sel_i[1]_pad ,
		_w1459_
	);
	LUT3 #(
		.INIT('h08)
	) name1218 (
		_w585_,
		_w1057_,
		_w1459_,
		_w1460_
	);
	LUT4 #(
		.INIT('h0001)
	) name1219 (
		_w1032_,
		_w1042_,
		_w1049_,
		_w1052_,
		_w1461_
	);
	LUT3 #(
		.INIT('h80)
	) name1220 (
		_w1350_,
		_w1352_,
		_w1461_,
		_w1462_
	);
	LUT4 #(
		.INIT('h1555)
	) name1221 (
		\shift_data_reg[73]/NET0131 ,
		_w1350_,
		_w1352_,
		_w1461_,
		_w1463_
	);
	LUT2 #(
		.INIT('h2)
	) name1222 (
		_w1354_,
		_w1463_,
		_w1464_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1223 (
		_w1165_,
		_w1262_,
		_w1462_,
		_w1464_,
		_w1465_
	);
	LUT3 #(
		.INIT('h80)
	) name1224 (
		\shift_data_reg[73]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1466_
	);
	LUT4 #(
		.INIT('hff54)
	) name1225 (
		_w1346_,
		_w1460_,
		_w1465_,
		_w1466_,
		_w1467_
	);
	LUT3 #(
		.INIT('h35)
	) name1226 (
		\shift_data_reg[76]/NET0131 ,
		\wb_dat_i[12]_pad ,
		\wb_sel_i[1]_pad ,
		_w1468_
	);
	LUT3 #(
		.INIT('h08)
	) name1227 (
		_w585_,
		_w1057_,
		_w1468_,
		_w1469_
	);
	LUT4 #(
		.INIT('h4000)
	) name1228 (
		_w1032_,
		_w1350_,
		_w1361_,
		_w1370_,
		_w1470_
	);
	LUT3 #(
		.INIT('hc8)
	) name1229 (
		\shift_data_reg[76]/NET0131 ,
		_w1354_,
		_w1470_,
		_w1471_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1230 (
		_w1165_,
		_w1262_,
		_w1470_,
		_w1471_,
		_w1472_
	);
	LUT3 #(
		.INIT('h80)
	) name1231 (
		\shift_data_reg[76]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1473_
	);
	LUT4 #(
		.INIT('hff54)
	) name1232 (
		_w1346_,
		_w1469_,
		_w1472_,
		_w1473_,
		_w1474_
	);
	LUT3 #(
		.INIT('h35)
	) name1233 (
		\shift_data_reg[77]/NET0131 ,
		\wb_dat_i[13]_pad ,
		\wb_sel_i[1]_pad ,
		_w1475_
	);
	LUT3 #(
		.INIT('h08)
	) name1234 (
		_w585_,
		_w1057_,
		_w1475_,
		_w1476_
	);
	LUT4 #(
		.INIT('h4000)
	) name1235 (
		_w1032_,
		_w1277_,
		_w1350_,
		_w1370_,
		_w1477_
	);
	LUT3 #(
		.INIT('hc8)
	) name1236 (
		\shift_data_reg[77]/NET0131 ,
		_w1354_,
		_w1477_,
		_w1478_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1237 (
		_w1165_,
		_w1262_,
		_w1477_,
		_w1478_,
		_w1479_
	);
	LUT3 #(
		.INIT('h80)
	) name1238 (
		\shift_data_reg[77]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1480_
	);
	LUT4 #(
		.INIT('hff54)
	) name1239 (
		_w1346_,
		_w1476_,
		_w1479_,
		_w1480_,
		_w1481_
	);
	LUT3 #(
		.INIT('h35)
	) name1240 (
		\shift_data_reg[78]/NET0131 ,
		\wb_dat_i[14]_pad ,
		\wb_sel_i[1]_pad ,
		_w1482_
	);
	LUT3 #(
		.INIT('h08)
	) name1241 (
		_w585_,
		_w1057_,
		_w1482_,
		_w1483_
	);
	LUT4 #(
		.INIT('h4000)
	) name1242 (
		_w1032_,
		_w1297_,
		_w1350_,
		_w1370_,
		_w1484_
	);
	LUT3 #(
		.INIT('hc8)
	) name1243 (
		\shift_data_reg[78]/NET0131 ,
		_w1354_,
		_w1484_,
		_w1485_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1244 (
		_w1165_,
		_w1262_,
		_w1484_,
		_w1485_,
		_w1486_
	);
	LUT3 #(
		.INIT('h80)
	) name1245 (
		\shift_data_reg[78]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1487_
	);
	LUT4 #(
		.INIT('hff54)
	) name1246 (
		_w1346_,
		_w1483_,
		_w1486_,
		_w1487_,
		_w1488_
	);
	LUT3 #(
		.INIT('h35)
	) name1247 (
		\shift_data_reg[79]/NET0131 ,
		\wb_dat_i[15]_pad ,
		\wb_sel_i[1]_pad ,
		_w1489_
	);
	LUT3 #(
		.INIT('h08)
	) name1248 (
		_w585_,
		_w1057_,
		_w1489_,
		_w1490_
	);
	LUT2 #(
		.INIT('h2)
	) name1249 (
		_w1025_,
		_w1032_,
		_w1491_
	);
	LUT3 #(
		.INIT('h80)
	) name1250 (
		_w1350_,
		_w1370_,
		_w1491_,
		_w1492_
	);
	LUT4 #(
		.INIT('h1555)
	) name1251 (
		\shift_data_reg[79]/NET0131 ,
		_w1350_,
		_w1370_,
		_w1491_,
		_w1493_
	);
	LUT2 #(
		.INIT('h2)
	) name1252 (
		_w1354_,
		_w1493_,
		_w1494_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1253 (
		_w1165_,
		_w1262_,
		_w1492_,
		_w1494_,
		_w1495_
	);
	LUT3 #(
		.INIT('h80)
	) name1254 (
		\shift_data_reg[79]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1496_
	);
	LUT4 #(
		.INIT('hff54)
	) name1255 (
		_w1346_,
		_w1490_,
		_w1495_,
		_w1496_,
		_w1497_
	);
	LUT2 #(
		.INIT('h8)
	) name1256 (
		\wb_dat_i[17]_pad ,
		\wb_sel_i[2]_pad ,
		_w1498_
	);
	LUT3 #(
		.INIT('h35)
	) name1257 (
		\shift_data_reg[81]/NET0131 ,
		\wb_dat_i[17]_pad ,
		\wb_sel_i[2]_pad ,
		_w1499_
	);
	LUT3 #(
		.INIT('h08)
	) name1258 (
		_w585_,
		_w1057_,
		_w1499_,
		_w1500_
	);
	LUT3 #(
		.INIT('h80)
	) name1259 (
		_w1350_,
		_w1351_,
		_w1379_,
		_w1501_
	);
	LUT4 #(
		.INIT('h1555)
	) name1260 (
		\shift_data_reg[81]/NET0131 ,
		_w1350_,
		_w1351_,
		_w1379_,
		_w1502_
	);
	LUT2 #(
		.INIT('h2)
	) name1261 (
		_w1354_,
		_w1502_,
		_w1503_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1262 (
		_w1165_,
		_w1262_,
		_w1501_,
		_w1503_,
		_w1504_
	);
	LUT3 #(
		.INIT('h80)
	) name1263 (
		\shift_data_reg[81]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1505_
	);
	LUT4 #(
		.INIT('hff54)
	) name1264 (
		_w1346_,
		_w1500_,
		_w1504_,
		_w1505_,
		_w1506_
	);
	LUT3 #(
		.INIT('h80)
	) name1265 (
		\shift_data_reg[82]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1507_
	);
	LUT2 #(
		.INIT('h8)
	) name1266 (
		\wb_dat_i[18]_pad ,
		\wb_sel_i[2]_pad ,
		_w1508_
	);
	LUT3 #(
		.INIT('h35)
	) name1267 (
		\shift_data_reg[82]/NET0131 ,
		\wb_dat_i[18]_pad ,
		\wb_sel_i[2]_pad ,
		_w1509_
	);
	LUT3 #(
		.INIT('h08)
	) name1268 (
		_w585_,
		_w1057_,
		_w1509_,
		_w1510_
	);
	LUT3 #(
		.INIT('h80)
	) name1269 (
		_w1350_,
		_w1351_,
		_w1389_,
		_w1511_
	);
	LUT4 #(
		.INIT('h1555)
	) name1270 (
		\shift_data_reg[82]/NET0131 ,
		_w1350_,
		_w1351_,
		_w1389_,
		_w1512_
	);
	LUT2 #(
		.INIT('h2)
	) name1271 (
		_w1354_,
		_w1512_,
		_w1513_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1272 (
		_w1165_,
		_w1262_,
		_w1511_,
		_w1513_,
		_w1514_
	);
	LUT4 #(
		.INIT('hdddc)
	) name1273 (
		_w1346_,
		_w1507_,
		_w1510_,
		_w1514_,
		_w1515_
	);
	LUT2 #(
		.INIT('h8)
	) name1274 (
		\wb_dat_i[16]_pad ,
		\wb_sel_i[2]_pad ,
		_w1516_
	);
	LUT3 #(
		.INIT('h35)
	) name1275 (
		\shift_data_reg[80]/NET0131 ,
		\wb_dat_i[16]_pad ,
		\wb_sel_i[2]_pad ,
		_w1517_
	);
	LUT3 #(
		.INIT('h08)
	) name1276 (
		_w585_,
		_w1057_,
		_w1517_,
		_w1518_
	);
	LUT4 #(
		.INIT('h8000)
	) name1277 (
		_w1032_,
		_w1306_,
		_w1350_,
		_w1351_,
		_w1519_
	);
	LUT3 #(
		.INIT('hc8)
	) name1278 (
		\shift_data_reg[80]/NET0131 ,
		_w1354_,
		_w1519_,
		_w1520_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1279 (
		_w1165_,
		_w1262_,
		_w1519_,
		_w1520_,
		_w1521_
	);
	LUT3 #(
		.INIT('h80)
	) name1280 (
		\shift_data_reg[80]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1522_
	);
	LUT4 #(
		.INIT('hff54)
	) name1281 (
		_w1346_,
		_w1518_,
		_w1521_,
		_w1522_,
		_w1523_
	);
	LUT2 #(
		.INIT('h8)
	) name1282 (
		\wb_dat_i[19]_pad ,
		\wb_sel_i[2]_pad ,
		_w1524_
	);
	LUT3 #(
		.INIT('h35)
	) name1283 (
		\shift_data_reg[83]/NET0131 ,
		\wb_dat_i[19]_pad ,
		\wb_sel_i[2]_pad ,
		_w1525_
	);
	LUT3 #(
		.INIT('h08)
	) name1284 (
		_w585_,
		_w1057_,
		_w1525_,
		_w1526_
	);
	LUT4 #(
		.INIT('h8000)
	) name1285 (
		_w1032_,
		_w1350_,
		_w1351_,
		_w1398_,
		_w1527_
	);
	LUT3 #(
		.INIT('hc8)
	) name1286 (
		\shift_data_reg[83]/NET0131 ,
		_w1354_,
		_w1527_,
		_w1528_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1287 (
		_w1165_,
		_w1262_,
		_w1527_,
		_w1528_,
		_w1529_
	);
	LUT3 #(
		.INIT('h80)
	) name1288 (
		\shift_data_reg[83]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1530_
	);
	LUT4 #(
		.INIT('hff54)
	) name1289 (
		_w1346_,
		_w1526_,
		_w1529_,
		_w1530_,
		_w1531_
	);
	LUT2 #(
		.INIT('h8)
	) name1290 (
		\wb_dat_i[20]_pad ,
		\wb_sel_i[2]_pad ,
		_w1532_
	);
	LUT3 #(
		.INIT('h35)
	) name1291 (
		\shift_data_reg[84]/NET0131 ,
		\wb_dat_i[20]_pad ,
		\wb_sel_i[2]_pad ,
		_w1533_
	);
	LUT3 #(
		.INIT('h08)
	) name1292 (
		_w585_,
		_w1057_,
		_w1533_,
		_w1534_
	);
	LUT3 #(
		.INIT('h80)
	) name1293 (
		_w1350_,
		_w1351_,
		_w1406_,
		_w1535_
	);
	LUT4 #(
		.INIT('h1555)
	) name1294 (
		\shift_data_reg[84]/NET0131 ,
		_w1350_,
		_w1351_,
		_w1406_,
		_w1536_
	);
	LUT2 #(
		.INIT('h2)
	) name1295 (
		_w1354_,
		_w1536_,
		_w1537_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1296 (
		_w1165_,
		_w1262_,
		_w1535_,
		_w1537_,
		_w1538_
	);
	LUT3 #(
		.INIT('h80)
	) name1297 (
		\shift_data_reg[84]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1539_
	);
	LUT4 #(
		.INIT('hff54)
	) name1298 (
		_w1346_,
		_w1534_,
		_w1538_,
		_w1539_,
		_w1540_
	);
	LUT2 #(
		.INIT('h8)
	) name1299 (
		\wb_dat_i[21]_pad ,
		\wb_sel_i[2]_pad ,
		_w1541_
	);
	LUT3 #(
		.INIT('h35)
	) name1300 (
		\shift_data_reg[85]/NET0131 ,
		\wb_dat_i[21]_pad ,
		\wb_sel_i[2]_pad ,
		_w1542_
	);
	LUT3 #(
		.INIT('h08)
	) name1301 (
		_w585_,
		_w1057_,
		_w1542_,
		_w1543_
	);
	LUT4 #(
		.INIT('h8000)
	) name1302 (
		_w1032_,
		_w1277_,
		_w1350_,
		_w1351_,
		_w1544_
	);
	LUT3 #(
		.INIT('hc8)
	) name1303 (
		\shift_data_reg[85]/NET0131 ,
		_w1354_,
		_w1544_,
		_w1545_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1304 (
		_w1165_,
		_w1262_,
		_w1544_,
		_w1545_,
		_w1546_
	);
	LUT3 #(
		.INIT('h80)
	) name1305 (
		\shift_data_reg[85]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1547_
	);
	LUT4 #(
		.INIT('hff54)
	) name1306 (
		_w1346_,
		_w1543_,
		_w1546_,
		_w1547_,
		_w1548_
	);
	LUT2 #(
		.INIT('h8)
	) name1307 (
		\wb_dat_i[22]_pad ,
		\wb_sel_i[2]_pad ,
		_w1549_
	);
	LUT3 #(
		.INIT('h35)
	) name1308 (
		\shift_data_reg[86]/NET0131 ,
		\wb_dat_i[22]_pad ,
		\wb_sel_i[2]_pad ,
		_w1550_
	);
	LUT3 #(
		.INIT('h08)
	) name1309 (
		_w585_,
		_w1057_,
		_w1550_,
		_w1551_
	);
	LUT4 #(
		.INIT('h8000)
	) name1310 (
		_w1032_,
		_w1297_,
		_w1350_,
		_w1351_,
		_w1552_
	);
	LUT3 #(
		.INIT('hc8)
	) name1311 (
		\shift_data_reg[86]/NET0131 ,
		_w1354_,
		_w1552_,
		_w1553_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1312 (
		_w1165_,
		_w1262_,
		_w1552_,
		_w1553_,
		_w1554_
	);
	LUT3 #(
		.INIT('h80)
	) name1313 (
		\shift_data_reg[86]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1555_
	);
	LUT4 #(
		.INIT('hff54)
	) name1314 (
		_w1346_,
		_w1551_,
		_w1554_,
		_w1555_,
		_w1556_
	);
	LUT3 #(
		.INIT('h35)
	) name1315 (
		\shift_data_reg[88]/NET0131 ,
		\wb_dat_i[24]_pad ,
		\wb_sel_i[3]_pad ,
		_w1557_
	);
	LUT3 #(
		.INIT('h08)
	) name1316 (
		_w585_,
		_w1057_,
		_w1557_,
		_w1558_
	);
	LUT4 #(
		.INIT('h4000)
	) name1317 (
		_w1032_,
		_w1306_,
		_w1350_,
		_w1351_,
		_w1559_
	);
	LUT3 #(
		.INIT('hc8)
	) name1318 (
		\shift_data_reg[88]/NET0131 ,
		_w1354_,
		_w1559_,
		_w1560_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1319 (
		_w1165_,
		_w1262_,
		_w1559_,
		_w1560_,
		_w1561_
	);
	LUT3 #(
		.INIT('h80)
	) name1320 (
		\shift_data_reg[88]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1562_
	);
	LUT4 #(
		.INIT('hff54)
	) name1321 (
		_w1346_,
		_w1558_,
		_w1561_,
		_w1562_,
		_w1563_
	);
	LUT3 #(
		.INIT('h35)
	) name1322 (
		\shift_data_reg[87]/NET0131 ,
		\wb_dat_i[23]_pad ,
		\wb_sel_i[2]_pad ,
		_w1564_
	);
	LUT3 #(
		.INIT('h08)
	) name1323 (
		_w585_,
		_w1057_,
		_w1564_,
		_w1565_
	);
	LUT3 #(
		.INIT('h80)
	) name1324 (
		_w1033_,
		_w1350_,
		_w1351_,
		_w1566_
	);
	LUT4 #(
		.INIT('h1555)
	) name1325 (
		\shift_data_reg[87]/NET0131 ,
		_w1033_,
		_w1350_,
		_w1351_,
		_w1567_
	);
	LUT2 #(
		.INIT('h2)
	) name1326 (
		_w1354_,
		_w1567_,
		_w1568_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1327 (
		_w1165_,
		_w1262_,
		_w1566_,
		_w1568_,
		_w1569_
	);
	LUT3 #(
		.INIT('h80)
	) name1328 (
		\shift_data_reg[87]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1570_
	);
	LUT4 #(
		.INIT('hff54)
	) name1329 (
		_w1346_,
		_w1565_,
		_w1569_,
		_w1570_,
		_w1571_
	);
	LUT2 #(
		.INIT('h8)
	) name1330 (
		\wb_dat_i[26]_pad ,
		\wb_sel_i[3]_pad ,
		_w1572_
	);
	LUT3 #(
		.INIT('h35)
	) name1331 (
		\shift_data_reg[90]/NET0131 ,
		\wb_dat_i[26]_pad ,
		\wb_sel_i[3]_pad ,
		_w1573_
	);
	LUT3 #(
		.INIT('h08)
	) name1332 (
		_w585_,
		_w1057_,
		_w1573_,
		_w1574_
	);
	LUT4 #(
		.INIT('h4000)
	) name1333 (
		_w1032_,
		_w1350_,
		_w1351_,
		_w1388_,
		_w1575_
	);
	LUT3 #(
		.INIT('hc8)
	) name1334 (
		\shift_data_reg[90]/NET0131 ,
		_w1354_,
		_w1575_,
		_w1576_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1335 (
		_w1165_,
		_w1262_,
		_w1575_,
		_w1576_,
		_w1577_
	);
	LUT3 #(
		.INIT('h80)
	) name1336 (
		\shift_data_reg[90]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1578_
	);
	LUT4 #(
		.INIT('hff54)
	) name1337 (
		_w1346_,
		_w1574_,
		_w1577_,
		_w1578_,
		_w1579_
	);
	LUT2 #(
		.INIT('h8)
	) name1338 (
		\wb_dat_i[27]_pad ,
		\wb_sel_i[3]_pad ,
		_w1580_
	);
	LUT3 #(
		.INIT('h35)
	) name1339 (
		\shift_data_reg[91]/NET0131 ,
		\wb_dat_i[27]_pad ,
		\wb_sel_i[3]_pad ,
		_w1581_
	);
	LUT3 #(
		.INIT('h08)
	) name1340 (
		_w585_,
		_w1057_,
		_w1581_,
		_w1582_
	);
	LUT4 #(
		.INIT('h4000)
	) name1341 (
		_w1032_,
		_w1350_,
		_w1351_,
		_w1398_,
		_w1583_
	);
	LUT3 #(
		.INIT('hc8)
	) name1342 (
		\shift_data_reg[91]/NET0131 ,
		_w1354_,
		_w1583_,
		_w1584_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1343 (
		_w1165_,
		_w1262_,
		_w1583_,
		_w1584_,
		_w1585_
	);
	LUT3 #(
		.INIT('h80)
	) name1344 (
		\shift_data_reg[91]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1586_
	);
	LUT4 #(
		.INIT('hff54)
	) name1345 (
		_w1346_,
		_w1582_,
		_w1585_,
		_w1586_,
		_w1587_
	);
	LUT2 #(
		.INIT('h8)
	) name1346 (
		\wb_dat_i[29]_pad ,
		\wb_sel_i[3]_pad ,
		_w1588_
	);
	LUT3 #(
		.INIT('h35)
	) name1347 (
		\shift_data_reg[93]/NET0131 ,
		\wb_dat_i[29]_pad ,
		\wb_sel_i[3]_pad ,
		_w1589_
	);
	LUT3 #(
		.INIT('h08)
	) name1348 (
		_w585_,
		_w1057_,
		_w1589_,
		_w1590_
	);
	LUT4 #(
		.INIT('h4000)
	) name1349 (
		_w1032_,
		_w1277_,
		_w1350_,
		_w1351_,
		_w1591_
	);
	LUT3 #(
		.INIT('hc8)
	) name1350 (
		\shift_data_reg[93]/NET0131 ,
		_w1354_,
		_w1591_,
		_w1592_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1351 (
		_w1165_,
		_w1262_,
		_w1591_,
		_w1592_,
		_w1593_
	);
	LUT3 #(
		.INIT('h80)
	) name1352 (
		\shift_data_reg[93]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1594_
	);
	LUT4 #(
		.INIT('hff54)
	) name1353 (
		_w1346_,
		_w1590_,
		_w1593_,
		_w1594_,
		_w1595_
	);
	LUT2 #(
		.INIT('h8)
	) name1354 (
		\wb_dat_i[30]_pad ,
		\wb_sel_i[3]_pad ,
		_w1596_
	);
	LUT3 #(
		.INIT('h35)
	) name1355 (
		\shift_data_reg[94]/NET0131 ,
		\wb_dat_i[30]_pad ,
		\wb_sel_i[3]_pad ,
		_w1597_
	);
	LUT3 #(
		.INIT('h08)
	) name1356 (
		_w585_,
		_w1057_,
		_w1597_,
		_w1598_
	);
	LUT4 #(
		.INIT('h4000)
	) name1357 (
		_w1032_,
		_w1297_,
		_w1350_,
		_w1351_,
		_w1599_
	);
	LUT3 #(
		.INIT('hc8)
	) name1358 (
		\shift_data_reg[94]/NET0131 ,
		_w1354_,
		_w1599_,
		_w1600_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1359 (
		_w1165_,
		_w1262_,
		_w1599_,
		_w1600_,
		_w1601_
	);
	LUT3 #(
		.INIT('h80)
	) name1360 (
		\shift_data_reg[94]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1602_
	);
	LUT4 #(
		.INIT('hff54)
	) name1361 (
		_w1346_,
		_w1598_,
		_w1601_,
		_w1602_,
		_w1603_
	);
	LUT3 #(
		.INIT('h35)
	) name1362 (
		\shift_data_reg[95]/NET0131 ,
		\wb_dat_i[31]_pad ,
		\wb_sel_i[3]_pad ,
		_w1604_
	);
	LUT3 #(
		.INIT('h08)
	) name1363 (
		_w585_,
		_w1057_,
		_w1604_,
		_w1605_
	);
	LUT3 #(
		.INIT('h80)
	) name1364 (
		_w1350_,
		_w1351_,
		_w1491_,
		_w1606_
	);
	LUT4 #(
		.INIT('h1555)
	) name1365 (
		\shift_data_reg[95]/NET0131 ,
		_w1350_,
		_w1351_,
		_w1491_,
		_w1607_
	);
	LUT2 #(
		.INIT('h2)
	) name1366 (
		_w1354_,
		_w1607_,
		_w1608_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1367 (
		_w1165_,
		_w1262_,
		_w1606_,
		_w1608_,
		_w1609_
	);
	LUT3 #(
		.INIT('h80)
	) name1368 (
		\shift_data_reg[95]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1610_
	);
	LUT4 #(
		.INIT('hff54)
	) name1369 (
		_w1346_,
		_w1605_,
		_w1609_,
		_w1610_,
		_w1611_
	);
	LUT3 #(
		.INIT('h35)
	) name1370 (
		\shift_data_reg[25]/NET0131 ,
		\wb_dat_i[25]_pad ,
		\wb_sel_i[3]_pad ,
		_w1612_
	);
	LUT4 #(
		.INIT('h0040)
	) name1371 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1612_,
		_w1613_
	);
	LUT2 #(
		.INIT('h4)
	) name1372 (
		_w1268_,
		_w1060_,
		_w1614_
	);
	LUT4 #(
		.INIT('h4000)
	) name1373 (
		_w1032_,
		_w1065_,
		_w1351_,
		_w1614_,
		_w1615_
	);
	LUT2 #(
		.INIT('h8)
	) name1374 (
		_w1352_,
		_w1615_,
		_w1616_
	);
	LUT4 #(
		.INIT('h3222)
	) name1375 (
		\shift_data_reg[25]/NET0131 ,
		_w1346_,
		_w1352_,
		_w1615_,
		_w1617_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1376 (
		_w1165_,
		_w1262_,
		_w1616_,
		_w1617_,
		_w1618_
	);
	LUT2 #(
		.INIT('he)
	) name1377 (
		_w1613_,
		_w1618_,
		_w1619_
	);
	LUT3 #(
		.INIT('h35)
	) name1378 (
		\shift_data_reg[27]/NET0131 ,
		\wb_dat_i[27]_pad ,
		\wb_sel_i[3]_pad ,
		_w1620_
	);
	LUT4 #(
		.INIT('h0040)
	) name1379 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1620_,
		_w1621_
	);
	LUT2 #(
		.INIT('h8)
	) name1380 (
		_w1398_,
		_w1615_,
		_w1622_
	);
	LUT4 #(
		.INIT('h3222)
	) name1381 (
		\shift_data_reg[27]/NET0131 ,
		_w1346_,
		_w1398_,
		_w1615_,
		_w1623_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1382 (
		_w1165_,
		_w1262_,
		_w1622_,
		_w1623_,
		_w1624_
	);
	LUT2 #(
		.INIT('he)
	) name1383 (
		_w1621_,
		_w1624_,
		_w1625_
	);
	LUT3 #(
		.INIT('h35)
	) name1384 (
		\shift_data_reg[26]/NET0131 ,
		\wb_dat_i[26]_pad ,
		\wb_sel_i[3]_pad ,
		_w1626_
	);
	LUT4 #(
		.INIT('h0040)
	) name1385 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1626_,
		_w1627_
	);
	LUT4 #(
		.INIT('h8000)
	) name1386 (
		_w1065_,
		_w1351_,
		_w1445_,
		_w1614_,
		_w1628_
	);
	LUT3 #(
		.INIT('h32)
	) name1387 (
		\shift_data_reg[26]/NET0131 ,
		_w1346_,
		_w1628_,
		_w1629_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1388 (
		_w1165_,
		_w1262_,
		_w1628_,
		_w1629_,
		_w1630_
	);
	LUT2 #(
		.INIT('he)
	) name1389 (
		_w1627_,
		_w1630_,
		_w1631_
	);
	LUT3 #(
		.INIT('h35)
	) name1390 (
		\shift_data_reg[28]/NET0131 ,
		\wb_dat_i[28]_pad ,
		\wb_sel_i[3]_pad ,
		_w1632_
	);
	LUT4 #(
		.INIT('h0040)
	) name1391 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1632_,
		_w1633_
	);
	LUT2 #(
		.INIT('h8)
	) name1392 (
		_w1361_,
		_w1615_,
		_w1634_
	);
	LUT4 #(
		.INIT('h3222)
	) name1393 (
		\shift_data_reg[28]/NET0131 ,
		_w1346_,
		_w1361_,
		_w1615_,
		_w1635_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1394 (
		_w1165_,
		_w1262_,
		_w1634_,
		_w1635_,
		_w1636_
	);
	LUT2 #(
		.INIT('he)
	) name1395 (
		_w1633_,
		_w1636_,
		_w1637_
	);
	LUT3 #(
		.INIT('h35)
	) name1396 (
		\shift_data_reg[29]/NET0131 ,
		\wb_dat_i[29]_pad ,
		\wb_sel_i[3]_pad ,
		_w1638_
	);
	LUT4 #(
		.INIT('h0040)
	) name1397 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1638_,
		_w1639_
	);
	LUT2 #(
		.INIT('h8)
	) name1398 (
		_w1277_,
		_w1615_,
		_w1640_
	);
	LUT4 #(
		.INIT('h0e0a)
	) name1399 (
		\shift_data_reg[29]/NET0131 ,
		_w1277_,
		_w1346_,
		_w1615_,
		_w1641_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1400 (
		_w1165_,
		_w1262_,
		_w1640_,
		_w1641_,
		_w1642_
	);
	LUT2 #(
		.INIT('he)
	) name1401 (
		_w1639_,
		_w1642_,
		_w1643_
	);
	LUT3 #(
		.INIT('h35)
	) name1402 (
		\shift_data_reg[2]/NET0131 ,
		\wb_dat_i[2]_pad ,
		\wb_sel_i[0]_pad ,
		_w1644_
	);
	LUT4 #(
		.INIT('h0040)
	) name1403 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1644_,
		_w1645_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name1404 (
		\shift_data_reg[2]/NET0131 ,
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1646_
	);
	LUT3 #(
		.INIT('h0b)
	) name1405 (
		_w1264_,
		_w1060_,
		_w1646_,
		_w1647_
	);
	LUT3 #(
		.INIT('h80)
	) name1406 (
		_w1065_,
		_w1388_,
		_w1429_,
		_w1648_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1407 (
		\shift_data_reg[2]/NET0131 ,
		_w1065_,
		_w1388_,
		_w1429_,
		_w1649_
	);
	LUT2 #(
		.INIT('h2)
	) name1408 (
		_w1614_,
		_w1649_,
		_w1650_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1409 (
		_w1165_,
		_w1262_,
		_w1648_,
		_w1650_,
		_w1651_
	);
	LUT3 #(
		.INIT('hab)
	) name1410 (
		_w1645_,
		_w1647_,
		_w1651_,
		_w1652_
	);
	LUT3 #(
		.INIT('h35)
	) name1411 (
		\shift_data_reg[30]/NET0131 ,
		\wb_dat_i[30]_pad ,
		\wb_sel_i[3]_pad ,
		_w1653_
	);
	LUT4 #(
		.INIT('h0040)
	) name1412 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1653_,
		_w1654_
	);
	LUT2 #(
		.INIT('h8)
	) name1413 (
		_w1297_,
		_w1615_,
		_w1655_
	);
	LUT4 #(
		.INIT('h0e0a)
	) name1414 (
		\shift_data_reg[30]/NET0131 ,
		_w1297_,
		_w1346_,
		_w1615_,
		_w1656_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1415 (
		_w1165_,
		_w1262_,
		_w1655_,
		_w1656_,
		_w1657_
	);
	LUT2 #(
		.INIT('he)
	) name1416 (
		_w1654_,
		_w1657_,
		_w1658_
	);
	LUT3 #(
		.INIT('h35)
	) name1417 (
		\shift_data_reg[31]/NET0131 ,
		\wb_dat_i[31]_pad ,
		\wb_sel_i[3]_pad ,
		_w1659_
	);
	LUT4 #(
		.INIT('h0040)
	) name1418 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1659_,
		_w1660_
	);
	LUT2 #(
		.INIT('h8)
	) name1419 (
		_w1025_,
		_w1615_,
		_w1661_
	);
	LUT4 #(
		.INIT('h0e0a)
	) name1420 (
		\shift_data_reg[31]/NET0131 ,
		_w1025_,
		_w1346_,
		_w1615_,
		_w1662_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1421 (
		_w1165_,
		_w1262_,
		_w1661_,
		_w1662_,
		_w1663_
	);
	LUT2 #(
		.INIT('he)
	) name1422 (
		_w1660_,
		_w1663_,
		_w1664_
	);
	LUT3 #(
		.INIT('h35)
	) name1423 (
		\shift_data_reg[3]/NET0131 ,
		\wb_dat_i[3]_pad ,
		\wb_sel_i[0]_pad ,
		_w1665_
	);
	LUT4 #(
		.INIT('h0040)
	) name1424 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1665_,
		_w1666_
	);
	LUT3 #(
		.INIT('h10)
	) name1425 (
		_w1062_,
		_w1064_,
		_w1614_,
		_w1667_
	);
	LUT4 #(
		.INIT('h1000)
	) name1426 (
		_w1062_,
		_w1064_,
		_w1398_,
		_w1614_,
		_w1668_
	);
	LUT2 #(
		.INIT('h8)
	) name1427 (
		_w1429_,
		_w1668_,
		_w1669_
	);
	LUT4 #(
		.INIT('h3222)
	) name1428 (
		\shift_data_reg[3]/NET0131 ,
		_w1346_,
		_w1429_,
		_w1668_,
		_w1670_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1429 (
		_w1165_,
		_w1262_,
		_w1669_,
		_w1670_,
		_w1671_
	);
	LUT2 #(
		.INIT('he)
	) name1430 (
		_w1666_,
		_w1671_,
		_w1672_
	);
	LUT3 #(
		.INIT('h35)
	) name1431 (
		\shift_data_reg[4]/NET0131 ,
		\wb_dat_i[4]_pad ,
		\wb_sel_i[0]_pad ,
		_w1673_
	);
	LUT4 #(
		.INIT('h0040)
	) name1432 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1673_,
		_w1674_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name1433 (
		\shift_data_reg[4]/NET0131 ,
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1675_
	);
	LUT3 #(
		.INIT('h0b)
	) name1434 (
		_w1264_,
		_w1060_,
		_w1675_,
		_w1676_
	);
	LUT3 #(
		.INIT('h80)
	) name1435 (
		_w1065_,
		_w1361_,
		_w1429_,
		_w1677_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1436 (
		\shift_data_reg[4]/NET0131 ,
		_w1065_,
		_w1361_,
		_w1429_,
		_w1678_
	);
	LUT2 #(
		.INIT('h2)
	) name1437 (
		_w1614_,
		_w1678_,
		_w1679_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1438 (
		_w1165_,
		_w1262_,
		_w1677_,
		_w1679_,
		_w1680_
	);
	LUT3 #(
		.INIT('hab)
	) name1439 (
		_w1674_,
		_w1676_,
		_w1680_,
		_w1681_
	);
	LUT3 #(
		.INIT('h35)
	) name1440 (
		\shift_data_reg[5]/NET0131 ,
		\wb_dat_i[5]_pad ,
		\wb_sel_i[0]_pad ,
		_w1682_
	);
	LUT4 #(
		.INIT('h0040)
	) name1441 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1682_,
		_w1683_
	);
	LUT3 #(
		.INIT('h80)
	) name1442 (
		_w1024_,
		_w1276_,
		_w1614_,
		_w1684_
	);
	LUT3 #(
		.INIT('h80)
	) name1443 (
		_w1065_,
		_w1429_,
		_w1684_,
		_w1685_
	);
	LUT4 #(
		.INIT('h1555)
	) name1444 (
		\shift_data_reg[5]/NET0131 ,
		_w1065_,
		_w1429_,
		_w1684_,
		_w1686_
	);
	LUT2 #(
		.INIT('h1)
	) name1445 (
		_w1346_,
		_w1686_,
		_w1687_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1446 (
		_w1165_,
		_w1262_,
		_w1685_,
		_w1687_,
		_w1688_
	);
	LUT2 #(
		.INIT('he)
	) name1447 (
		_w1683_,
		_w1688_,
		_w1689_
	);
	LUT3 #(
		.INIT('h35)
	) name1448 (
		\shift_data_reg[6]/NET0131 ,
		\wb_dat_i[6]_pad ,
		\wb_sel_i[0]_pad ,
		_w1690_
	);
	LUT4 #(
		.INIT('h0040)
	) name1449 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1690_,
		_w1691_
	);
	LUT3 #(
		.INIT('h80)
	) name1450 (
		_w1024_,
		_w1296_,
		_w1614_,
		_w1692_
	);
	LUT3 #(
		.INIT('h80)
	) name1451 (
		_w1065_,
		_w1429_,
		_w1692_,
		_w1693_
	);
	LUT4 #(
		.INIT('h1555)
	) name1452 (
		\shift_data_reg[6]/NET0131 ,
		_w1065_,
		_w1429_,
		_w1692_,
		_w1694_
	);
	LUT2 #(
		.INIT('h1)
	) name1453 (
		_w1346_,
		_w1694_,
		_w1695_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1454 (
		_w1165_,
		_w1262_,
		_w1693_,
		_w1695_,
		_w1696_
	);
	LUT2 #(
		.INIT('he)
	) name1455 (
		_w1691_,
		_w1696_,
		_w1697_
	);
	LUT3 #(
		.INIT('h35)
	) name1456 (
		\shift_data_reg[0]/NET0131 ,
		\wb_dat_i[0]_pad ,
		\wb_sel_i[0]_pad ,
		_w1698_
	);
	LUT4 #(
		.INIT('h0040)
	) name1457 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1698_,
		_w1699_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name1458 (
		\shift_data_reg[0]/NET0131 ,
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1700_
	);
	LUT3 #(
		.INIT('h0b)
	) name1459 (
		_w1264_,
		_w1060_,
		_w1700_,
		_w1701_
	);
	LUT3 #(
		.INIT('h80)
	) name1460 (
		_w1065_,
		_w1306_,
		_w1429_,
		_w1702_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1461 (
		\shift_data_reg[0]/NET0131 ,
		_w1065_,
		_w1306_,
		_w1429_,
		_w1703_
	);
	LUT2 #(
		.INIT('h2)
	) name1462 (
		_w1614_,
		_w1703_,
		_w1704_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1463 (
		_w1165_,
		_w1262_,
		_w1702_,
		_w1704_,
		_w1705_
	);
	LUT3 #(
		.INIT('hab)
	) name1464 (
		_w1699_,
		_w1701_,
		_w1705_,
		_w1706_
	);
	LUT3 #(
		.INIT('h35)
	) name1465 (
		\shift_data_reg[10]/NET0131 ,
		\wb_dat_i[10]_pad ,
		\wb_sel_i[1]_pad ,
		_w1707_
	);
	LUT4 #(
		.INIT('h0040)
	) name1466 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1707_,
		_w1708_
	);
	LUT2 #(
		.INIT('h8)
	) name1467 (
		\shift_data_reg[10]/NET0131 ,
		\wb_adr_i[2]_pad ,
		_w1709_
	);
	LUT3 #(
		.INIT('h08)
	) name1468 (
		_w1055_,
		_w1263_,
		_w1709_,
		_w1710_
	);
	LUT3 #(
		.INIT('h80)
	) name1469 (
		_w1065_,
		_w1388_,
		_w1461_,
		_w1711_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1470 (
		_w1060_,
		_w1165_,
		_w1262_,
		_w1711_,
		_w1712_
	);
	LUT4 #(
		.INIT('h8000)
	) name1471 (
		_w1065_,
		_w1388_,
		_w1461_,
		_w1614_,
		_w1713_
	);
	LUT2 #(
		.INIT('h2)
	) name1472 (
		\shift_data_reg[10]/NET0131 ,
		_w1713_,
		_w1714_
	);
	LUT4 #(
		.INIT('hbbba)
	) name1473 (
		_w1708_,
		_w1710_,
		_w1712_,
		_w1714_,
		_w1715_
	);
	LUT3 #(
		.INIT('h35)
	) name1474 (
		\shift_data_reg[7]/NET0131 ,
		\wb_dat_i[7]_pad ,
		\wb_sel_i[0]_pad ,
		_w1716_
	);
	LUT4 #(
		.INIT('h0040)
	) name1475 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1716_,
		_w1717_
	);
	LUT3 #(
		.INIT('h80)
	) name1476 (
		_w1025_,
		_w1429_,
		_w1667_,
		_w1718_
	);
	LUT4 #(
		.INIT('h1555)
	) name1477 (
		\shift_data_reg[7]/NET0131 ,
		_w1025_,
		_w1429_,
		_w1667_,
		_w1719_
	);
	LUT2 #(
		.INIT('h1)
	) name1478 (
		_w1346_,
		_w1719_,
		_w1720_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1479 (
		_w1165_,
		_w1262_,
		_w1718_,
		_w1720_,
		_w1721_
	);
	LUT2 #(
		.INIT('he)
	) name1480 (
		_w1717_,
		_w1721_,
		_w1722_
	);
	LUT3 #(
		.INIT('h35)
	) name1481 (
		\shift_data_reg[11]/NET0131 ,
		\wb_dat_i[11]_pad ,
		\wb_sel_i[1]_pad ,
		_w1723_
	);
	LUT4 #(
		.INIT('h0040)
	) name1482 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1723_,
		_w1724_
	);
	LUT2 #(
		.INIT('h8)
	) name1483 (
		_w1461_,
		_w1668_,
		_w1725_
	);
	LUT4 #(
		.INIT('h3222)
	) name1484 (
		\shift_data_reg[11]/NET0131 ,
		_w1346_,
		_w1461_,
		_w1668_,
		_w1726_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1485 (
		_w1165_,
		_w1262_,
		_w1725_,
		_w1726_,
		_w1727_
	);
	LUT2 #(
		.INIT('he)
	) name1486 (
		_w1724_,
		_w1727_,
		_w1728_
	);
	LUT3 #(
		.INIT('h35)
	) name1487 (
		\shift_data_reg[8]/NET0131 ,
		\wb_dat_i[8]_pad ,
		\wb_sel_i[1]_pad ,
		_w1729_
	);
	LUT4 #(
		.INIT('h0040)
	) name1488 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1729_,
		_w1730_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name1489 (
		\shift_data_reg[8]/NET0131 ,
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1731_
	);
	LUT3 #(
		.INIT('h0b)
	) name1490 (
		_w1264_,
		_w1060_,
		_w1731_,
		_w1732_
	);
	LUT3 #(
		.INIT('h80)
	) name1491 (
		_w1065_,
		_w1306_,
		_w1461_,
		_w1733_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1492 (
		\shift_data_reg[8]/NET0131 ,
		_w1065_,
		_w1306_,
		_w1461_,
		_w1734_
	);
	LUT2 #(
		.INIT('h2)
	) name1493 (
		_w1614_,
		_w1734_,
		_w1735_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1494 (
		_w1165_,
		_w1262_,
		_w1733_,
		_w1735_,
		_w1736_
	);
	LUT3 #(
		.INIT('hab)
	) name1495 (
		_w1730_,
		_w1732_,
		_w1736_,
		_w1737_
	);
	LUT3 #(
		.INIT('h35)
	) name1496 (
		\shift_data_reg[9]/NET0131 ,
		\wb_dat_i[9]_pad ,
		\wb_sel_i[1]_pad ,
		_w1738_
	);
	LUT4 #(
		.INIT('h0040)
	) name1497 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1738_,
		_w1739_
	);
	LUT3 #(
		.INIT('h80)
	) name1498 (
		_w1352_,
		_w1461_,
		_w1667_,
		_w1740_
	);
	LUT4 #(
		.INIT('h1555)
	) name1499 (
		\shift_data_reg[9]/NET0131 ,
		_w1352_,
		_w1461_,
		_w1667_,
		_w1741_
	);
	LUT2 #(
		.INIT('h1)
	) name1500 (
		_w1346_,
		_w1741_,
		_w1742_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1501 (
		_w1165_,
		_w1262_,
		_w1740_,
		_w1742_,
		_w1743_
	);
	LUT2 #(
		.INIT('he)
	) name1502 (
		_w1739_,
		_w1743_,
		_w1744_
	);
	LUT3 #(
		.INIT('h35)
	) name1503 (
		\shift_data_reg[12]/NET0131 ,
		\wb_dat_i[12]_pad ,
		\wb_sel_i[1]_pad ,
		_w1745_
	);
	LUT4 #(
		.INIT('h0040)
	) name1504 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1745_,
		_w1746_
	);
	LUT2 #(
		.INIT('h8)
	) name1505 (
		\shift_data_reg[12]/NET0131 ,
		\wb_adr_i[2]_pad ,
		_w1747_
	);
	LUT3 #(
		.INIT('h08)
	) name1506 (
		_w1055_,
		_w1263_,
		_w1747_,
		_w1748_
	);
	LUT3 #(
		.INIT('h80)
	) name1507 (
		_w1065_,
		_w1361_,
		_w1461_,
		_w1749_
	);
	LUT4 #(
		.INIT('h8000)
	) name1508 (
		_w1065_,
		_w1361_,
		_w1461_,
		_w1614_,
		_w1750_
	);
	LUT2 #(
		.INIT('h2)
	) name1509 (
		\shift_data_reg[12]/NET0131 ,
		_w1750_,
		_w1751_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1510 (
		_w1060_,
		_w1165_,
		_w1262_,
		_w1749_,
		_w1752_
	);
	LUT4 #(
		.INIT('hbbba)
	) name1511 (
		_w1746_,
		_w1748_,
		_w1751_,
		_w1752_,
		_w1753_
	);
	LUT3 #(
		.INIT('h35)
	) name1512 (
		\shift_data_reg[14]/NET0131 ,
		\wb_dat_i[14]_pad ,
		\wb_sel_i[1]_pad ,
		_w1754_
	);
	LUT4 #(
		.INIT('h0040)
	) name1513 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1754_,
		_w1755_
	);
	LUT3 #(
		.INIT('h80)
	) name1514 (
		_w1065_,
		_w1461_,
		_w1692_,
		_w1756_
	);
	LUT4 #(
		.INIT('h1555)
	) name1515 (
		\shift_data_reg[14]/NET0131 ,
		_w1065_,
		_w1461_,
		_w1692_,
		_w1757_
	);
	LUT2 #(
		.INIT('h1)
	) name1516 (
		_w1346_,
		_w1757_,
		_w1758_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1517 (
		_w1165_,
		_w1262_,
		_w1756_,
		_w1758_,
		_w1759_
	);
	LUT2 #(
		.INIT('he)
	) name1518 (
		_w1755_,
		_w1759_,
		_w1760_
	);
	LUT3 #(
		.INIT('h35)
	) name1519 (
		\shift_data_reg[13]/NET0131 ,
		\wb_dat_i[13]_pad ,
		\wb_sel_i[1]_pad ,
		_w1761_
	);
	LUT4 #(
		.INIT('h0040)
	) name1520 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1761_,
		_w1762_
	);
	LUT3 #(
		.INIT('h80)
	) name1521 (
		_w1065_,
		_w1461_,
		_w1684_,
		_w1763_
	);
	LUT4 #(
		.INIT('h1555)
	) name1522 (
		\shift_data_reg[13]/NET0131 ,
		_w1065_,
		_w1461_,
		_w1684_,
		_w1764_
	);
	LUT2 #(
		.INIT('h1)
	) name1523 (
		_w1346_,
		_w1764_,
		_w1765_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1524 (
		_w1165_,
		_w1262_,
		_w1763_,
		_w1765_,
		_w1766_
	);
	LUT2 #(
		.INIT('he)
	) name1525 (
		_w1762_,
		_w1766_,
		_w1767_
	);
	LUT3 #(
		.INIT('h35)
	) name1526 (
		\shift_data_reg[15]/NET0131 ,
		\wb_dat_i[15]_pad ,
		\wb_sel_i[1]_pad ,
		_w1768_
	);
	LUT4 #(
		.INIT('h0040)
	) name1527 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1768_,
		_w1769_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name1528 (
		\shift_data_reg[15]/NET0131 ,
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1770_
	);
	LUT3 #(
		.INIT('h0b)
	) name1529 (
		_w1264_,
		_w1060_,
		_w1770_,
		_w1771_
	);
	LUT3 #(
		.INIT('h80)
	) name1530 (
		_w1025_,
		_w1065_,
		_w1461_,
		_w1772_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1531 (
		\shift_data_reg[15]/NET0131 ,
		_w1025_,
		_w1065_,
		_w1461_,
		_w1773_
	);
	LUT2 #(
		.INIT('h2)
	) name1532 (
		_w1614_,
		_w1773_,
		_w1774_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1533 (
		_w1165_,
		_w1262_,
		_w1772_,
		_w1774_,
		_w1775_
	);
	LUT3 #(
		.INIT('hab)
	) name1534 (
		_w1769_,
		_w1771_,
		_w1775_,
		_w1776_
	);
	LUT3 #(
		.INIT('h35)
	) name1535 (
		\shift_data_reg[16]/NET0131 ,
		\wb_dat_i[16]_pad ,
		\wb_sel_i[2]_pad ,
		_w1777_
	);
	LUT4 #(
		.INIT('h0040)
	) name1536 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1777_,
		_w1778_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name1537 (
		\shift_data_reg[16]/NET0131 ,
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1779_
	);
	LUT3 #(
		.INIT('h0b)
	) name1538 (
		_w1264_,
		_w1060_,
		_w1779_,
		_w1780_
	);
	LUT3 #(
		.INIT('h80)
	) name1539 (
		_w1065_,
		_w1351_,
		_w1369_,
		_w1781_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1540 (
		\shift_data_reg[16]/NET0131 ,
		_w1065_,
		_w1351_,
		_w1369_,
		_w1782_
	);
	LUT2 #(
		.INIT('h2)
	) name1541 (
		_w1614_,
		_w1782_,
		_w1783_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1542 (
		_w1165_,
		_w1262_,
		_w1781_,
		_w1783_,
		_w1784_
	);
	LUT3 #(
		.INIT('hab)
	) name1543 (
		_w1778_,
		_w1780_,
		_w1784_,
		_w1785_
	);
	LUT3 #(
		.INIT('h35)
	) name1544 (
		\shift_data_reg[17]/NET0131 ,
		\wb_dat_i[17]_pad ,
		\wb_sel_i[2]_pad ,
		_w1786_
	);
	LUT4 #(
		.INIT('h0040)
	) name1545 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1786_,
		_w1787_
	);
	LUT4 #(
		.INIT('h8000)
	) name1546 (
		_w1032_,
		_w1065_,
		_w1351_,
		_w1614_,
		_w1788_
	);
	LUT2 #(
		.INIT('h8)
	) name1547 (
		_w1352_,
		_w1788_,
		_w1789_
	);
	LUT4 #(
		.INIT('h3222)
	) name1548 (
		\shift_data_reg[17]/NET0131 ,
		_w1346_,
		_w1352_,
		_w1788_,
		_w1790_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1549 (
		_w1165_,
		_w1262_,
		_w1789_,
		_w1790_,
		_w1791_
	);
	LUT2 #(
		.INIT('he)
	) name1550 (
		_w1787_,
		_w1791_,
		_w1792_
	);
	LUT3 #(
		.INIT('h35)
	) name1551 (
		\shift_data_reg[18]/NET0131 ,
		\wb_dat_i[18]_pad ,
		\wb_sel_i[2]_pad ,
		_w1793_
	);
	LUT4 #(
		.INIT('h0040)
	) name1552 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1793_,
		_w1794_
	);
	LUT4 #(
		.INIT('h8000)
	) name1553 (
		_w1065_,
		_w1351_,
		_w1389_,
		_w1614_,
		_w1795_
	);
	LUT3 #(
		.INIT('h32)
	) name1554 (
		\shift_data_reg[18]/NET0131 ,
		_w1346_,
		_w1795_,
		_w1796_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1555 (
		_w1165_,
		_w1262_,
		_w1795_,
		_w1796_,
		_w1797_
	);
	LUT2 #(
		.INIT('he)
	) name1556 (
		_w1794_,
		_w1797_,
		_w1798_
	);
	LUT3 #(
		.INIT('h35)
	) name1557 (
		\shift_data_reg[19]/NET0131 ,
		\wb_dat_i[19]_pad ,
		\wb_sel_i[2]_pad ,
		_w1799_
	);
	LUT4 #(
		.INIT('h0040)
	) name1558 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1799_,
		_w1800_
	);
	LUT2 #(
		.INIT('h8)
	) name1559 (
		_w1398_,
		_w1788_,
		_w1801_
	);
	LUT4 #(
		.INIT('h3222)
	) name1560 (
		\shift_data_reg[19]/NET0131 ,
		_w1346_,
		_w1398_,
		_w1788_,
		_w1802_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1561 (
		_w1165_,
		_w1262_,
		_w1801_,
		_w1802_,
		_w1803_
	);
	LUT2 #(
		.INIT('he)
	) name1562 (
		_w1800_,
		_w1803_,
		_w1804_
	);
	LUT3 #(
		.INIT('h35)
	) name1563 (
		\shift_data_reg[1]/NET0131 ,
		\wb_dat_i[1]_pad ,
		\wb_sel_i[0]_pad ,
		_w1805_
	);
	LUT4 #(
		.INIT('h0040)
	) name1564 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1805_,
		_w1806_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name1565 (
		\shift_data_reg[1]/NET0131 ,
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1807_
	);
	LUT3 #(
		.INIT('h0b)
	) name1566 (
		_w1264_,
		_w1060_,
		_w1807_,
		_w1808_
	);
	LUT3 #(
		.INIT('h80)
	) name1567 (
		_w1065_,
		_w1352_,
		_w1429_,
		_w1809_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1568 (
		\shift_data_reg[1]/NET0131 ,
		_w1065_,
		_w1352_,
		_w1429_,
		_w1810_
	);
	LUT2 #(
		.INIT('h2)
	) name1569 (
		_w1614_,
		_w1810_,
		_w1811_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1570 (
		_w1165_,
		_w1262_,
		_w1809_,
		_w1811_,
		_w1812_
	);
	LUT3 #(
		.INIT('hab)
	) name1571 (
		_w1806_,
		_w1808_,
		_w1812_,
		_w1813_
	);
	LUT3 #(
		.INIT('h35)
	) name1572 (
		\shift_data_reg[20]/NET0131 ,
		\wb_dat_i[20]_pad ,
		\wb_sel_i[2]_pad ,
		_w1814_
	);
	LUT4 #(
		.INIT('h0040)
	) name1573 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1814_,
		_w1815_
	);
	LUT2 #(
		.INIT('h8)
	) name1574 (
		_w1361_,
		_w1788_,
		_w1816_
	);
	LUT4 #(
		.INIT('h3222)
	) name1575 (
		\shift_data_reg[20]/NET0131 ,
		_w1346_,
		_w1361_,
		_w1788_,
		_w1817_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1576 (
		_w1165_,
		_w1262_,
		_w1816_,
		_w1817_,
		_w1818_
	);
	LUT2 #(
		.INIT('he)
	) name1577 (
		_w1815_,
		_w1818_,
		_w1819_
	);
	LUT3 #(
		.INIT('h35)
	) name1578 (
		\shift_data_reg[21]/NET0131 ,
		\wb_dat_i[21]_pad ,
		\wb_sel_i[2]_pad ,
		_w1820_
	);
	LUT4 #(
		.INIT('h0040)
	) name1579 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1820_,
		_w1821_
	);
	LUT2 #(
		.INIT('h8)
	) name1580 (
		_w1277_,
		_w1788_,
		_w1822_
	);
	LUT4 #(
		.INIT('h0e0a)
	) name1581 (
		\shift_data_reg[21]/NET0131 ,
		_w1277_,
		_w1346_,
		_w1788_,
		_w1823_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1582 (
		_w1165_,
		_w1262_,
		_w1822_,
		_w1823_,
		_w1824_
	);
	LUT2 #(
		.INIT('he)
	) name1583 (
		_w1821_,
		_w1824_,
		_w1825_
	);
	LUT3 #(
		.INIT('h35)
	) name1584 (
		\shift_data_reg[22]/NET0131 ,
		\wb_dat_i[22]_pad ,
		\wb_sel_i[2]_pad ,
		_w1826_
	);
	LUT4 #(
		.INIT('h0040)
	) name1585 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1826_,
		_w1827_
	);
	LUT2 #(
		.INIT('h8)
	) name1586 (
		_w1297_,
		_w1788_,
		_w1828_
	);
	LUT4 #(
		.INIT('h0e0a)
	) name1587 (
		\shift_data_reg[22]/NET0131 ,
		_w1297_,
		_w1346_,
		_w1788_,
		_w1829_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1588 (
		_w1165_,
		_w1262_,
		_w1828_,
		_w1829_,
		_w1830_
	);
	LUT2 #(
		.INIT('he)
	) name1589 (
		_w1827_,
		_w1830_,
		_w1831_
	);
	LUT3 #(
		.INIT('h35)
	) name1590 (
		\shift_data_reg[23]/NET0131 ,
		\wb_dat_i[23]_pad ,
		\wb_sel_i[2]_pad ,
		_w1832_
	);
	LUT4 #(
		.INIT('h0040)
	) name1591 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1832_,
		_w1833_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name1592 (
		\shift_data_reg[23]/NET0131 ,
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1834_
	);
	LUT3 #(
		.INIT('h0b)
	) name1593 (
		_w1264_,
		_w1060_,
		_w1834_,
		_w1835_
	);
	LUT3 #(
		.INIT('h80)
	) name1594 (
		_w1033_,
		_w1065_,
		_w1351_,
		_w1836_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1595 (
		\shift_data_reg[23]/NET0131 ,
		_w1033_,
		_w1065_,
		_w1351_,
		_w1837_
	);
	LUT2 #(
		.INIT('h2)
	) name1596 (
		_w1614_,
		_w1837_,
		_w1838_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1597 (
		_w1165_,
		_w1262_,
		_w1836_,
		_w1838_,
		_w1839_
	);
	LUT3 #(
		.INIT('hab)
	) name1598 (
		_w1833_,
		_w1835_,
		_w1839_,
		_w1840_
	);
	LUT3 #(
		.INIT('h35)
	) name1599 (
		\shift_data_reg[24]/NET0131 ,
		\wb_dat_i[24]_pad ,
		\wb_sel_i[3]_pad ,
		_w1841_
	);
	LUT4 #(
		.INIT('h0040)
	) name1600 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1841_,
		_w1842_
	);
	LUT2 #(
		.INIT('h4)
	) name1601 (
		_w1032_,
		_w1306_,
		_w1843_
	);
	LUT4 #(
		.INIT('h8000)
	) name1602 (
		_w1065_,
		_w1351_,
		_w1614_,
		_w1843_,
		_w1844_
	);
	LUT3 #(
		.INIT('h32)
	) name1603 (
		\shift_data_reg[24]/NET0131 ,
		_w1346_,
		_w1844_,
		_w1845_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1604 (
		_w1165_,
		_w1262_,
		_w1844_,
		_w1845_,
		_w1846_
	);
	LUT2 #(
		.INIT('he)
	) name1605 (
		_w1842_,
		_w1846_,
		_w1847_
	);
	LUT3 #(
		.INIT('h80)
	) name1606 (
		_w1278_,
		_w1307_,
		_w1352_,
		_w1848_
	);
	LUT4 #(
		.INIT('h1555)
	) name1607 (
		\shift_data_reg[33]/NET0131 ,
		_w1278_,
		_w1307_,
		_w1352_,
		_w1849_
	);
	LUT2 #(
		.INIT('h1)
	) name1608 (
		_w1264_,
		_w1849_,
		_w1850_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1609 (
		_w1165_,
		_w1262_,
		_w1848_,
		_w1850_,
		_w1851_
	);
	LUT4 #(
		.INIT('h8000)
	) name1610 (
		\wb_adr_i[2]_pad ,
		_w858_,
		_w1055_,
		_w1263_,
		_w1852_
	);
	LUT4 #(
		.INIT('h0080)
	) name1611 (
		\shift_data_reg[33]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1313_,
		_w1853_
	);
	LUT2 #(
		.INIT('h1)
	) name1612 (
		_w1852_,
		_w1853_,
		_w1854_
	);
	LUT2 #(
		.INIT('hb)
	) name1613 (
		_w1851_,
		_w1854_,
		_w1855_
	);
	LUT3 #(
		.INIT('h80)
	) name1614 (
		_w1278_,
		_w1307_,
		_w1388_,
		_w1856_
	);
	LUT4 #(
		.INIT('h1555)
	) name1615 (
		\shift_data_reg[34]/NET0131 ,
		_w1278_,
		_w1307_,
		_w1388_,
		_w1857_
	);
	LUT2 #(
		.INIT('h1)
	) name1616 (
		_w1264_,
		_w1857_,
		_w1858_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1617 (
		_w1165_,
		_w1262_,
		_w1856_,
		_w1858_,
		_w1859_
	);
	LUT4 #(
		.INIT('h8000)
	) name1618 (
		\wb_adr_i[2]_pad ,
		_w833_,
		_w1055_,
		_w1263_,
		_w1860_
	);
	LUT4 #(
		.INIT('h0080)
	) name1619 (
		\shift_data_reg[34]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1313_,
		_w1861_
	);
	LUT2 #(
		.INIT('h1)
	) name1620 (
		_w1860_,
		_w1861_,
		_w1862_
	);
	LUT2 #(
		.INIT('hb)
	) name1621 (
		_w1859_,
		_w1862_,
		_w1863_
	);
	LUT3 #(
		.INIT('h80)
	) name1622 (
		_w1278_,
		_w1307_,
		_w1398_,
		_w1864_
	);
	LUT4 #(
		.INIT('h1555)
	) name1623 (
		\shift_data_reg[35]/NET0131 ,
		_w1278_,
		_w1307_,
		_w1398_,
		_w1865_
	);
	LUT2 #(
		.INIT('h1)
	) name1624 (
		_w1264_,
		_w1865_,
		_w1866_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1625 (
		_w1165_,
		_w1262_,
		_w1864_,
		_w1866_,
		_w1867_
	);
	LUT4 #(
		.INIT('h8000)
	) name1626 (
		\wb_adr_i[2]_pad ,
		_w868_,
		_w1055_,
		_w1263_,
		_w1868_
	);
	LUT4 #(
		.INIT('h0080)
	) name1627 (
		\shift_data_reg[35]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1313_,
		_w1869_
	);
	LUT2 #(
		.INIT('h1)
	) name1628 (
		_w1868_,
		_w1869_,
		_w1870_
	);
	LUT2 #(
		.INIT('hb)
	) name1629 (
		_w1867_,
		_w1870_,
		_w1871_
	);
	LUT3 #(
		.INIT('h80)
	) name1630 (
		_w1278_,
		_w1307_,
		_w1361_,
		_w1872_
	);
	LUT4 #(
		.INIT('h1555)
	) name1631 (
		\shift_data_reg[36]/NET0131 ,
		_w1278_,
		_w1307_,
		_w1361_,
		_w1873_
	);
	LUT2 #(
		.INIT('h1)
	) name1632 (
		_w1264_,
		_w1873_,
		_w1874_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1633 (
		_w1165_,
		_w1262_,
		_w1872_,
		_w1874_,
		_w1875_
	);
	LUT4 #(
		.INIT('h8000)
	) name1634 (
		\wb_adr_i[2]_pad ,
		_w806_,
		_w1055_,
		_w1263_,
		_w1876_
	);
	LUT4 #(
		.INIT('h0080)
	) name1635 (
		\shift_data_reg[36]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1313_,
		_w1877_
	);
	LUT2 #(
		.INIT('h1)
	) name1636 (
		_w1876_,
		_w1877_,
		_w1878_
	);
	LUT2 #(
		.INIT('hb)
	) name1637 (
		_w1875_,
		_w1878_,
		_w1879_
	);
	LUT3 #(
		.INIT('h80)
	) name1638 (
		_w1277_,
		_w1278_,
		_w1307_,
		_w1880_
	);
	LUT4 #(
		.INIT('h1555)
	) name1639 (
		\shift_data_reg[37]/NET0131 ,
		_w1277_,
		_w1278_,
		_w1307_,
		_w1881_
	);
	LUT2 #(
		.INIT('h1)
	) name1640 (
		_w1264_,
		_w1881_,
		_w1882_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1641 (
		_w1165_,
		_w1262_,
		_w1880_,
		_w1882_,
		_w1883_
	);
	LUT4 #(
		.INIT('h8000)
	) name1642 (
		\wb_adr_i[2]_pad ,
		_w826_,
		_w1055_,
		_w1263_,
		_w1884_
	);
	LUT4 #(
		.INIT('h0080)
	) name1643 (
		\shift_data_reg[37]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1313_,
		_w1885_
	);
	LUT2 #(
		.INIT('h1)
	) name1644 (
		_w1884_,
		_w1885_,
		_w1886_
	);
	LUT2 #(
		.INIT('hb)
	) name1645 (
		_w1883_,
		_w1886_,
		_w1887_
	);
	LUT3 #(
		.INIT('h80)
	) name1646 (
		_w1278_,
		_w1297_,
		_w1307_,
		_w1888_
	);
	LUT4 #(
		.INIT('h1555)
	) name1647 (
		\shift_data_reg[38]/NET0131 ,
		_w1278_,
		_w1297_,
		_w1307_,
		_w1889_
	);
	LUT2 #(
		.INIT('h1)
	) name1648 (
		_w1264_,
		_w1889_,
		_w1890_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1649 (
		_w1165_,
		_w1262_,
		_w1888_,
		_w1890_,
		_w1891_
	);
	LUT4 #(
		.INIT('h8000)
	) name1650 (
		\wb_adr_i[2]_pad ,
		_w848_,
		_w1055_,
		_w1263_,
		_w1892_
	);
	LUT4 #(
		.INIT('h0080)
	) name1651 (
		\shift_data_reg[38]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1313_,
		_w1893_
	);
	LUT2 #(
		.INIT('h1)
	) name1652 (
		_w1892_,
		_w1893_,
		_w1894_
	);
	LUT2 #(
		.INIT('hb)
	) name1653 (
		_w1891_,
		_w1894_,
		_w1895_
	);
	LUT3 #(
		.INIT('h80)
	) name1654 (
		_w1278_,
		_w1306_,
		_w1325_,
		_w1896_
	);
	LUT4 #(
		.INIT('h1555)
	) name1655 (
		\shift_data_reg[40]/NET0131 ,
		_w1278_,
		_w1306_,
		_w1325_,
		_w1897_
	);
	LUT2 #(
		.INIT('h1)
	) name1656 (
		_w1264_,
		_w1897_,
		_w1898_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1657 (
		_w1165_,
		_w1262_,
		_w1896_,
		_w1898_,
		_w1899_
	);
	LUT4 #(
		.INIT('h8000)
	) name1658 (
		\wb_adr_i[2]_pad ,
		_w583_,
		_w1055_,
		_w1263_,
		_w1900_
	);
	LUT2 #(
		.INIT('h8)
	) name1659 (
		\wb_adr_i[2]_pad ,
		\wb_sel_i[1]_pad ,
		_w1901_
	);
	LUT4 #(
		.INIT('h0080)
	) name1660 (
		\shift_data_reg[40]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1901_,
		_w1902_
	);
	LUT2 #(
		.INIT('h1)
	) name1661 (
		_w1900_,
		_w1902_,
		_w1903_
	);
	LUT2 #(
		.INIT('hb)
	) name1662 (
		_w1899_,
		_w1903_,
		_w1904_
	);
	LUT3 #(
		.INIT('h80)
	) name1663 (
		_w1278_,
		_w1325_,
		_w1352_,
		_w1905_
	);
	LUT4 #(
		.INIT('h1555)
	) name1664 (
		\shift_data_reg[41]/NET0131 ,
		_w1278_,
		_w1325_,
		_w1352_,
		_w1906_
	);
	LUT2 #(
		.INIT('h1)
	) name1665 (
		_w1264_,
		_w1906_,
		_w1907_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1666 (
		_w1165_,
		_w1262_,
		_w1905_,
		_w1907_,
		_w1908_
	);
	LUT4 #(
		.INIT('h8000)
	) name1667 (
		\wb_adr_i[2]_pad ,
		_w885_,
		_w1055_,
		_w1263_,
		_w1909_
	);
	LUT4 #(
		.INIT('h0080)
	) name1668 (
		\shift_data_reg[41]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1901_,
		_w1910_
	);
	LUT2 #(
		.INIT('h1)
	) name1669 (
		_w1909_,
		_w1910_,
		_w1911_
	);
	LUT2 #(
		.INIT('hb)
	) name1670 (
		_w1908_,
		_w1911_,
		_w1912_
	);
	LUT3 #(
		.INIT('h80)
	) name1671 (
		_w1278_,
		_w1325_,
		_w1388_,
		_w1913_
	);
	LUT4 #(
		.INIT('h1555)
	) name1672 (
		\shift_data_reg[42]/NET0131 ,
		_w1278_,
		_w1325_,
		_w1388_,
		_w1914_
	);
	LUT2 #(
		.INIT('h1)
	) name1673 (
		_w1264_,
		_w1914_,
		_w1915_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1674 (
		_w1165_,
		_w1262_,
		_w1913_,
		_w1915_,
		_w1916_
	);
	LUT4 #(
		.INIT('h8000)
	) name1675 (
		\wb_adr_i[2]_pad ,
		_w814_,
		_w1055_,
		_w1263_,
		_w1917_
	);
	LUT4 #(
		.INIT('h0080)
	) name1676 (
		\shift_data_reg[42]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1901_,
		_w1918_
	);
	LUT2 #(
		.INIT('h1)
	) name1677 (
		_w1917_,
		_w1918_,
		_w1919_
	);
	LUT2 #(
		.INIT('hb)
	) name1678 (
		_w1916_,
		_w1919_,
		_w1920_
	);
	LUT3 #(
		.INIT('h80)
	) name1679 (
		_w1278_,
		_w1325_,
		_w1398_,
		_w1921_
	);
	LUT4 #(
		.INIT('h1555)
	) name1680 (
		\shift_data_reg[43]/NET0131 ,
		_w1278_,
		_w1325_,
		_w1398_,
		_w1922_
	);
	LUT2 #(
		.INIT('h1)
	) name1681 (
		_w1264_,
		_w1922_,
		_w1923_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1682 (
		_w1165_,
		_w1262_,
		_w1921_,
		_w1923_,
		_w1924_
	);
	LUT4 #(
		.INIT('h8000)
	) name1683 (
		\wb_adr_i[2]_pad ,
		_w840_,
		_w1055_,
		_w1263_,
		_w1925_
	);
	LUT4 #(
		.INIT('h0080)
	) name1684 (
		\shift_data_reg[43]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1901_,
		_w1926_
	);
	LUT2 #(
		.INIT('h1)
	) name1685 (
		_w1925_,
		_w1926_,
		_w1927_
	);
	LUT2 #(
		.INIT('hb)
	) name1686 (
		_w1924_,
		_w1927_,
		_w1928_
	);
	LUT3 #(
		.INIT('h80)
	) name1687 (
		_w1278_,
		_w1325_,
		_w1361_,
		_w1929_
	);
	LUT4 #(
		.INIT('h1555)
	) name1688 (
		\shift_data_reg[44]/NET0131 ,
		_w1278_,
		_w1325_,
		_w1361_,
		_w1930_
	);
	LUT2 #(
		.INIT('h1)
	) name1689 (
		_w1264_,
		_w1930_,
		_w1931_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1690 (
		_w1165_,
		_w1262_,
		_w1929_,
		_w1931_,
		_w1932_
	);
	LUT4 #(
		.INIT('h8000)
	) name1691 (
		\wb_adr_i[2]_pad ,
		_w878_,
		_w1055_,
		_w1263_,
		_w1933_
	);
	LUT4 #(
		.INIT('h0080)
	) name1692 (
		\shift_data_reg[44]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1901_,
		_w1934_
	);
	LUT2 #(
		.INIT('h1)
	) name1693 (
		_w1933_,
		_w1934_,
		_w1935_
	);
	LUT2 #(
		.INIT('hb)
	) name1694 (
		_w1932_,
		_w1935_,
		_w1936_
	);
	LUT3 #(
		.INIT('h80)
	) name1695 (
		_w1277_,
		_w1278_,
		_w1325_,
		_w1937_
	);
	LUT4 #(
		.INIT('h1555)
	) name1696 (
		\shift_data_reg[45]/NET0131 ,
		_w1277_,
		_w1278_,
		_w1325_,
		_w1938_
	);
	LUT2 #(
		.INIT('h1)
	) name1697 (
		_w1264_,
		_w1938_,
		_w1939_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1698 (
		_w1165_,
		_w1262_,
		_w1937_,
		_w1939_,
		_w1940_
	);
	LUT4 #(
		.INIT('h8000)
	) name1699 (
		\wb_adr_i[2]_pad ,
		_w822_,
		_w1055_,
		_w1263_,
		_w1941_
	);
	LUT4 #(
		.INIT('h0080)
	) name1700 (
		\shift_data_reg[45]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1901_,
		_w1942_
	);
	LUT2 #(
		.INIT('h1)
	) name1701 (
		_w1941_,
		_w1942_,
		_w1943_
	);
	LUT2 #(
		.INIT('hb)
	) name1702 (
		_w1940_,
		_w1943_,
		_w1944_
	);
	LUT3 #(
		.INIT('h80)
	) name1703 (
		_w1278_,
		_w1297_,
		_w1325_,
		_w1945_
	);
	LUT4 #(
		.INIT('h1555)
	) name1704 (
		\shift_data_reg[46]/NET0131 ,
		_w1278_,
		_w1297_,
		_w1325_,
		_w1946_
	);
	LUT2 #(
		.INIT('h1)
	) name1705 (
		_w1264_,
		_w1946_,
		_w1947_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1706 (
		_w1165_,
		_w1262_,
		_w1945_,
		_w1947_,
		_w1948_
	);
	LUT4 #(
		.INIT('h8000)
	) name1707 (
		\wb_adr_i[2]_pad ,
		_w844_,
		_w1055_,
		_w1263_,
		_w1949_
	);
	LUT4 #(
		.INIT('h0080)
	) name1708 (
		\shift_data_reg[46]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1901_,
		_w1950_
	);
	LUT2 #(
		.INIT('h1)
	) name1709 (
		_w1949_,
		_w1950_,
		_w1951_
	);
	LUT2 #(
		.INIT('hb)
	) name1710 (
		_w1948_,
		_w1951_,
		_w1952_
	);
	LUT3 #(
		.INIT('h80)
	) name1711 (
		_w1025_,
		_w1278_,
		_w1325_,
		_w1953_
	);
	LUT4 #(
		.INIT('h1555)
	) name1712 (
		\shift_data_reg[47]/NET0131 ,
		_w1025_,
		_w1278_,
		_w1325_,
		_w1954_
	);
	LUT2 #(
		.INIT('h1)
	) name1713 (
		_w1264_,
		_w1954_,
		_w1955_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1714 (
		_w1165_,
		_w1262_,
		_w1953_,
		_w1955_,
		_w1956_
	);
	LUT4 #(
		.INIT('h8000)
	) name1715 (
		\wb_adr_i[2]_pad ,
		_w899_,
		_w1055_,
		_w1263_,
		_w1957_
	);
	LUT4 #(
		.INIT('h0080)
	) name1716 (
		\shift_data_reg[47]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1901_,
		_w1958_
	);
	LUT2 #(
		.INIT('h1)
	) name1717 (
		_w1957_,
		_w1958_,
		_w1959_
	);
	LUT2 #(
		.INIT('hb)
	) name1718 (
		_w1956_,
		_w1959_,
		_w1960_
	);
	LUT3 #(
		.INIT('h80)
	) name1719 (
		_w1054_,
		_w1066_,
		_w1369_,
		_w1961_
	);
	LUT4 #(
		.INIT('h1555)
	) name1720 (
		\shift_data_reg[48]/NET0131 ,
		_w1054_,
		_w1066_,
		_w1369_,
		_w1962_
	);
	LUT2 #(
		.INIT('h1)
	) name1721 (
		_w1264_,
		_w1962_,
		_w1963_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1722 (
		_w1165_,
		_w1262_,
		_w1961_,
		_w1963_,
		_w1964_
	);
	LUT4 #(
		.INIT('h8000)
	) name1723 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1516_,
		_w1965_
	);
	LUT4 #(
		.INIT('h0080)
	) name1724 (
		\shift_data_reg[48]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1271_,
		_w1966_
	);
	LUT2 #(
		.INIT('h1)
	) name1725 (
		_w1965_,
		_w1966_,
		_w1967_
	);
	LUT2 #(
		.INIT('hb)
	) name1726 (
		_w1964_,
		_w1967_,
		_w1968_
	);
	LUT3 #(
		.INIT('h80)
	) name1727 (
		_w1054_,
		_w1066_,
		_w1379_,
		_w1969_
	);
	LUT4 #(
		.INIT('h1555)
	) name1728 (
		\shift_data_reg[49]/NET0131 ,
		_w1054_,
		_w1066_,
		_w1379_,
		_w1970_
	);
	LUT2 #(
		.INIT('h1)
	) name1729 (
		_w1264_,
		_w1970_,
		_w1971_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1730 (
		_w1165_,
		_w1262_,
		_w1969_,
		_w1971_,
		_w1972_
	);
	LUT4 #(
		.INIT('h8000)
	) name1731 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1498_,
		_w1973_
	);
	LUT4 #(
		.INIT('h0080)
	) name1732 (
		\shift_data_reg[49]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1271_,
		_w1974_
	);
	LUT2 #(
		.INIT('h1)
	) name1733 (
		_w1973_,
		_w1974_,
		_w1975_
	);
	LUT2 #(
		.INIT('hb)
	) name1734 (
		_w1972_,
		_w1975_,
		_w1976_
	);
	LUT3 #(
		.INIT('h80)
	) name1735 (
		_w1054_,
		_w1066_,
		_w1389_,
		_w1977_
	);
	LUT4 #(
		.INIT('h1555)
	) name1736 (
		\shift_data_reg[50]/NET0131 ,
		_w1054_,
		_w1066_,
		_w1389_,
		_w1978_
	);
	LUT2 #(
		.INIT('h1)
	) name1737 (
		_w1264_,
		_w1978_,
		_w1979_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1738 (
		_w1165_,
		_w1262_,
		_w1977_,
		_w1979_,
		_w1980_
	);
	LUT4 #(
		.INIT('h8000)
	) name1739 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1508_,
		_w1981_
	);
	LUT4 #(
		.INIT('h0080)
	) name1740 (
		\shift_data_reg[50]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1271_,
		_w1982_
	);
	LUT2 #(
		.INIT('h1)
	) name1741 (
		_w1981_,
		_w1982_,
		_w1983_
	);
	LUT2 #(
		.INIT('hb)
	) name1742 (
		_w1980_,
		_w1983_,
		_w1984_
	);
	LUT4 #(
		.INIT('ha800)
	) name1743 (
		_w1042_,
		_w1049_,
		_w1052_,
		_w1398_,
		_w1985_
	);
	LUT2 #(
		.INIT('h8)
	) name1744 (
		_w1307_,
		_w1985_,
		_w1986_
	);
	LUT4 #(
		.INIT('h3222)
	) name1745 (
		\shift_data_reg[51]/NET0131 ,
		_w1264_,
		_w1307_,
		_w1985_,
		_w1987_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1746 (
		_w1165_,
		_w1262_,
		_w1986_,
		_w1987_,
		_w1988_
	);
	LUT4 #(
		.INIT('h8000)
	) name1747 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1524_,
		_w1989_
	);
	LUT4 #(
		.INIT('h0080)
	) name1748 (
		\shift_data_reg[51]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1271_,
		_w1990_
	);
	LUT2 #(
		.INIT('h1)
	) name1749 (
		_w1989_,
		_w1990_,
		_w1991_
	);
	LUT2 #(
		.INIT('hb)
	) name1750 (
		_w1988_,
		_w1991_,
		_w1992_
	);
	LUT3 #(
		.INIT('h80)
	) name1751 (
		_w1054_,
		_w1066_,
		_w1406_,
		_w1993_
	);
	LUT4 #(
		.INIT('h1555)
	) name1752 (
		\shift_data_reg[52]/NET0131 ,
		_w1054_,
		_w1066_,
		_w1406_,
		_w1994_
	);
	LUT2 #(
		.INIT('h1)
	) name1753 (
		_w1264_,
		_w1994_,
		_w1995_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1754 (
		_w1165_,
		_w1262_,
		_w1993_,
		_w1995_,
		_w1996_
	);
	LUT4 #(
		.INIT('h8000)
	) name1755 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1532_,
		_w1997_
	);
	LUT4 #(
		.INIT('h0080)
	) name1756 (
		\shift_data_reg[52]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1271_,
		_w1998_
	);
	LUT2 #(
		.INIT('h1)
	) name1757 (
		_w1997_,
		_w1998_,
		_w1999_
	);
	LUT2 #(
		.INIT('hb)
	) name1758 (
		_w1996_,
		_w1999_,
		_w2000_
	);
	LUT4 #(
		.INIT('ha800)
	) name1759 (
		_w1042_,
		_w1049_,
		_w1052_,
		_w1277_,
		_w2001_
	);
	LUT2 #(
		.INIT('h8)
	) name1760 (
		_w1307_,
		_w2001_,
		_w2002_
	);
	LUT4 #(
		.INIT('h3222)
	) name1761 (
		\shift_data_reg[53]/NET0131 ,
		_w1264_,
		_w1307_,
		_w2001_,
		_w2003_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1762 (
		_w1165_,
		_w1262_,
		_w2002_,
		_w2003_,
		_w2004_
	);
	LUT4 #(
		.INIT('h8000)
	) name1763 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1541_,
		_w2005_
	);
	LUT4 #(
		.INIT('h0080)
	) name1764 (
		\shift_data_reg[53]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1271_,
		_w2006_
	);
	LUT2 #(
		.INIT('h1)
	) name1765 (
		_w2005_,
		_w2006_,
		_w2007_
	);
	LUT2 #(
		.INIT('hb)
	) name1766 (
		_w2004_,
		_w2007_,
		_w2008_
	);
	LUT4 #(
		.INIT('ha800)
	) name1767 (
		_w1042_,
		_w1049_,
		_w1052_,
		_w1297_,
		_w2009_
	);
	LUT2 #(
		.INIT('h8)
	) name1768 (
		_w1307_,
		_w2009_,
		_w2010_
	);
	LUT4 #(
		.INIT('h3222)
	) name1769 (
		\shift_data_reg[54]/NET0131 ,
		_w1264_,
		_w1307_,
		_w2009_,
		_w2011_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1770 (
		_w1165_,
		_w1262_,
		_w2010_,
		_w2011_,
		_w2012_
	);
	LUT4 #(
		.INIT('h8000)
	) name1771 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1549_,
		_w2013_
	);
	LUT4 #(
		.INIT('h0080)
	) name1772 (
		\shift_data_reg[54]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1271_,
		_w2014_
	);
	LUT2 #(
		.INIT('h1)
	) name1773 (
		_w2013_,
		_w2014_,
		_w2015_
	);
	LUT2 #(
		.INIT('hb)
	) name1774 (
		_w2012_,
		_w2015_,
		_w2016_
	);
	LUT3 #(
		.INIT('h80)
	) name1775 (
		_w1054_,
		_w1325_,
		_w1352_,
		_w2017_
	);
	LUT4 #(
		.INIT('h1555)
	) name1776 (
		\shift_data_reg[57]/NET0131 ,
		_w1054_,
		_w1325_,
		_w1352_,
		_w2018_
	);
	LUT2 #(
		.INIT('h1)
	) name1777 (
		_w1264_,
		_w2018_,
		_w2019_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1778 (
		_w1165_,
		_w1262_,
		_w2017_,
		_w2019_,
		_w2020_
	);
	LUT4 #(
		.INIT('h8000)
	) name1779 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1347_,
		_w2021_
	);
	LUT4 #(
		.INIT('h0080)
	) name1780 (
		\shift_data_reg[57]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1332_,
		_w2022_
	);
	LUT2 #(
		.INIT('h1)
	) name1781 (
		_w2021_,
		_w2022_,
		_w2023_
	);
	LUT2 #(
		.INIT('hb)
	) name1782 (
		_w2020_,
		_w2023_,
		_w2024_
	);
	LUT3 #(
		.INIT('h80)
	) name1783 (
		_w1054_,
		_w1325_,
		_w1388_,
		_w2025_
	);
	LUT4 #(
		.INIT('h1555)
	) name1784 (
		\shift_data_reg[58]/NET0131 ,
		_w1054_,
		_w1325_,
		_w1388_,
		_w2026_
	);
	LUT2 #(
		.INIT('h1)
	) name1785 (
		_w1264_,
		_w2026_,
		_w2027_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1786 (
		_w1165_,
		_w1262_,
		_w2025_,
		_w2027_,
		_w2028_
	);
	LUT4 #(
		.INIT('h8000)
	) name1787 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1572_,
		_w2029_
	);
	LUT4 #(
		.INIT('h0080)
	) name1788 (
		\shift_data_reg[58]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1332_,
		_w2030_
	);
	LUT2 #(
		.INIT('h1)
	) name1789 (
		_w2029_,
		_w2030_,
		_w2031_
	);
	LUT2 #(
		.INIT('hb)
	) name1790 (
		_w2028_,
		_w2031_,
		_w2032_
	);
	LUT2 #(
		.INIT('h8)
	) name1791 (
		_w1325_,
		_w1985_,
		_w2033_
	);
	LUT4 #(
		.INIT('h3222)
	) name1792 (
		\shift_data_reg[59]/NET0131 ,
		_w1264_,
		_w1325_,
		_w1985_,
		_w2034_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1793 (
		_w1165_,
		_w1262_,
		_w2033_,
		_w2034_,
		_w2035_
	);
	LUT4 #(
		.INIT('h8000)
	) name1794 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1580_,
		_w2036_
	);
	LUT4 #(
		.INIT('h0080)
	) name1795 (
		\shift_data_reg[59]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1332_,
		_w2037_
	);
	LUT2 #(
		.INIT('h1)
	) name1796 (
		_w2036_,
		_w2037_,
		_w2038_
	);
	LUT2 #(
		.INIT('hb)
	) name1797 (
		_w2035_,
		_w2038_,
		_w2039_
	);
	LUT3 #(
		.INIT('h80)
	) name1798 (
		_w1054_,
		_w1325_,
		_w1361_,
		_w2040_
	);
	LUT4 #(
		.INIT('h1555)
	) name1799 (
		\shift_data_reg[60]/NET0131 ,
		_w1054_,
		_w1325_,
		_w1361_,
		_w2041_
	);
	LUT2 #(
		.INIT('h1)
	) name1800 (
		_w1264_,
		_w2041_,
		_w2042_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1801 (
		_w1165_,
		_w1262_,
		_w2040_,
		_w2042_,
		_w2043_
	);
	LUT4 #(
		.INIT('h8000)
	) name1802 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1358_,
		_w2044_
	);
	LUT4 #(
		.INIT('h0080)
	) name1803 (
		\shift_data_reg[60]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1332_,
		_w2045_
	);
	LUT2 #(
		.INIT('h1)
	) name1804 (
		_w2044_,
		_w2045_,
		_w2046_
	);
	LUT2 #(
		.INIT('hb)
	) name1805 (
		_w2043_,
		_w2046_,
		_w2047_
	);
	LUT2 #(
		.INIT('h8)
	) name1806 (
		_w1325_,
		_w2001_,
		_w2048_
	);
	LUT4 #(
		.INIT('h3222)
	) name1807 (
		\shift_data_reg[61]/NET0131 ,
		_w1264_,
		_w1325_,
		_w2001_,
		_w2049_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1808 (
		_w1165_,
		_w1262_,
		_w2048_,
		_w2049_,
		_w2050_
	);
	LUT4 #(
		.INIT('h8000)
	) name1809 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1588_,
		_w2051_
	);
	LUT4 #(
		.INIT('h0080)
	) name1810 (
		\shift_data_reg[61]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1332_,
		_w2052_
	);
	LUT2 #(
		.INIT('h1)
	) name1811 (
		_w2051_,
		_w2052_,
		_w2053_
	);
	LUT2 #(
		.INIT('hb)
	) name1812 (
		_w2050_,
		_w2053_,
		_w2054_
	);
	LUT2 #(
		.INIT('h8)
	) name1813 (
		_w1325_,
		_w2009_,
		_w2055_
	);
	LUT4 #(
		.INIT('h3222)
	) name1814 (
		\shift_data_reg[62]/NET0131 ,
		_w1264_,
		_w1325_,
		_w2009_,
		_w2056_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1815 (
		_w1165_,
		_w1262_,
		_w2055_,
		_w2056_,
		_w2057_
	);
	LUT4 #(
		.INIT('h8000)
	) name1816 (
		\wb_adr_i[2]_pad ,
		_w1055_,
		_w1263_,
		_w1596_,
		_w2058_
	);
	LUT4 #(
		.INIT('h0080)
	) name1817 (
		\shift_data_reg[62]/NET0131 ,
		_w1055_,
		_w1263_,
		_w1332_,
		_w2059_
	);
	LUT2 #(
		.INIT('h1)
	) name1818 (
		_w2058_,
		_w2059_,
		_w2060_
	);
	LUT2 #(
		.INIT('hb)
	) name1819 (
		_w2057_,
		_w2060_,
		_w2061_
	);
	LUT3 #(
		.INIT('h35)
	) name1820 (
		\shift_data_reg[105]/NET0131 ,
		\wb_dat_i[9]_pad ,
		\wb_sel_i[1]_pad ,
		_w2062_
	);
	LUT3 #(
		.INIT('h08)
	) name1821 (
		_w804_,
		_w1057_,
		_w2062_,
		_w2063_
	);
	LUT4 #(
		.INIT('h1000)
	) name1822 (
		_w1032_,
		_w1065_,
		_w1278_,
		_w1352_,
		_w2064_
	);
	LUT3 #(
		.INIT('hc8)
	) name1823 (
		\shift_data_reg[105]/NET0131 ,
		_w1060_,
		_w2064_,
		_w2065_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1824 (
		_w1165_,
		_w1262_,
		_w2064_,
		_w2065_,
		_w2066_
	);
	LUT2 #(
		.INIT('h2)
	) name1825 (
		\shift_data_reg[105]/NET0131 ,
		_w1283_,
		_w2067_
	);
	LUT4 #(
		.INIT('hff54)
	) name1826 (
		_w1264_,
		_w2063_,
		_w2066_,
		_w2067_,
		_w2068_
	);
	LUT3 #(
		.INIT('h35)
	) name1827 (
		\shift_data_reg[113]/NET0131 ,
		\wb_dat_i[17]_pad ,
		\wb_sel_i[2]_pad ,
		_w2069_
	);
	LUT3 #(
		.INIT('h08)
	) name1828 (
		_w804_,
		_w1057_,
		_w2069_,
		_w2070_
	);
	LUT3 #(
		.INIT('h20)
	) name1829 (
		_w1054_,
		_w1065_,
		_w1379_,
		_w2071_
	);
	LUT4 #(
		.INIT('h5155)
	) name1830 (
		\shift_data_reg[113]/NET0131 ,
		_w1054_,
		_w1065_,
		_w1379_,
		_w2072_
	);
	LUT2 #(
		.INIT('h2)
	) name1831 (
		_w1060_,
		_w2072_,
		_w2073_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1832 (
		_w1165_,
		_w1262_,
		_w2071_,
		_w2073_,
		_w2074_
	);
	LUT2 #(
		.INIT('h2)
	) name1833 (
		\shift_data_reg[113]/NET0131 ,
		_w1283_,
		_w2075_
	);
	LUT4 #(
		.INIT('hff54)
	) name1834 (
		_w1264_,
		_w2070_,
		_w2074_,
		_w2075_,
		_w2076_
	);
	LUT3 #(
		.INIT('h35)
	) name1835 (
		\shift_data_reg[108]/NET0131 ,
		\wb_dat_i[12]_pad ,
		\wb_sel_i[1]_pad ,
		_w2077_
	);
	LUT3 #(
		.INIT('h08)
	) name1836 (
		_w804_,
		_w1057_,
		_w2077_,
		_w2078_
	);
	LUT4 #(
		.INIT('h1000)
	) name1837 (
		_w1032_,
		_w1065_,
		_w1278_,
		_w1361_,
		_w2079_
	);
	LUT3 #(
		.INIT('hc8)
	) name1838 (
		\shift_data_reg[108]/NET0131 ,
		_w1060_,
		_w2079_,
		_w2080_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1839 (
		_w1165_,
		_w1262_,
		_w2079_,
		_w2080_,
		_w2081_
	);
	LUT2 #(
		.INIT('h2)
	) name1840 (
		\shift_data_reg[108]/NET0131 ,
		_w1283_,
		_w2082_
	);
	LUT4 #(
		.INIT('hff54)
	) name1841 (
		_w1264_,
		_w2078_,
		_w2081_,
		_w2082_,
		_w2083_
	);
	LUT3 #(
		.INIT('h35)
	) name1842 (
		\shift_data_reg[116]/NET0131 ,
		\wb_dat_i[20]_pad ,
		\wb_sel_i[2]_pad ,
		_w2084_
	);
	LUT3 #(
		.INIT('h08)
	) name1843 (
		_w804_,
		_w1057_,
		_w2084_,
		_w2085_
	);
	LUT3 #(
		.INIT('h20)
	) name1844 (
		_w1054_,
		_w1065_,
		_w1406_,
		_w2086_
	);
	LUT4 #(
		.INIT('h5155)
	) name1845 (
		\shift_data_reg[116]/NET0131 ,
		_w1054_,
		_w1065_,
		_w1406_,
		_w2087_
	);
	LUT2 #(
		.INIT('h2)
	) name1846 (
		_w1060_,
		_w2087_,
		_w2088_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1847 (
		_w1165_,
		_w1262_,
		_w2086_,
		_w2088_,
		_w2089_
	);
	LUT2 #(
		.INIT('h2)
	) name1848 (
		\shift_data_reg[116]/NET0131 ,
		_w1283_,
		_w2090_
	);
	LUT4 #(
		.INIT('hff54)
	) name1849 (
		_w1264_,
		_w2085_,
		_w2089_,
		_w2090_,
		_w2091_
	);
	LUT3 #(
		.INIT('h20)
	) name1850 (
		_w1054_,
		_w1065_,
		_w1843_,
		_w2092_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1851 (
		_w1060_,
		_w1165_,
		_w1262_,
		_w2092_,
		_w2093_
	);
	LUT3 #(
		.INIT('h35)
	) name1852 (
		\shift_data_reg[120]/NET0131 ,
		\wb_dat_i[24]_pad ,
		\wb_sel_i[3]_pad ,
		_w2094_
	);
	LUT3 #(
		.INIT('h08)
	) name1853 (
		_w804_,
		_w1057_,
		_w2094_,
		_w2095_
	);
	LUT4 #(
		.INIT('h02aa)
	) name1854 (
		\shift_data_reg[120]/NET0131 ,
		_w585_,
		_w804_,
		_w1057_,
		_w2096_
	);
	LUT4 #(
		.INIT('hdf00)
	) name1855 (
		_w1054_,
		_w1065_,
		_w1843_,
		_w2096_,
		_w2097_
	);
	LUT2 #(
		.INIT('h1)
	) name1856 (
		_w2095_,
		_w2097_,
		_w2098_
	);
	LUT2 #(
		.INIT('h2)
	) name1857 (
		\shift_data_reg[120]/NET0131 ,
		_w1283_,
		_w2099_
	);
	LUT4 #(
		.INIT('hff45)
	) name1858 (
		_w1264_,
		_w2093_,
		_w2098_,
		_w2099_,
		_w2100_
	);
	LUT3 #(
		.INIT('h80)
	) name1859 (
		_w804_,
		_w848_,
		_w1057_,
		_w2101_
	);
	LUT3 #(
		.INIT('h80)
	) name1860 (
		_w1278_,
		_w1279_,
		_w1297_,
		_w2102_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1861 (
		_w1060_,
		_w1165_,
		_w1262_,
		_w2102_,
		_w2103_
	);
	LUT4 #(
		.INIT('h1555)
	) name1862 (
		_w1059_,
		_w1278_,
		_w1279_,
		_w1297_,
		_w2104_
	);
	LUT3 #(
		.INIT('ha2)
	) name1863 (
		\shift_data_reg[102]/NET0131 ,
		_w1285_,
		_w2104_,
		_w2105_
	);
	LUT4 #(
		.INIT('hff54)
	) name1864 (
		_w1264_,
		_w2101_,
		_w2103_,
		_w2105_,
		_w2106_
	);
	LUT3 #(
		.INIT('h35)
	) name1865 (
		\shift_data_reg[107]/NET0131 ,
		\wb_dat_i[11]_pad ,
		\wb_sel_i[1]_pad ,
		_w2107_
	);
	LUT3 #(
		.INIT('h08)
	) name1866 (
		_w804_,
		_w1057_,
		_w2107_,
		_w2108_
	);
	LUT4 #(
		.INIT('h1000)
	) name1867 (
		_w1032_,
		_w1065_,
		_w1278_,
		_w1398_,
		_w2109_
	);
	LUT3 #(
		.INIT('hc8)
	) name1868 (
		\shift_data_reg[107]/NET0131 ,
		_w1060_,
		_w2109_,
		_w2110_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1869 (
		_w1165_,
		_w1262_,
		_w2109_,
		_w2110_,
		_w2111_
	);
	LUT2 #(
		.INIT('h2)
	) name1870 (
		\shift_data_reg[107]/NET0131 ,
		_w1283_,
		_w2112_
	);
	LUT4 #(
		.INIT('hff54)
	) name1871 (
		_w1264_,
		_w2108_,
		_w2111_,
		_w2112_,
		_w2113_
	);
	LUT2 #(
		.INIT('h2)
	) name1872 (
		\shift_data_reg[115]/NET0131 ,
		_w1283_,
		_w2114_
	);
	LUT2 #(
		.INIT('h8)
	) name1873 (
		_w1279_,
		_w1985_,
		_w2115_
	);
	LUT3 #(
		.INIT('h35)
	) name1874 (
		\shift_data_reg[115]/NET0131 ,
		\wb_dat_i[19]_pad ,
		\wb_sel_i[2]_pad ,
		_w2116_
	);
	LUT3 #(
		.INIT('h08)
	) name1875 (
		_w804_,
		_w1057_,
		_w2116_,
		_w2117_
	);
	LUT4 #(
		.INIT('h00d5)
	) name1876 (
		\shift_data_reg[115]/NET0131 ,
		_w1279_,
		_w1985_,
		_w2117_,
		_w2118_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1877 (
		_w1165_,
		_w1262_,
		_w2115_,
		_w2118_,
		_w2119_
	);
	LUT4 #(
		.INIT('he020)
	) name1878 (
		_w585_,
		_w804_,
		_w1057_,
		_w2116_,
		_w2120_
	);
	LUT2 #(
		.INIT('h1)
	) name1879 (
		_w1264_,
		_w2120_,
		_w2121_
	);
	LUT3 #(
		.INIT('hba)
	) name1880 (
		_w2114_,
		_w2119_,
		_w2121_,
		_w2122_
	);
	LUT3 #(
		.INIT('h35)
	) name1881 (
		\shift_data_reg[118]/NET0131 ,
		\wb_dat_i[22]_pad ,
		\wb_sel_i[2]_pad ,
		_w2123_
	);
	LUT3 #(
		.INIT('h08)
	) name1882 (
		_w804_,
		_w1057_,
		_w2123_,
		_w2124_
	);
	LUT2 #(
		.INIT('h8)
	) name1883 (
		_w1279_,
		_w2009_,
		_w2125_
	);
	LUT4 #(
		.INIT('hc888)
	) name1884 (
		\shift_data_reg[118]/NET0131 ,
		_w1060_,
		_w1279_,
		_w2009_,
		_w2126_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1885 (
		_w1165_,
		_w1262_,
		_w2125_,
		_w2126_,
		_w2127_
	);
	LUT2 #(
		.INIT('h2)
	) name1886 (
		\shift_data_reg[118]/NET0131 ,
		_w1283_,
		_w2128_
	);
	LUT4 #(
		.INIT('hff54)
	) name1887 (
		_w1264_,
		_w2124_,
		_w2127_,
		_w2128_,
		_w2129_
	);
	LUT3 #(
		.INIT('h35)
	) name1888 (
		\shift_data_reg[117]/NET0131 ,
		\wb_dat_i[21]_pad ,
		\wb_sel_i[2]_pad ,
		_w2130_
	);
	LUT3 #(
		.INIT('h08)
	) name1889 (
		_w804_,
		_w1057_,
		_w2130_,
		_w2131_
	);
	LUT2 #(
		.INIT('h8)
	) name1890 (
		_w1279_,
		_w2001_,
		_w2132_
	);
	LUT4 #(
		.INIT('hc888)
	) name1891 (
		\shift_data_reg[117]/NET0131 ,
		_w1060_,
		_w1279_,
		_w2001_,
		_w2133_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1892 (
		_w1165_,
		_w1262_,
		_w2132_,
		_w2133_,
		_w2134_
	);
	LUT2 #(
		.INIT('h2)
	) name1893 (
		\shift_data_reg[117]/NET0131 ,
		_w1283_,
		_w2135_
	);
	LUT4 #(
		.INIT('hff54)
	) name1894 (
		_w1264_,
		_w2131_,
		_w2134_,
		_w2135_,
		_w2136_
	);
	LUT3 #(
		.INIT('h35)
	) name1895 (
		\shift_data_reg[122]/NET0131 ,
		\wb_dat_i[26]_pad ,
		\wb_sel_i[3]_pad ,
		_w2137_
	);
	LUT3 #(
		.INIT('h08)
	) name1896 (
		_w804_,
		_w1057_,
		_w2137_,
		_w2138_
	);
	LUT3 #(
		.INIT('h20)
	) name1897 (
		_w1054_,
		_w1065_,
		_w1445_,
		_w2139_
	);
	LUT4 #(
		.INIT('h5155)
	) name1898 (
		\shift_data_reg[122]/NET0131 ,
		_w1054_,
		_w1065_,
		_w1445_,
		_w2140_
	);
	LUT2 #(
		.INIT('h2)
	) name1899 (
		_w1060_,
		_w2140_,
		_w2141_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1900 (
		_w1165_,
		_w1262_,
		_w2139_,
		_w2141_,
		_w2142_
	);
	LUT2 #(
		.INIT('h2)
	) name1901 (
		\shift_data_reg[122]/NET0131 ,
		_w1283_,
		_w2143_
	);
	LUT4 #(
		.INIT('hff54)
	) name1902 (
		_w1264_,
		_w2138_,
		_w2142_,
		_w2143_,
		_w2144_
	);
	LUT3 #(
		.INIT('h35)
	) name1903 (
		\shift_data_reg[127]/NET0131 ,
		\wb_dat_i[31]_pad ,
		\wb_sel_i[3]_pad ,
		_w2145_
	);
	LUT3 #(
		.INIT('h08)
	) name1904 (
		_w804_,
		_w1057_,
		_w2145_,
		_w2146_
	);
	LUT3 #(
		.INIT('h20)
	) name1905 (
		_w1054_,
		_w1065_,
		_w1491_,
		_w2147_
	);
	LUT4 #(
		.INIT('h5155)
	) name1906 (
		\shift_data_reg[127]/NET0131 ,
		_w1054_,
		_w1065_,
		_w1491_,
		_w2148_
	);
	LUT2 #(
		.INIT('h2)
	) name1907 (
		_w1060_,
		_w2148_,
		_w2149_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1908 (
		_w1165_,
		_w1262_,
		_w2147_,
		_w2149_,
		_w2150_
	);
	LUT2 #(
		.INIT('h2)
	) name1909 (
		\shift_data_reg[127]/NET0131 ,
		_w1283_,
		_w2151_
	);
	LUT4 #(
		.INIT('hff54)
	) name1910 (
		_w1264_,
		_w2146_,
		_w2150_,
		_w2151_,
		_w2152_
	);
	LUT3 #(
		.INIT('h80)
	) name1911 (
		_w804_,
		_w806_,
		_w1057_,
		_w2153_
	);
	LUT3 #(
		.INIT('h80)
	) name1912 (
		_w1278_,
		_w1279_,
		_w1361_,
		_w2154_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1913 (
		_w1060_,
		_w1165_,
		_w1262_,
		_w2154_,
		_w2155_
	);
	LUT4 #(
		.INIT('h1555)
	) name1914 (
		_w1059_,
		_w1278_,
		_w1279_,
		_w1361_,
		_w2156_
	);
	LUT3 #(
		.INIT('ha2)
	) name1915 (
		\shift_data_reg[100]/NET0131 ,
		_w1285_,
		_w2156_,
		_w2157_
	);
	LUT4 #(
		.INIT('hff54)
	) name1916 (
		_w1264_,
		_w2153_,
		_w2155_,
		_w2157_,
		_w2158_
	);
	LUT3 #(
		.INIT('h80)
	) name1917 (
		_w804_,
		_w818_,
		_w1057_,
		_w2159_
	);
	LUT3 #(
		.INIT('h20)
	) name1918 (
		_w1033_,
		_w1065_,
		_w1278_,
		_w2160_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1919 (
		_w1060_,
		_w1165_,
		_w1262_,
		_w2160_,
		_w2161_
	);
	LUT4 #(
		.INIT('h3133)
	) name1920 (
		_w1033_,
		_w1059_,
		_w1065_,
		_w1278_,
		_w2162_
	);
	LUT3 #(
		.INIT('ha2)
	) name1921 (
		\shift_data_reg[103]/NET0131 ,
		_w1285_,
		_w2162_,
		_w2163_
	);
	LUT4 #(
		.INIT('hff54)
	) name1922 (
		_w1264_,
		_w2159_,
		_w2161_,
		_w2163_,
		_w2164_
	);
	LUT3 #(
		.INIT('h35)
	) name1923 (
		\shift_data_reg[104]/NET0131 ,
		\wb_dat_i[8]_pad ,
		\wb_sel_i[1]_pad ,
		_w2165_
	);
	LUT3 #(
		.INIT('h08)
	) name1924 (
		_w804_,
		_w1057_,
		_w2165_,
		_w2166_
	);
	LUT4 #(
		.INIT('h1000)
	) name1925 (
		_w1032_,
		_w1065_,
		_w1278_,
		_w1306_,
		_w2167_
	);
	LUT3 #(
		.INIT('hc8)
	) name1926 (
		\shift_data_reg[104]/NET0131 ,
		_w1060_,
		_w2167_,
		_w2168_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1927 (
		_w1165_,
		_w1262_,
		_w2167_,
		_w2168_,
		_w2169_
	);
	LUT2 #(
		.INIT('h2)
	) name1928 (
		\shift_data_reg[104]/NET0131 ,
		_w1283_,
		_w2170_
	);
	LUT4 #(
		.INIT('hff54)
	) name1929 (
		_w1264_,
		_w2166_,
		_w2169_,
		_w2170_,
		_w2171_
	);
	LUT3 #(
		.INIT('h35)
	) name1930 (
		\shift_data_reg[106]/NET0131 ,
		\wb_dat_i[10]_pad ,
		\wb_sel_i[1]_pad ,
		_w2172_
	);
	LUT3 #(
		.INIT('h08)
	) name1931 (
		_w804_,
		_w1057_,
		_w2172_,
		_w2173_
	);
	LUT3 #(
		.INIT('h40)
	) name1932 (
		_w1065_,
		_w1278_,
		_w1445_,
		_w2174_
	);
	LUT4 #(
		.INIT('h4555)
	) name1933 (
		\shift_data_reg[106]/NET0131 ,
		_w1065_,
		_w1278_,
		_w1445_,
		_w2175_
	);
	LUT2 #(
		.INIT('h2)
	) name1934 (
		_w1060_,
		_w2175_,
		_w2176_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1935 (
		_w1165_,
		_w1262_,
		_w2174_,
		_w2176_,
		_w2177_
	);
	LUT2 #(
		.INIT('h2)
	) name1936 (
		\shift_data_reg[106]/NET0131 ,
		_w1283_,
		_w2178_
	);
	LUT4 #(
		.INIT('hff54)
	) name1937 (
		_w1264_,
		_w2173_,
		_w2177_,
		_w2178_,
		_w2179_
	);
	LUT3 #(
		.INIT('h35)
	) name1938 (
		\shift_data_reg[111]/NET0131 ,
		\wb_dat_i[15]_pad ,
		\wb_sel_i[1]_pad ,
		_w2180_
	);
	LUT3 #(
		.INIT('h08)
	) name1939 (
		_w804_,
		_w1057_,
		_w2180_,
		_w2181_
	);
	LUT4 #(
		.INIT('h0200)
	) name1940 (
		_w1025_,
		_w1032_,
		_w1065_,
		_w1278_,
		_w2182_
	);
	LUT3 #(
		.INIT('hc8)
	) name1941 (
		\shift_data_reg[111]/NET0131 ,
		_w1060_,
		_w2182_,
		_w2183_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1942 (
		_w1165_,
		_w1262_,
		_w2182_,
		_w2183_,
		_w2184_
	);
	LUT2 #(
		.INIT('h2)
	) name1943 (
		\shift_data_reg[111]/NET0131 ,
		_w1283_,
		_w2185_
	);
	LUT4 #(
		.INIT('hff54)
	) name1944 (
		_w1264_,
		_w2181_,
		_w2184_,
		_w2185_,
		_w2186_
	);
	LUT3 #(
		.INIT('h35)
	) name1945 (
		\shift_data_reg[112]/NET0131 ,
		\wb_dat_i[16]_pad ,
		\wb_sel_i[2]_pad ,
		_w2187_
	);
	LUT3 #(
		.INIT('h08)
	) name1946 (
		_w804_,
		_w1057_,
		_w2187_,
		_w2188_
	);
	LUT3 #(
		.INIT('h20)
	) name1947 (
		_w1054_,
		_w1065_,
		_w1369_,
		_w2189_
	);
	LUT4 #(
		.INIT('h5155)
	) name1948 (
		\shift_data_reg[112]/NET0131 ,
		_w1054_,
		_w1065_,
		_w1369_,
		_w2190_
	);
	LUT2 #(
		.INIT('h2)
	) name1949 (
		_w1060_,
		_w2190_,
		_w2191_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1950 (
		_w1165_,
		_w1262_,
		_w2189_,
		_w2191_,
		_w2192_
	);
	LUT2 #(
		.INIT('h2)
	) name1951 (
		\shift_data_reg[112]/NET0131 ,
		_w1283_,
		_w2193_
	);
	LUT4 #(
		.INIT('hff54)
	) name1952 (
		_w1264_,
		_w2188_,
		_w2192_,
		_w2193_,
		_w2194_
	);
	LUT3 #(
		.INIT('h35)
	) name1953 (
		\shift_data_reg[114]/NET0131 ,
		\wb_dat_i[18]_pad ,
		\wb_sel_i[2]_pad ,
		_w2195_
	);
	LUT3 #(
		.INIT('h08)
	) name1954 (
		_w804_,
		_w1057_,
		_w2195_,
		_w2196_
	);
	LUT3 #(
		.INIT('h20)
	) name1955 (
		_w1054_,
		_w1065_,
		_w1389_,
		_w2197_
	);
	LUT4 #(
		.INIT('h5155)
	) name1956 (
		\shift_data_reg[114]/NET0131 ,
		_w1054_,
		_w1065_,
		_w1389_,
		_w2198_
	);
	LUT2 #(
		.INIT('h2)
	) name1957 (
		_w1060_,
		_w2198_,
		_w2199_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1958 (
		_w1165_,
		_w1262_,
		_w2197_,
		_w2199_,
		_w2200_
	);
	LUT2 #(
		.INIT('h2)
	) name1959 (
		\shift_data_reg[114]/NET0131 ,
		_w1283_,
		_w2201_
	);
	LUT4 #(
		.INIT('hff54)
	) name1960 (
		_w1264_,
		_w2196_,
		_w2200_,
		_w2201_,
		_w2202_
	);
	LUT3 #(
		.INIT('h35)
	) name1961 (
		\shift_data_reg[119]/NET0131 ,
		\wb_dat_i[23]_pad ,
		\wb_sel_i[2]_pad ,
		_w2203_
	);
	LUT3 #(
		.INIT('h08)
	) name1962 (
		_w804_,
		_w1057_,
		_w2203_,
		_w2204_
	);
	LUT3 #(
		.INIT('h08)
	) name1963 (
		_w1033_,
		_w1054_,
		_w1065_,
		_w2205_
	);
	LUT4 #(
		.INIT('h5515)
	) name1964 (
		\shift_data_reg[119]/NET0131 ,
		_w1033_,
		_w1054_,
		_w1065_,
		_w2206_
	);
	LUT2 #(
		.INIT('h2)
	) name1965 (
		_w1060_,
		_w2206_,
		_w2207_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1966 (
		_w1165_,
		_w1262_,
		_w2205_,
		_w2207_,
		_w2208_
	);
	LUT2 #(
		.INIT('h2)
	) name1967 (
		\shift_data_reg[119]/NET0131 ,
		_w1283_,
		_w2209_
	);
	LUT4 #(
		.INIT('hff54)
	) name1968 (
		_w1264_,
		_w2204_,
		_w2208_,
		_w2209_,
		_w2210_
	);
	LUT3 #(
		.INIT('h35)
	) name1969 (
		\shift_data_reg[121]/NET0131 ,
		\wb_dat_i[25]_pad ,
		\wb_sel_i[3]_pad ,
		_w2211_
	);
	LUT3 #(
		.INIT('h08)
	) name1970 (
		_w804_,
		_w1057_,
		_w2211_,
		_w2212_
	);
	LUT4 #(
		.INIT('h0400)
	) name1971 (
		_w1032_,
		_w1054_,
		_w1065_,
		_w1352_,
		_w2213_
	);
	LUT3 #(
		.INIT('hc8)
	) name1972 (
		\shift_data_reg[121]/NET0131 ,
		_w1060_,
		_w2213_,
		_w2214_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1973 (
		_w1165_,
		_w1262_,
		_w2213_,
		_w2214_,
		_w2215_
	);
	LUT2 #(
		.INIT('h2)
	) name1974 (
		\shift_data_reg[121]/NET0131 ,
		_w1283_,
		_w2216_
	);
	LUT4 #(
		.INIT('hff54)
	) name1975 (
		_w1264_,
		_w2212_,
		_w2215_,
		_w2216_,
		_w2217_
	);
	LUT3 #(
		.INIT('h80)
	) name1976 (
		_w804_,
		_w889_,
		_w1057_,
		_w2218_
	);
	LUT3 #(
		.INIT('h40)
	) name1977 (
		_w1065_,
		_w1278_,
		_w1369_,
		_w2219_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1978 (
		_w1060_,
		_w1165_,
		_w1262_,
		_w2219_,
		_w2220_
	);
	LUT4 #(
		.INIT('h4555)
	) name1979 (
		_w1059_,
		_w1065_,
		_w1278_,
		_w1369_,
		_w2221_
	);
	LUT3 #(
		.INIT('ha2)
	) name1980 (
		\shift_data_reg[96]/NET0131 ,
		_w1285_,
		_w2221_,
		_w2222_
	);
	LUT4 #(
		.INIT('hff54)
	) name1981 (
		_w1264_,
		_w2218_,
		_w2220_,
		_w2222_,
		_w2223_
	);
	LUT3 #(
		.INIT('h80)
	) name1982 (
		_w804_,
		_w858_,
		_w1057_,
		_w2224_
	);
	LUT3 #(
		.INIT('h40)
	) name1983 (
		_w1065_,
		_w1278_,
		_w1379_,
		_w2225_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1984 (
		_w1060_,
		_w1165_,
		_w1262_,
		_w2225_,
		_w2226_
	);
	LUT4 #(
		.INIT('h4555)
	) name1985 (
		_w1059_,
		_w1065_,
		_w1278_,
		_w1379_,
		_w2227_
	);
	LUT3 #(
		.INIT('ha2)
	) name1986 (
		\shift_data_reg[97]/NET0131 ,
		_w1285_,
		_w2227_,
		_w2228_
	);
	LUT4 #(
		.INIT('hff54)
	) name1987 (
		_w1264_,
		_w2224_,
		_w2226_,
		_w2228_,
		_w2229_
	);
	LUT3 #(
		.INIT('h80)
	) name1988 (
		_w804_,
		_w833_,
		_w1057_,
		_w2230_
	);
	LUT3 #(
		.INIT('h80)
	) name1989 (
		_w1278_,
		_w1279_,
		_w1388_,
		_w2231_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1990 (
		_w1060_,
		_w1165_,
		_w1262_,
		_w2231_,
		_w2232_
	);
	LUT4 #(
		.INIT('h1555)
	) name1991 (
		_w1059_,
		_w1278_,
		_w1279_,
		_w1388_,
		_w2233_
	);
	LUT3 #(
		.INIT('ha2)
	) name1992 (
		\shift_data_reg[98]/NET0131 ,
		_w1285_,
		_w2233_,
		_w2234_
	);
	LUT4 #(
		.INIT('hff54)
	) name1993 (
		_w1264_,
		_w2230_,
		_w2232_,
		_w2234_,
		_w2235_
	);
	LUT3 #(
		.INIT('h80)
	) name1994 (
		_w804_,
		_w868_,
		_w1057_,
		_w2236_
	);
	LUT3 #(
		.INIT('h80)
	) name1995 (
		_w1278_,
		_w1279_,
		_w1398_,
		_w2237_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1996 (
		_w1060_,
		_w1165_,
		_w1262_,
		_w2237_,
		_w2238_
	);
	LUT4 #(
		.INIT('h1555)
	) name1997 (
		_w1059_,
		_w1278_,
		_w1279_,
		_w1398_,
		_w2239_
	);
	LUT3 #(
		.INIT('ha2)
	) name1998 (
		\shift_data_reg[99]/NET0131 ,
		_w1285_,
		_w2239_,
		_w2240_
	);
	LUT4 #(
		.INIT('hff54)
	) name1999 (
		_w1264_,
		_w2236_,
		_w2238_,
		_w2240_,
		_w2241_
	);
	LUT3 #(
		.INIT('h35)
	) name2000 (
		\shift_data_reg[123]/NET0131 ,
		\wb_dat_i[27]_pad ,
		\wb_sel_i[3]_pad ,
		_w2242_
	);
	LUT3 #(
		.INIT('h08)
	) name2001 (
		_w804_,
		_w1057_,
		_w2242_,
		_w2243_
	);
	LUT3 #(
		.INIT('h54)
	) name2002 (
		_w1032_,
		_w1062_,
		_w1064_,
		_w2244_
	);
	LUT2 #(
		.INIT('h8)
	) name2003 (
		_w1985_,
		_w2244_,
		_w2245_
	);
	LUT4 #(
		.INIT('hc888)
	) name2004 (
		\shift_data_reg[123]/NET0131 ,
		_w1060_,
		_w1985_,
		_w2244_,
		_w2246_
	);
	LUT4 #(
		.INIT('hbf00)
	) name2005 (
		_w1165_,
		_w1262_,
		_w2245_,
		_w2246_,
		_w2247_
	);
	LUT2 #(
		.INIT('h2)
	) name2006 (
		\shift_data_reg[123]/NET0131 ,
		_w1283_,
		_w2248_
	);
	LUT4 #(
		.INIT('hff54)
	) name2007 (
		_w1264_,
		_w2243_,
		_w2247_,
		_w2248_,
		_w2249_
	);
	LUT3 #(
		.INIT('h35)
	) name2008 (
		\shift_data_reg[124]/NET0131 ,
		\wb_dat_i[28]_pad ,
		\wb_sel_i[3]_pad ,
		_w2250_
	);
	LUT3 #(
		.INIT('h08)
	) name2009 (
		_w804_,
		_w1057_,
		_w2250_,
		_w2251_
	);
	LUT4 #(
		.INIT('h0400)
	) name2010 (
		_w1032_,
		_w1054_,
		_w1065_,
		_w1361_,
		_w2252_
	);
	LUT3 #(
		.INIT('hc8)
	) name2011 (
		\shift_data_reg[124]/NET0131 ,
		_w1060_,
		_w2252_,
		_w2253_
	);
	LUT4 #(
		.INIT('hbf00)
	) name2012 (
		_w1165_,
		_w1262_,
		_w2252_,
		_w2253_,
		_w2254_
	);
	LUT2 #(
		.INIT('h2)
	) name2013 (
		\shift_data_reg[124]/NET0131 ,
		_w1283_,
		_w2255_
	);
	LUT4 #(
		.INIT('hff54)
	) name2014 (
		_w1264_,
		_w2251_,
		_w2254_,
		_w2255_,
		_w2256_
	);
	LUT3 #(
		.INIT('h35)
	) name2015 (
		\shift_data_reg[125]/NET0131 ,
		\wb_dat_i[29]_pad ,
		\wb_sel_i[3]_pad ,
		_w2257_
	);
	LUT3 #(
		.INIT('h08)
	) name2016 (
		_w804_,
		_w1057_,
		_w2257_,
		_w2258_
	);
	LUT2 #(
		.INIT('h8)
	) name2017 (
		_w2001_,
		_w2244_,
		_w2259_
	);
	LUT4 #(
		.INIT('hc888)
	) name2018 (
		\shift_data_reg[125]/NET0131 ,
		_w1060_,
		_w2001_,
		_w2244_,
		_w2260_
	);
	LUT4 #(
		.INIT('hbf00)
	) name2019 (
		_w1165_,
		_w1262_,
		_w2259_,
		_w2260_,
		_w2261_
	);
	LUT2 #(
		.INIT('h2)
	) name2020 (
		\shift_data_reg[125]/NET0131 ,
		_w1283_,
		_w2262_
	);
	LUT4 #(
		.INIT('hff54)
	) name2021 (
		_w1264_,
		_w2258_,
		_w2261_,
		_w2262_,
		_w2263_
	);
	LUT3 #(
		.INIT('h35)
	) name2022 (
		\shift_data_reg[126]/NET0131 ,
		\wb_dat_i[30]_pad ,
		\wb_sel_i[3]_pad ,
		_w2264_
	);
	LUT3 #(
		.INIT('h08)
	) name2023 (
		_w804_,
		_w1057_,
		_w2264_,
		_w2265_
	);
	LUT4 #(
		.INIT('h0400)
	) name2024 (
		_w1032_,
		_w1054_,
		_w1065_,
		_w1297_,
		_w2266_
	);
	LUT3 #(
		.INIT('hc8)
	) name2025 (
		\shift_data_reg[126]/NET0131 ,
		_w1060_,
		_w2266_,
		_w2267_
	);
	LUT4 #(
		.INIT('hbf00)
	) name2026 (
		_w1165_,
		_w1262_,
		_w2266_,
		_w2267_,
		_w2268_
	);
	LUT2 #(
		.INIT('h2)
	) name2027 (
		\shift_data_reg[126]/NET0131 ,
		_w1283_,
		_w2269_
	);
	LUT4 #(
		.INIT('hff54)
	) name2028 (
		_w1264_,
		_w2265_,
		_w2268_,
		_w2269_,
		_w2270_
	);
	LUT3 #(
		.INIT('h2f)
	) name2029 (
		\ctrl_reg[13]/NET0131 ,
		\shift_tip_reg/NET0131 ,
		\ss_reg[0]/NET0131 ,
		_w2271_
	);
	LUT3 #(
		.INIT('h2f)
	) name2030 (
		\ctrl_reg[13]/NET0131 ,
		\shift_tip_reg/NET0131 ,
		\ss_reg[1]/NET0131 ,
		_w2272_
	);
	LUT3 #(
		.INIT('h2f)
	) name2031 (
		\ctrl_reg[13]/NET0131 ,
		\shift_tip_reg/NET0131 ,
		\ss_reg[2]/NET0131 ,
		_w2273_
	);
	LUT3 #(
		.INIT('h2f)
	) name2032 (
		\ctrl_reg[13]/NET0131 ,
		\shift_tip_reg/NET0131 ,
		\ss_reg[3]/NET0131 ,
		_w2274_
	);
	LUT3 #(
		.INIT('h2f)
	) name2033 (
		\ctrl_reg[13]/NET0131 ,
		\shift_tip_reg/NET0131 ,
		\ss_reg[4]/NET0131 ,
		_w2275_
	);
	LUT3 #(
		.INIT('h2f)
	) name2034 (
		\ctrl_reg[13]/NET0131 ,
		\shift_tip_reg/NET0131 ,
		\ss_reg[5]/NET0131 ,
		_w2276_
	);
	LUT3 #(
		.INIT('h2f)
	) name2035 (
		\ctrl_reg[13]/NET0131 ,
		\shift_tip_reg/NET0131 ,
		\ss_reg[6]/NET0131 ,
		_w2277_
	);
	LUT3 #(
		.INIT('h2f)
	) name2036 (
		\ctrl_reg[13]/NET0131 ,
		\shift_tip_reg/NET0131 ,
		\ss_reg[7]/NET0131 ,
		_w2278_
	);
	assign \_al_n1  = 1'b1;
	assign \g10384/_0_  = _w539_ ;
	assign \g10421/_0_  = _w554_ ;
	assign \g10487/_0_  = _w556_ ;
	assign \g10622/_0_  = _w559_ ;
	assign \g10625/_0_  = _w561_ ;
	assign \g10631/_3_  = _w562_ ;
	assign \g10641/_0_  = _w568_ ;
	assign \g10677/_3_  = _w570_ ;
	assign \g10695/_0_  = _w573_ ;
	assign \g10699/_3_  = _w577_ ;
	assign \g10796/_0_  = _w579_ ;
	assign \g10814/_00_  = _w582_ ;
	assign \g10815/_0_  = _w591_ ;
	assign \g10819/_0_  = _w595_ ;
	assign \g10821/_0_  = _w598_ ;
	assign \g10824/_3_  = _w600_ ;
	assign \g10858/_0_  = _w604_ ;
	assign \g11042/_00_  = _w606_ ;
	assign \g11067/_0_  = _w616_ ;
	assign \g11071/_00_  = _w618_ ;
	assign \g11074/_0_  = _w620_ ;
	assign \g11075/_0_  = _w624_ ;
	assign \g11076/_0_  = _w626_ ;
	assign \g11077/_0_  = _w630_ ;
	assign \g11078/_0_  = _w634_ ;
	assign \g11079/_0_  = _w637_ ;
	assign \g11080/_0_  = _w639_ ;
	assign \g11149/_0_  = _w643_ ;
	assign \g11151/_0_  = _w647_ ;
	assign \g11190/_00_  = _w650_ ;
	assign \g11297/_0_  = _w660_ ;
	assign \g11298/_0_  = _w670_ ;
	assign \g11300/_0_  = _w679_ ;
	assign \g11301/_0_  = _w688_ ;
	assign \g11303/_0_  = _w697_ ;
	assign \g11346/_0_  = _w706_ ;
	assign \g11347/_0_  = _w715_ ;
	assign \g11348/_0_  = _w724_ ;
	assign \g11358/_0_  = _w734_ ;
	assign \g11359/_0_  = _w744_ ;
	assign \g11360/_0_  = _w754_ ;
	assign \g11361/_0_  = _w764_ ;
	assign \g11362/_0_  = _w774_ ;
	assign \g11363/_0_  = _w784_ ;
	assign \g11470/_0_  = _w792_ ;
	assign \g11499/_0_  = _w800_ ;
	assign \g11501/_0_  = _w801_ ;
	assign \g11502/_0_  = _w803_ ;
	assign \g11503/_0_  = _w808_ ;
	assign \g11504/_0_  = _w812_ ;
	assign \g11505/_0_  = _w816_ ;
	assign \g11506/_0_  = _w820_ ;
	assign \g11507/_0_  = _w824_ ;
	assign \g11508/_0_  = _w828_ ;
	assign \g11509/_0_  = _w831_ ;
	assign \g11510/_0_  = _w835_ ;
	assign \g11511/_0_  = _w838_ ;
	assign \g11512/_0_  = _w842_ ;
	assign \g11513/_0_  = _w846_ ;
	assign \g11514/_0_  = _w850_ ;
	assign \g11515/_0_  = _w853_ ;
	assign \g11516/_0_  = _w856_ ;
	assign \g11517/_0_  = _w860_ ;
	assign \g11519/_0_  = _w863_ ;
	assign \g11520/_0_  = _w866_ ;
	assign \g11521/_0_  = _w870_ ;
	assign \g11522/_0_  = _w873_ ;
	assign \g11523/_0_  = _w876_ ;
	assign \g11524/_0_  = _w880_ ;
	assign \g11525/_0_  = _w883_ ;
	assign \g11526/_0_  = _w887_ ;
	assign \g11527/_0_  = _w891_ ;
	assign \g11528/_0_  = _w894_ ;
	assign \g11529/_0_  = _w897_ ;
	assign \g11530/_0_  = _w901_ ;
	assign \g11531/_0_  = _w904_ ;
	assign \g11532/_0_  = _w907_ ;
	assign \g11533/_0_  = _w910_ ;
	assign \g11534/_0_  = _w913_ ;
	assign \g11535/_0_  = _w916_ ;
	assign \g11536/_0_  = _w919_ ;
	assign \g11537/_0_  = _w922_ ;
	assign \g11538/_0_  = _w925_ ;
	assign \g11539/_0_  = _w928_ ;
	assign \g11655/_0_  = _w933_ ;
	assign \g11658/_0_  = _w938_ ;
	assign \g11659/_0_  = _w943_ ;
	assign \g11661/_0_  = _w948_ ;
	assign \g11662/_0_  = _w953_ ;
	assign \g11680/_0_  = _w958_ ;
	assign \g11723/_0_  = _w963_ ;
	assign \g11726/_0_  = _w968_ ;
	assign \g11730/_0_  = _w973_ ;
	assign \g11739/_0_  = _w978_ ;
	assign \g11750/_0_  = _w983_ ;
	assign \g11759/_0_  = _w988_ ;
	assign \g11760/_0_  = _w993_ ;
	assign \g11761/_0_  = _w998_ ;
	assign \g11764/_0_  = _w1003_ ;
	assign \g11765/_0_  = _w1008_ ;
	assign \g12212/_0_  = _w1009_ ;
	assign \g13497/_0_  = _w1274_ ;
	assign \g13884/_0_  = _w1287_ ;
	assign \g13982/_0_  = _w1295_ ;
	assign \g13999/_0_  = _w1304_ ;
	assign \g9305/_0_  = _w1316_ ;
	assign \g9306/_0_  = _w1324_ ;
	assign \g9307/_0_  = _w1335_ ;
	assign \g9308/_0_  = _w1344_ ;
	assign \g9309/_0_  = _w1357_ ;
	assign \g9310/_0_  = _w1366_ ;
	assign \g9346/_0_  = _w1376_ ;
	assign \g9347/_0_  = _w1385_ ;
	assign \g9348/_0_  = _w1395_ ;
	assign \g9349/_0_  = _w1403_ ;
	assign \g9350/_0_  = _w1412_ ;
	assign \g9351/_0_  = _w1419_ ;
	assign \g9352/_0_  = _w1426_ ;
	assign \g9353/_0_  = _w1435_ ;
	assign \g9354/_0_  = _w1442_ ;
	assign \g9355/_0_  = _w1451_ ;
	assign \g9356/_0_  = _w1458_ ;
	assign \g9357/_0_  = _w1467_ ;
	assign \g9358/_0_  = _w1474_ ;
	assign \g9359/_0_  = _w1481_ ;
	assign \g9360/_0_  = _w1488_ ;
	assign \g9361/_0_  = _w1497_ ;
	assign \g9362/_0_  = _w1506_ ;
	assign \g9363/_0_  = _w1515_ ;
	assign \g9364/_0_  = _w1523_ ;
	assign \g9365/_0_  = _w1531_ ;
	assign \g9366/_0_  = _w1540_ ;
	assign \g9367/_0_  = _w1548_ ;
	assign \g9368/_0_  = _w1556_ ;
	assign \g9369/_0_  = _w1563_ ;
	assign \g9370/_0_  = _w1571_ ;
	assign \g9371/_0_  = _w1579_ ;
	assign \g9372/_0_  = _w1587_ ;
	assign \g9373/_0_  = _w1595_ ;
	assign \g9374/_0_  = _w1603_ ;
	assign \g9375/_0_  = _w1611_ ;
	assign \g9380/_0_  = _w1619_ ;
	assign \g9381/_0_  = _w1625_ ;
	assign \g9382/_0_  = _w1631_ ;
	assign \g9383/_0_  = _w1637_ ;
	assign \g9384/_0_  = _w1643_ ;
	assign \g9385/_0_  = _w1652_ ;
	assign \g9386/_0_  = _w1658_ ;
	assign \g9387/_0_  = _w1664_ ;
	assign \g9388/_0_  = _w1672_ ;
	assign \g9389/_0_  = _w1681_ ;
	assign \g9390/_0_  = _w1689_ ;
	assign \g9391/_0_  = _w1697_ ;
	assign \g9392/_0_  = _w1706_ ;
	assign \g9393/_0_  = _w1715_ ;
	assign \g9394/_0_  = _w1722_ ;
	assign \g9395/_0_  = _w1728_ ;
	assign \g9396/_0_  = _w1737_ ;
	assign \g9397/_0_  = _w1744_ ;
	assign \g9398/_0_  = _w1753_ ;
	assign \g9399/_0_  = _w1760_ ;
	assign \g9400/_0_  = _w1767_ ;
	assign \g9401/_0_  = _w1776_ ;
	assign \g9402/_0_  = _w1785_ ;
	assign \g9403/_0_  = _w1792_ ;
	assign \g9404/_0_  = _w1798_ ;
	assign \g9405/_0_  = _w1804_ ;
	assign \g9406/_0_  = _w1813_ ;
	assign \g9407/_0_  = _w1819_ ;
	assign \g9408/_0_  = _w1825_ ;
	assign \g9409/_0_  = _w1831_ ;
	assign \g9410/_0_  = _w1840_ ;
	assign \g9411/_0_  = _w1847_ ;
	assign \g9439/_0_  = _w1855_ ;
	assign \g9440/_0_  = _w1863_ ;
	assign \g9441/_0_  = _w1871_ ;
	assign \g9442/_0_  = _w1879_ ;
	assign \g9443/_0_  = _w1887_ ;
	assign \g9444/_0_  = _w1895_ ;
	assign \g9445/_0_  = _w1904_ ;
	assign \g9446/_0_  = _w1912_ ;
	assign \g9447/_0_  = _w1920_ ;
	assign \g9448/_0_  = _w1928_ ;
	assign \g9449/_0_  = _w1936_ ;
	assign \g9450/_0_  = _w1944_ ;
	assign \g9451/_0_  = _w1952_ ;
	assign \g9452/_0_  = _w1960_ ;
	assign \g9453/_0_  = _w1968_ ;
	assign \g9454/_0_  = _w1976_ ;
	assign \g9455/_0_  = _w1984_ ;
	assign \g9456/_0_  = _w1992_ ;
	assign \g9457/_0_  = _w2000_ ;
	assign \g9458/_0_  = _w2008_ ;
	assign \g9459/_0_  = _w2016_ ;
	assign \g9461/_0_  = _w2024_ ;
	assign \g9462/_0_  = _w2032_ ;
	assign \g9463/_0_  = _w2039_ ;
	assign \g9464/_0_  = _w2047_ ;
	assign \g9465/_0_  = _w2054_ ;
	assign \g9466/_0_  = _w2061_ ;
	assign \g9529/_0_  = _w2068_ ;
	assign \g9530/_0_  = _w2076_ ;
	assign \g9531/_0_  = _w2083_ ;
	assign \g9532/_0_  = _w2091_ ;
	assign \g9535/_0_  = _w2100_ ;
	assign \g9542/_0_  = _w2106_ ;
	assign \g9543/_0_  = _w2113_ ;
	assign \g9546/_0_  = _w2122_ ;
	assign \g9547/_0_  = _w2129_ ;
	assign \g9548/_0_  = _w2136_ ;
	assign \g9549/_0_  = _w2144_ ;
	assign \g9550/_0_  = _w2152_ ;
	assign \g9551/_0_  = _w2158_ ;
	assign \g9552/_0_  = _w2164_ ;
	assign \g9553/_0_  = _w2171_ ;
	assign \g9559/_0_  = _w2179_ ;
	assign \g9568/_0_  = _w2186_ ;
	assign \g9571/_0_  = _w2194_ ;
	assign \g9573/_0_  = _w2202_ ;
	assign \g9583/_0_  = _w2210_ ;
	assign \g9589/_0_  = _w2217_ ;
	assign \g9590/_0_  = _w2223_ ;
	assign \g9591/_0_  = _w2229_ ;
	assign \g9592/_0_  = _w2235_ ;
	assign \g9593/_0_  = _w2241_ ;
	assign \g9594/_0_  = _w2249_ ;
	assign \g9595/_0_  = _w2256_ ;
	assign \g9596/_0_  = _w2263_ ;
	assign \g9597/_0_  = _w2270_ ;
	assign \ss_pad_o[0]_pad  = _w2271_ ;
	assign \ss_pad_o[1]_pad  = _w2272_ ;
	assign \ss_pad_o[2]_pad  = _w2273_ ;
	assign \ss_pad_o[3]_pad  = _w2274_ ;
	assign \ss_pad_o[4]_pad  = _w2275_ ;
	assign \ss_pad_o[5]_pad  = _w2276_ ;
	assign \ss_pad_o[6]_pad  = _w2277_ ;
	assign \ss_pad_o[7]_pad  = _w2278_ ;
	assign wb_err_o_pad = 1'b0;
endmodule;