module top( a_pad , b_pad , c_pad , d_pad , e_pad , f_pad , g_pad , h_pad , i_pad , j_pad , k_pad , l_pad , m_pad , n_pad , o_pad , p_pad , q_pad , r_pad , s_pad , t_pad , u_pad );
  input a_pad ;
  input b_pad ;
  input c_pad ;
  input d_pad ;
  input e_pad ;
  output f_pad ;
  output g_pad ;
  output h_pad ;
  output i_pad ;
  output j_pad ;
  output k_pad ;
  output l_pad ;
  output m_pad ;
  output n_pad ;
  output o_pad ;
  output p_pad ;
  output q_pad ;
  output r_pad ;
  output s_pad ;
  output t_pad ;
  output u_pad ;
  wire n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 ;
  assign n6 = a_pad & e_pad ;
  assign n7 = c_pad & d_pad ;
  assign n8 = b_pad & n7 ;
  assign n9 = n6 & n8 ;
  assign n10 = c_pad & ~d_pad ;
  assign n11 = b_pad & n10 ;
  assign n12 = n6 & n11 ;
  assign n13 = ~c_pad & d_pad ;
  assign n14 = b_pad & n13 ;
  assign n15 = n6 & n14 ;
  assign n16 = ~c_pad & ~d_pad ;
  assign n17 = b_pad & n16 ;
  assign n18 = n6 & n17 ;
  assign n19 = ~b_pad & n7 ;
  assign n20 = n6 & n19 ;
  assign n21 = ~b_pad & n10 ;
  assign n22 = n6 & n21 ;
  assign n23 = ~b_pad & n13 ;
  assign n24 = n6 & n23 ;
  assign n25 = ~b_pad & n16 ;
  assign n26 = n6 & n25 ;
  assign n27 = ~a_pad & e_pad ;
  assign n28 = n8 & n27 ;
  assign n29 = n11 & n27 ;
  assign n30 = n14 & n27 ;
  assign n31 = n17 & n27 ;
  assign n32 = n19 & n27 ;
  assign n33 = n21 & n27 ;
  assign n34 = n23 & n27 ;
  assign n35 = n25 & n27 ;
  assign f_pad = n9 ;
  assign g_pad = n12 ;
  assign h_pad = n15 ;
  assign i_pad = n18 ;
  assign j_pad = n20 ;
  assign k_pad = n22 ;
  assign l_pad = n24 ;
  assign m_pad = n26 ;
  assign n_pad = n28 ;
  assign o_pad = n29 ;
  assign p_pad = n30 ;
  assign q_pad = n31 ;
  assign r_pad = n32 ;
  assign s_pad = n33 ;
  assign t_pad = n34 ;
  assign u_pad = n35 ;
endmodule
