module top (\a0_pad , a_pad, \b0_pad , b_pad, \c0_pad , c_pad, \d0_pad , d_pad, \e0_pad , e_pad, \f0_pad , f_pad, g_pad, h_pad, i_pad, j_pad, k_pad, l_pad, m_pad, n_pad, o_pad, p_pad, q_pad, r_pad, s_pad, t_pad, u_pad, v_pad, w_pad, x_pad, y_pad, z_pad, \g0_pad , \h0_pad , \i0_pad );
	input \a0_pad  ;
	input a_pad ;
	input \b0_pad  ;
	input b_pad ;
	input \c0_pad  ;
	input c_pad ;
	input \d0_pad  ;
	input d_pad ;
	input \e0_pad  ;
	input e_pad ;
	input \f0_pad  ;
	input f_pad ;
	input g_pad ;
	input h_pad ;
	input i_pad ;
	input j_pad ;
	input k_pad ;
	input l_pad ;
	input m_pad ;
	input n_pad ;
	input o_pad ;
	input p_pad ;
	input q_pad ;
	input r_pad ;
	input s_pad ;
	input t_pad ;
	input u_pad ;
	input v_pad ;
	input w_pad ;
	input x_pad ;
	input y_pad ;
	input z_pad ;
	output \g0_pad  ;
	output \h0_pad  ;
	output \i0_pad  ;
	wire _w68_ ;
	wire _w67_ ;
	wire _w66_ ;
	wire _w65_ ;
	wire _w64_ ;
	wire _w63_ ;
	wire _w46_ ;
	wire _w45_ ;
	wire _w44_ ;
	wire _w43_ ;
	wire _w42_ ;
	wire _w41_ ;
	wire _w40_ ;
	wire _w39_ ;
	wire _w38_ ;
	wire _w37_ ;
	wire _w36_ ;
	wire _w35_ ;
	wire _w34_ ;
	wire _w47_ ;
	wire _w48_ ;
	wire _w49_ ;
	wire _w50_ ;
	wire _w51_ ;
	wire _w52_ ;
	wire _w53_ ;
	wire _w54_ ;
	wire _w55_ ;
	wire _w56_ ;
	wire _w57_ ;
	wire _w58_ ;
	wire _w59_ ;
	wire _w60_ ;
	wire _w61_ ;
	wire _w62_ ;
	LUT2 #(
		.INIT('h4)
	) name0 (
		i_pad,
		y_pad,
		_w34_
	);
	LUT4 #(
		.INIT('hf531)
	) name1 (
		\b0_pad ,
		\c0_pad ,
		l_pad,
		m_pad,
		_w35_
	);
	LUT2 #(
		.INIT('h4)
	) name2 (
		_w34_,
		_w35_,
		_w36_
	);
	LUT4 #(
		.INIT('h8caf)
	) name3 (
		\a0_pad ,
		\b0_pad ,
		k_pad,
		l_pad,
		_w37_
	);
	LUT4 #(
		.INIT('hf531)
	) name4 (
		i_pad,
		j_pad,
		y_pad,
		z_pad,
		_w38_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name5 (
		\a0_pad ,
		j_pad,
		k_pad,
		z_pad,
		_w39_
	);
	LUT3 #(
		.INIT('h80)
	) name6 (
		_w38_,
		_w39_,
		_w37_,
		_w40_
	);
	LUT4 #(
		.INIT('h8caf)
	) name7 (
		\e0_pad ,
		\f0_pad ,
		o_pad,
		p_pad,
		_w41_
	);
	LUT4 #(
		.INIT('hf531)
	) name8 (
		\d0_pad ,
		\e0_pad ,
		n_pad,
		o_pad,
		_w42_
	);
	LUT4 #(
		.INIT('h8caf)
	) name9 (
		\c0_pad ,
		\d0_pad ,
		m_pad,
		n_pad,
		_w43_
	);
	LUT3 #(
		.INIT('hb0)
	) name10 (
		_w41_,
		_w42_,
		_w43_,
		_w44_
	);
	LUT4 #(
		.INIT('h1131)
	) name11 (
		_w38_,
		_w34_,
		_w39_,
		_w37_,
		_w45_
	);
	LUT4 #(
		.INIT('h00f7)
	) name12 (
		_w36_,
		_w40_,
		_w44_,
		_w45_,
		_w46_
	);
	LUT2 #(
		.INIT('h4)
	) name13 (
		a_pad,
		q_pad,
		_w47_
	);
	LUT4 #(
		.INIT('hf531)
	) name14 (
		a_pad,
		b_pad,
		q_pad,
		r_pad,
		_w48_
	);
	LUT4 #(
		.INIT('hf531)
	) name15 (
		c_pad,
		d_pad,
		s_pad,
		t_pad,
		_w49_
	);
	LUT4 #(
		.INIT('h8caf)
	) name16 (
		b_pad,
		c_pad,
		r_pad,
		s_pad,
		_w50_
	);
	LUT4 #(
		.INIT('h1311)
	) name17 (
		_w48_,
		_w47_,
		_w49_,
		_w50_,
		_w51_
	);
	LUT2 #(
		.INIT('h4)
	) name18 (
		e_pad,
		u_pad,
		_w52_
	);
	LUT4 #(
		.INIT('hf531)
	) name19 (
		e_pad,
		f_pad,
		u_pad,
		v_pad,
		_w53_
	);
	LUT4 #(
		.INIT('hf531)
	) name20 (
		g_pad,
		h_pad,
		w_pad,
		x_pad,
		_w54_
	);
	LUT4 #(
		.INIT('h8caf)
	) name21 (
		f_pad,
		g_pad,
		v_pad,
		w_pad,
		_w55_
	);
	LUT4 #(
		.INIT('h1511)
	) name22 (
		_w52_,
		_w53_,
		_w54_,
		_w55_,
		_w56_
	);
	LUT4 #(
		.INIT('h8caf)
	) name23 (
		a_pad,
		d_pad,
		q_pad,
		t_pad,
		_w57_
	);
	LUT4 #(
		.INIT('h8000)
	) name24 (
		_w48_,
		_w49_,
		_w50_,
		_w57_,
		_w58_
	);
	LUT4 #(
		.INIT('h8caf)
	) name25 (
		e_pad,
		h_pad,
		u_pad,
		x_pad,
		_w59_
	);
	LUT4 #(
		.INIT('h8000)
	) name26 (
		_w53_,
		_w54_,
		_w55_,
		_w59_,
		_w60_
	);
	LUT4 #(
		.INIT('h0400)
	) name27 (
		_w56_,
		_w58_,
		_w51_,
		_w60_,
		_w61_
	);
	LUT3 #(
		.INIT('h07)
	) name28 (
		_w56_,
		_w58_,
		_w51_,
		_w62_
	);
	LUT3 #(
		.INIT('h4f)
	) name29 (
		_w46_,
		_w61_,
		_w62_,
		_w63_
	);
	LUT2 #(
		.INIT('h2)
	) name30 (
		\f0_pad ,
		p_pad,
		_w64_
	);
	LUT4 #(
		.INIT('h0080)
	) name31 (
		_w41_,
		_w42_,
		_w43_,
		_w64_,
		_w65_
	);
	LUT4 #(
		.INIT('h0800)
	) name32 (
		_w36_,
		_w40_,
		_w45_,
		_w65_,
		_w66_
	);
	LUT2 #(
		.INIT('h8)
	) name33 (
		_w61_,
		_w66_,
		_w67_
	);
	LUT4 #(
		.INIT('h30b0)
	) name34 (
		_w46_,
		_w61_,
		_w62_,
		_w66_,
		_w68_
	);
	assign \g0_pad  = _w68_ ;
	assign \h0_pad  = _w67_ ;
	assign \i0_pad  = _w63_ ;
endmodule;