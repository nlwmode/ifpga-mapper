module top (a_pad, b_pad, d_pad, \e0_pad , f_pad, \g0_pad , g_pad, h_pad, i_pad, j_pad, k_pad, l_pad, m_pad, n_pad, o_pad, p_pad, q_pad, r_pad, s_pad, \a0_pad , \b0_pad , \c0_pad , \d0_pad , \f0_pad , \h0_pad , t_pad, u_pad, v_pad, w_pad, x_pad, y_pad, z_pad);
	input a_pad ;
	input b_pad ;
	input d_pad ;
	input \e0_pad  ;
	input f_pad ;
	input \g0_pad  ;
	input g_pad ;
	input h_pad ;
	input i_pad ;
	input j_pad ;
	input k_pad ;
	input l_pad ;
	input m_pad ;
	input n_pad ;
	input o_pad ;
	input p_pad ;
	input q_pad ;
	input r_pad ;
	input s_pad ;
	output \a0_pad  ;
	output \b0_pad  ;
	output \c0_pad  ;
	output \d0_pad  ;
	output \f0_pad  ;
	output \h0_pad  ;
	output t_pad ;
	output u_pad ;
	output v_pad ;
	output w_pad ;
	output x_pad ;
	output y_pad ;
	output z_pad ;
	wire _w71_ ;
	wire _w70_ ;
	wire _w69_ ;
	wire _w68_ ;
	wire _w67_ ;
	wire _w66_ ;
	wire _w65_ ;
	wire _w64_ ;
	wire _w63_ ;
	wire _w62_ ;
	wire _w61_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w56_ ;
	wire _w55_ ;
	wire _w54_ ;
	wire _w53_ ;
	wire _w52_ ;
	wire _w51_ ;
	wire _w50_ ;
	wire _w49_ ;
	wire _w32_ ;
	wire _w31_ ;
	wire _w30_ ;
	wire _w29_ ;
	wire _w28_ ;
	wire _w27_ ;
	wire _w26_ ;
	wire _w25_ ;
	wire _w24_ ;
	wire _w23_ ;
	wire _w22_ ;
	wire _w21_ ;
	wire _w20_ ;
	wire _w33_ ;
	wire _w34_ ;
	wire _w35_ ;
	wire _w36_ ;
	wire _w37_ ;
	wire _w38_ ;
	wire _w39_ ;
	wire _w40_ ;
	wire _w41_ ;
	wire _w42_ ;
	wire _w43_ ;
	wire _w44_ ;
	wire _w45_ ;
	wire _w46_ ;
	wire _w47_ ;
	wire _w48_ ;
	LUT2 #(
		.INIT('h8)
	) name0 (
		g_pad,
		h_pad,
		_w20_
	);
	LUT2 #(
		.INIT('h8)
	) name1 (
		i_pad,
		_w20_,
		_w21_
	);
	LUT2 #(
		.INIT('h4)
	) name2 (
		j_pad,
		_w21_,
		_w22_
	);
	LUT2 #(
		.INIT('h1)
	) name3 (
		k_pad,
		l_pad,
		_w23_
	);
	LUT2 #(
		.INIT('h8)
	) name4 (
		_w22_,
		_w23_,
		_w24_
	);
	LUT2 #(
		.INIT('h4)
	) name5 (
		k_pad,
		_w22_,
		_w25_
	);
	LUT2 #(
		.INIT('h2)
	) name6 (
		l_pad,
		_w25_,
		_w26_
	);
	LUT2 #(
		.INIT('h4)
	) name7 (
		d_pad,
		\e0_pad ,
		_w27_
	);
	LUT2 #(
		.INIT('h2)
	) name8 (
		q_pad,
		_w27_,
		_w28_
	);
	LUT2 #(
		.INIT('h2)
	) name9 (
		\g0_pad ,
		_w28_,
		_w29_
	);
	LUT2 #(
		.INIT('h4)
	) name10 (
		_w24_,
		_w29_,
		_w30_
	);
	LUT2 #(
		.INIT('h4)
	) name11 (
		_w26_,
		_w30_,
		_w31_
	);
	LUT2 #(
		.INIT('h4)
	) name12 (
		m_pad,
		_w24_,
		_w32_
	);
	LUT2 #(
		.INIT('h2)
	) name13 (
		m_pad,
		_w24_,
		_w33_
	);
	LUT2 #(
		.INIT('h2)
	) name14 (
		_w29_,
		_w32_,
		_w34_
	);
	LUT2 #(
		.INIT('h4)
	) name15 (
		_w33_,
		_w34_,
		_w35_
	);
	LUT2 #(
		.INIT('h2)
	) name16 (
		n_pad,
		_w32_,
		_w36_
	);
	LUT2 #(
		.INIT('h1)
	) name17 (
		m_pad,
		n_pad,
		_w37_
	);
	LUT2 #(
		.INIT('h8)
	) name18 (
		_w23_,
		_w37_,
		_w38_
	);
	LUT2 #(
		.INIT('h8)
	) name19 (
		_w22_,
		_w38_,
		_w39_
	);
	LUT2 #(
		.INIT('h2)
	) name20 (
		_w29_,
		_w39_,
		_w40_
	);
	LUT2 #(
		.INIT('h4)
	) name21 (
		_w36_,
		_w40_,
		_w41_
	);
	LUT2 #(
		.INIT('h8)
	) name22 (
		o_pad,
		_w28_,
		_w42_
	);
	LUT2 #(
		.INIT('h1)
	) name23 (
		a_pad,
		_w38_,
		_w43_
	);
	LUT2 #(
		.INIT('h2)
	) name24 (
		_w22_,
		_w28_,
		_w44_
	);
	LUT2 #(
		.INIT('h4)
	) name25 (
		_w43_,
		_w44_,
		_w45_
	);
	LUT2 #(
		.INIT('h1)
	) name26 (
		_w42_,
		_w45_,
		_w46_
	);
	LUT2 #(
		.INIT('h2)
	) name27 (
		\g0_pad ,
		_w46_,
		_w47_
	);
	LUT2 #(
		.INIT('h4)
	) name28 (
		\e0_pad ,
		q_pad,
		_w48_
	);
	LUT2 #(
		.INIT('h1)
	) name29 (
		d_pad,
		_w48_,
		_w49_
	);
	LUT2 #(
		.INIT('h2)
	) name30 (
		\g0_pad ,
		_w49_,
		_w50_
	);
	LUT2 #(
		.INIT('h8)
	) name31 (
		\g0_pad ,
		r_pad,
		_w51_
	);
	LUT2 #(
		.INIT('h8)
	) name32 (
		b_pad,
		\e0_pad ,
		_w52_
	);
	LUT2 #(
		.INIT('h4)
	) name33 (
		b_pad,
		o_pad,
		_w53_
	);
	LUT2 #(
		.INIT('h1)
	) name34 (
		_w52_,
		_w53_,
		_w54_
	);
	LUT2 #(
		.INIT('h4)
	) name35 (
		p_pad,
		s_pad,
		_w55_
	);
	LUT2 #(
		.INIT('h1)
	) name36 (
		f_pad,
		_w55_,
		_w56_
	);
	LUT2 #(
		.INIT('h2)
	) name37 (
		f_pad,
		\g0_pad ,
		_w57_
	);
	LUT2 #(
		.INIT('h1)
	) name38 (
		_w56_,
		_w57_,
		_w58_
	);
	LUT2 #(
		.INIT('h4)
	) name39 (
		g_pad,
		_w29_,
		_w59_
	);
	LUT2 #(
		.INIT('h1)
	) name40 (
		g_pad,
		h_pad,
		_w60_
	);
	LUT2 #(
		.INIT('h1)
	) name41 (
		_w20_,
		_w60_,
		_w61_
	);
	LUT2 #(
		.INIT('h8)
	) name42 (
		_w29_,
		_w61_,
		_w62_
	);
	LUT2 #(
		.INIT('h1)
	) name43 (
		i_pad,
		_w20_,
		_w63_
	);
	LUT2 #(
		.INIT('h1)
	) name44 (
		_w21_,
		_w63_,
		_w64_
	);
	LUT2 #(
		.INIT('h8)
	) name45 (
		_w29_,
		_w64_,
		_w65_
	);
	LUT2 #(
		.INIT('h2)
	) name46 (
		j_pad,
		_w21_,
		_w66_
	);
	LUT2 #(
		.INIT('h4)
	) name47 (
		_w22_,
		_w29_,
		_w67_
	);
	LUT2 #(
		.INIT('h4)
	) name48 (
		_w66_,
		_w67_,
		_w68_
	);
	LUT2 #(
		.INIT('h8)
	) name49 (
		k_pad,
		_w67_,
		_w69_
	);
	LUT2 #(
		.INIT('h4)
	) name50 (
		_w25_,
		_w29_,
		_w70_
	);
	LUT2 #(
		.INIT('h4)
	) name51 (
		_w69_,
		_w70_,
		_w71_
	);
	assign \a0_pad  = _w31_ ;
	assign \b0_pad  = _w35_ ;
	assign \c0_pad  = _w41_ ;
	assign \d0_pad  = _w47_ ;
	assign \f0_pad  = _w50_ ;
	assign \h0_pad  = _w51_ ;
	assign t_pad = _w54_ ;
	assign u_pad = _w58_ ;
	assign v_pad = _w59_ ;
	assign w_pad = _w62_ ;
	assign x_pad = _w65_ ;
	assign y_pad = _w68_ ;
	assign z_pad = _w71_ ;
endmodule;