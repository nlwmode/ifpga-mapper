module top( dma_ack_o_pad , dma_nd_i_pad , dma_req_i_pad , \u0_csr_r_reg[0]/NET0131  , \u0_int_maska_r_reg[0]/NET0131  , \u0_int_maska_r_reg[10]/NET0131  , \u0_int_maska_r_reg[11]/NET0131  , \u0_int_maska_r_reg[12]/NET0131  , \u0_int_maska_r_reg[13]/NET0131  , \u0_int_maska_r_reg[14]/NET0131  , \u0_int_maska_r_reg[15]/NET0131  , \u0_int_maska_r_reg[16]/NET0131  , \u0_int_maska_r_reg[17]/NET0131  , \u0_int_maska_r_reg[18]/NET0131  , \u0_int_maska_r_reg[19]/NET0131  , \u0_int_maska_r_reg[1]/NET0131  , \u0_int_maska_r_reg[20]/NET0131  , \u0_int_maska_r_reg[21]/NET0131  , \u0_int_maska_r_reg[22]/NET0131  , \u0_int_maska_r_reg[23]/NET0131  , \u0_int_maska_r_reg[24]/NET0131  , \u0_int_maska_r_reg[25]/NET0131  , \u0_int_maska_r_reg[26]/NET0131  , \u0_int_maska_r_reg[27]/NET0131  , \u0_int_maska_r_reg[28]/NET0131  , \u0_int_maska_r_reg[29]/NET0131  , \u0_int_maska_r_reg[2]/NET0131  , \u0_int_maska_r_reg[30]/NET0131  , \u0_int_maska_r_reg[3]/NET0131  , \u0_int_maska_r_reg[4]/NET0131  , \u0_int_maska_r_reg[5]/NET0131  , \u0_int_maska_r_reg[6]/NET0131  , \u0_int_maska_r_reg[7]/NET0131  , \u0_int_maska_r_reg[8]/NET0131  , \u0_int_maska_r_reg[9]/NET0131  , \u0_int_maskb_r_reg[0]/NET0131  , \u0_int_maskb_r_reg[10]/NET0131  , \u0_int_maskb_r_reg[11]/NET0131  , \u0_int_maskb_r_reg[12]/NET0131  , \u0_int_maskb_r_reg[13]/NET0131  , \u0_int_maskb_r_reg[14]/NET0131  , \u0_int_maskb_r_reg[15]/NET0131  , \u0_int_maskb_r_reg[16]/NET0131  , \u0_int_maskb_r_reg[17]/NET0131  , \u0_int_maskb_r_reg[18]/NET0131  , \u0_int_maskb_r_reg[19]/NET0131  , \u0_int_maskb_r_reg[1]/NET0131  , \u0_int_maskb_r_reg[20]/NET0131  , \u0_int_maskb_r_reg[21]/NET0131  , \u0_int_maskb_r_reg[22]/NET0131  , \u0_int_maskb_r_reg[23]/NET0131  , \u0_int_maskb_r_reg[24]/NET0131  , \u0_int_maskb_r_reg[25]/NET0131  , \u0_int_maskb_r_reg[26]/NET0131  , \u0_int_maskb_r_reg[27]/NET0131  , \u0_int_maskb_r_reg[28]/NET0131  , \u0_int_maskb_r_reg[29]/NET0131  , \u0_int_maskb_r_reg[2]/NET0131  , \u0_int_maskb_r_reg[30]/NET0131  , \u0_int_maskb_r_reg[3]/NET0131  , \u0_int_maskb_r_reg[4]/NET0131  , \u0_int_maskb_r_reg[5]/NET0131  , \u0_int_maskb_r_reg[6]/NET0131  , \u0_int_maskb_r_reg[7]/NET0131  , \u0_int_maskb_r_reg[8]/NET0131  , \u0_int_maskb_r_reg[9]/NET0131  , \u0_u0_ch_adr0_r_reg[0]/P0001  , \u0_u0_ch_adr0_r_reg[10]/P0001  , \u0_u0_ch_adr0_r_reg[11]/P0001  , \u0_u0_ch_adr0_r_reg[12]/P0001  , \u0_u0_ch_adr0_r_reg[13]/P0001  , \u0_u0_ch_adr0_r_reg[14]/P0001  , \u0_u0_ch_adr0_r_reg[15]/P0001  , \u0_u0_ch_adr0_r_reg[16]/P0001  , \u0_u0_ch_adr0_r_reg[17]/P0001  , \u0_u0_ch_adr0_r_reg[18]/P0001  , \u0_u0_ch_adr0_r_reg[19]/P0001  , \u0_u0_ch_adr0_r_reg[1]/P0001  , \u0_u0_ch_adr0_r_reg[20]/P0001  , \u0_u0_ch_adr0_r_reg[21]/P0001  , \u0_u0_ch_adr0_r_reg[22]/P0001  , \u0_u0_ch_adr0_r_reg[23]/P0001  , \u0_u0_ch_adr0_r_reg[24]/P0001  , \u0_u0_ch_adr0_r_reg[25]/P0001  , \u0_u0_ch_adr0_r_reg[26]/P0001  , \u0_u0_ch_adr0_r_reg[27]/P0001  , \u0_u0_ch_adr0_r_reg[28]/P0001  , \u0_u0_ch_adr0_r_reg[29]/P0001  , \u0_u0_ch_adr0_r_reg[2]/P0001  , \u0_u0_ch_adr0_r_reg[3]/P0001  , \u0_u0_ch_adr0_r_reg[4]/P0001  , \u0_u0_ch_adr0_r_reg[5]/P0001  , \u0_u0_ch_adr0_r_reg[6]/P0001  , \u0_u0_ch_adr0_r_reg[7]/P0001  , \u0_u0_ch_adr0_r_reg[8]/P0001  , \u0_u0_ch_adr0_r_reg[9]/P0001  , \u0_u0_ch_adr1_r_reg[0]/P0001  , \u0_u0_ch_adr1_r_reg[10]/P0001  , \u0_u0_ch_adr1_r_reg[11]/P0001  , \u0_u0_ch_adr1_r_reg[12]/P0001  , \u0_u0_ch_adr1_r_reg[13]/P0001  , \u0_u0_ch_adr1_r_reg[14]/P0001  , \u0_u0_ch_adr1_r_reg[15]/P0001  , \u0_u0_ch_adr1_r_reg[16]/P0001  , \u0_u0_ch_adr1_r_reg[17]/P0001  , \u0_u0_ch_adr1_r_reg[18]/P0001  , \u0_u0_ch_adr1_r_reg[19]/P0001  , \u0_u0_ch_adr1_r_reg[1]/P0001  , \u0_u0_ch_adr1_r_reg[20]/P0001  , \u0_u0_ch_adr1_r_reg[21]/P0001  , \u0_u0_ch_adr1_r_reg[22]/P0001  , \u0_u0_ch_adr1_r_reg[23]/P0001  , \u0_u0_ch_adr1_r_reg[24]/P0001  , \u0_u0_ch_adr1_r_reg[25]/P0001  , \u0_u0_ch_adr1_r_reg[26]/P0001  , \u0_u0_ch_adr1_r_reg[27]/P0001  , \u0_u0_ch_adr1_r_reg[28]/P0001  , \u0_u0_ch_adr1_r_reg[29]/P0001  , \u0_u0_ch_adr1_r_reg[2]/P0001  , \u0_u0_ch_adr1_r_reg[3]/P0001  , \u0_u0_ch_adr1_r_reg[4]/P0001  , \u0_u0_ch_adr1_r_reg[5]/P0001  , \u0_u0_ch_adr1_r_reg[6]/P0001  , \u0_u0_ch_adr1_r_reg[7]/P0001  , \u0_u0_ch_adr1_r_reg[8]/P0001  , \u0_u0_ch_adr1_r_reg[9]/P0001  , \u0_u0_ch_busy_reg/P0001  , \u0_u0_ch_chk_sz_r_reg[0]/P0001  , \u0_u0_ch_chk_sz_r_reg[10]/P0001  , \u0_u0_ch_chk_sz_r_reg[1]/P0001  , \u0_u0_ch_chk_sz_r_reg[2]/P0001  , \u0_u0_ch_chk_sz_r_reg[3]/P0001  , \u0_u0_ch_chk_sz_r_reg[4]/P0001  , \u0_u0_ch_chk_sz_r_reg[5]/P0001  , \u0_u0_ch_chk_sz_r_reg[6]/P0001  , \u0_u0_ch_chk_sz_r_reg[7]/P0001  , \u0_u0_ch_chk_sz_r_reg[8]/P0001  , \u0_u0_ch_chk_sz_r_reg[9]/P0001  , \u0_u0_ch_csr_r2_reg[0]/NET0131  , \u0_u0_ch_csr_r2_reg[1]/NET0131  , \u0_u0_ch_csr_r2_reg[2]/NET0131  , \u0_u0_ch_csr_r3_reg[0]/NET0131  , \u0_u0_ch_csr_r3_reg[1]/NET0131  , \u0_u0_ch_csr_r3_reg[2]/NET0131  , \u0_u0_ch_csr_r_reg[0]/NET0131  , \u0_u0_ch_csr_r_reg[1]/NET0131  , \u0_u0_ch_csr_r_reg[2]/NET0131  , \u0_u0_ch_csr_r_reg[3]/NET0131  , \u0_u0_ch_csr_r_reg[4]/NET0131  , \u0_u0_ch_csr_r_reg[5]/NET0131  , \u0_u0_ch_csr_r_reg[6]/NET0131  , \u0_u0_ch_csr_r_reg[7]/NET0131  , \u0_u0_ch_csr_r_reg[8]/NET0131  , \u0_u0_ch_done_reg/P0002  , \u0_u0_ch_err_reg/NET0131  , \u0_u0_ch_stop_reg/P0001  , \u0_u0_ch_sz_inf_reg/NET0131  , \u0_u0_ch_tot_sz_r_reg[0]/P0001  , \u0_u0_ch_tot_sz_r_reg[10]/P0001  , \u0_u0_ch_tot_sz_r_reg[11]/P0001  , \u0_u0_ch_tot_sz_r_reg[1]/P0001  , \u0_u0_ch_tot_sz_r_reg[2]/P0001  , \u0_u0_ch_tot_sz_r_reg[3]/P0001  , \u0_u0_ch_tot_sz_r_reg[4]/P0001  , \u0_u0_ch_tot_sz_r_reg[5]/P0001  , \u0_u0_ch_tot_sz_r_reg[6]/P0001  , \u0_u0_ch_tot_sz_r_reg[7]/P0001  , \u0_u0_ch_tot_sz_r_reg[8]/P0001  , \u0_u0_ch_tot_sz_r_reg[9]/P0001  , \u0_u0_int_src_r_reg[1]/NET0131  , \u0_u0_int_src_r_reg[2]/NET0131  , \u0_u0_rest_en_reg/NET0131  , \u0_wb_rf_dout_reg[0]/P0001  , \u0_wb_rf_dout_reg[10]/P0001  , \u0_wb_rf_dout_reg[11]/P0001  , \u0_wb_rf_dout_reg[12]/P0001  , \u0_wb_rf_dout_reg[13]/P0001  , \u0_wb_rf_dout_reg[14]/P0001  , \u0_wb_rf_dout_reg[15]/P0001  , \u0_wb_rf_dout_reg[16]/P0001  , \u0_wb_rf_dout_reg[17]/P0001  , \u0_wb_rf_dout_reg[18]/P0001  , \u0_wb_rf_dout_reg[19]/P0001  , \u0_wb_rf_dout_reg[1]/P0001  , \u0_wb_rf_dout_reg[20]/P0001  , \u0_wb_rf_dout_reg[21]/P0001  , \u0_wb_rf_dout_reg[22]/P0001  , \u0_wb_rf_dout_reg[23]/P0001  , \u0_wb_rf_dout_reg[24]/P0001  , \u0_wb_rf_dout_reg[25]/P0001  , \u0_wb_rf_dout_reg[26]/P0001  , \u0_wb_rf_dout_reg[27]/P0001  , \u0_wb_rf_dout_reg[28]/P0001  , \u0_wb_rf_dout_reg[29]/P0001  , \u0_wb_rf_dout_reg[2]/P0001  , \u0_wb_rf_dout_reg[30]/P0001  , \u0_wb_rf_dout_reg[31]/P0001  , \u0_wb_rf_dout_reg[3]/P0001  , \u0_wb_rf_dout_reg[4]/P0001  , \u0_wb_rf_dout_reg[5]/P0001  , \u0_wb_rf_dout_reg[6]/P0001  , \u0_wb_rf_dout_reg[7]/P0001  , \u0_wb_rf_dout_reg[8]/P0001  , \u0_wb_rf_dout_reg[9]/P0001  , \u1_de_start_r_reg/P0001  , \u1_ndnr_reg[0]/P0001  , \u1_ndr_r_reg[0]/NET0131  , \u1_next_start_reg/P0001  , \u1_req_r_reg[0]/P0001  , \u2_adr0_cnt_reg[0]/P0001  , \u2_adr0_cnt_reg[10]/P0001  , \u2_adr0_cnt_reg[11]/P0001  , \u2_adr0_cnt_reg[12]/P0001  , \u2_adr0_cnt_reg[13]/P0001  , \u2_adr0_cnt_reg[14]/P0001  , \u2_adr0_cnt_reg[15]/P0001  , \u2_adr0_cnt_reg[16]/NET0131  , \u2_adr0_cnt_reg[17]/P0001  , \u2_adr0_cnt_reg[18]/P0001  , \u2_adr0_cnt_reg[19]/P0001  , \u2_adr0_cnt_reg[1]/P0001  , \u2_adr0_cnt_reg[20]/P0001  , \u2_adr0_cnt_reg[21]/P0001  , \u2_adr0_cnt_reg[22]/P0001  , \u2_adr0_cnt_reg[23]/P0001  , \u2_adr0_cnt_reg[24]/P0001  , \u2_adr0_cnt_reg[25]/P0001  , \u2_adr0_cnt_reg[26]/P0001  , \u2_adr0_cnt_reg[27]/P0001  , \u2_adr0_cnt_reg[28]/P0001  , \u2_adr0_cnt_reg[29]/P0001  , \u2_adr0_cnt_reg[2]/P0001  , \u2_adr0_cnt_reg[3]/P0001  , \u2_adr0_cnt_reg[4]/P0001  , \u2_adr0_cnt_reg[5]/P0001  , \u2_adr0_cnt_reg[6]/P0001  , \u2_adr0_cnt_reg[7]/P0001  , \u2_adr0_cnt_reg[8]/P0001  , \u2_adr0_cnt_reg[9]/P0001  , \u2_adr1_cnt_reg[0]/P0001  , \u2_adr1_cnt_reg[10]/P0001  , \u2_adr1_cnt_reg[11]/P0001  , \u2_adr1_cnt_reg[12]/P0001  , \u2_adr1_cnt_reg[13]/P0001  , \u2_adr1_cnt_reg[14]/P0001  , \u2_adr1_cnt_reg[15]/P0001  , \u2_adr1_cnt_reg[16]/NET0131  , \u2_adr1_cnt_reg[17]/P0001  , \u2_adr1_cnt_reg[18]/P0001  , \u2_adr1_cnt_reg[19]/P0001  , \u2_adr1_cnt_reg[1]/P0001  , \u2_adr1_cnt_reg[20]/P0001  , \u2_adr1_cnt_reg[21]/P0001  , \u2_adr1_cnt_reg[22]/P0001  , \u2_adr1_cnt_reg[23]/P0001  , \u2_adr1_cnt_reg[24]/P0001  , \u2_adr1_cnt_reg[25]/P0001  , \u2_adr1_cnt_reg[26]/P0001  , \u2_adr1_cnt_reg[27]/P0001  , \u2_adr1_cnt_reg[28]/P0001  , \u2_adr1_cnt_reg[29]/P0001  , \u2_adr1_cnt_reg[2]/P0001  , \u2_adr1_cnt_reg[3]/P0001  , \u2_adr1_cnt_reg[4]/P0001  , \u2_adr1_cnt_reg[5]/P0001  , \u2_adr1_cnt_reg[6]/P0001  , \u2_adr1_cnt_reg[7]/P0001  , \u2_adr1_cnt_reg[8]/P0001  , \u2_adr1_cnt_reg[9]/P0001  , \u2_chunk_0_reg/P0001  , \u2_chunk_cnt_is_0_r_reg/P0001  , \u2_chunk_cnt_reg[0]/NET0131  , \u2_chunk_cnt_reg[1]/NET0131  , \u2_chunk_cnt_reg[2]/NET0131  , \u2_chunk_cnt_reg[3]/NET0131  , \u2_chunk_cnt_reg[4]/NET0131  , \u2_chunk_cnt_reg[5]/NET0131  , \u2_chunk_cnt_reg[6]/NET0131  , \u2_chunk_cnt_reg[7]/NET0131  , \u2_chunk_cnt_reg[8]/NET0131  , \u2_chunk_dec_reg/P0001  , \u2_dma_abort_r_reg/NET0131  , \u2_mast0_adr_reg[10]/P0001  , \u2_mast0_adr_reg[11]/P0001  , \u2_mast0_adr_reg[12]/P0001  , \u2_mast0_adr_reg[13]/P0001  , \u2_mast0_adr_reg[14]/P0001  , \u2_mast0_adr_reg[15]/P0001  , \u2_mast0_adr_reg[16]/P0001  , \u2_mast0_adr_reg[17]/P0001  , \u2_mast0_adr_reg[18]/P0001  , \u2_mast0_adr_reg[19]/P0001  , \u2_mast0_adr_reg[20]/P0001  , \u2_mast0_adr_reg[21]/P0001  , \u2_mast0_adr_reg[22]/P0001  , \u2_mast0_adr_reg[23]/P0001  , \u2_mast0_adr_reg[24]/P0001  , \u2_mast0_adr_reg[25]/P0001  , \u2_mast0_adr_reg[26]/P0001  , \u2_mast0_adr_reg[27]/P0001  , \u2_mast0_adr_reg[28]/P0001  , \u2_mast0_adr_reg[29]/P0001  , \u2_mast0_adr_reg[2]/P0001  , \u2_mast0_adr_reg[30]/P0001  , \u2_mast0_adr_reg[31]/P0001  , \u2_mast0_adr_reg[3]/NET0131  , \u2_mast0_adr_reg[4]/P0001  , \u2_mast0_adr_reg[5]/P0001  , \u2_mast0_adr_reg[6]/P0001  , \u2_mast0_adr_reg[7]/P0001  , \u2_mast0_adr_reg[8]/P0001  , \u2_mast0_adr_reg[9]/P0001  , \u2_mast0_drdy_r_reg/P0001  , \u2_mast1_adr_reg[10]/P0001  , \u2_mast1_adr_reg[11]/P0001  , \u2_mast1_adr_reg[12]/P0001  , \u2_mast1_adr_reg[13]/P0001  , \u2_mast1_adr_reg[14]/P0001  , \u2_mast1_adr_reg[15]/P0001  , \u2_mast1_adr_reg[16]/P0001  , \u2_mast1_adr_reg[17]/P0001  , \u2_mast1_adr_reg[18]/P0001  , \u2_mast1_adr_reg[19]/P0001  , \u2_mast1_adr_reg[20]/P0001  , \u2_mast1_adr_reg[21]/P0001  , \u2_mast1_adr_reg[22]/P0001  , \u2_mast1_adr_reg[23]/P0001  , \u2_mast1_adr_reg[24]/P0001  , \u2_mast1_adr_reg[25]/P0001  , \u2_mast1_adr_reg[26]/P0001  , \u2_mast1_adr_reg[27]/P0001  , \u2_mast1_adr_reg[28]/P0001  , \u2_mast1_adr_reg[29]/P0001  , \u2_mast1_adr_reg[2]/P0001  , \u2_mast1_adr_reg[30]/P0001  , \u2_mast1_adr_reg[31]/P0001  , \u2_mast1_adr_reg[3]/P0001  , \u2_mast1_adr_reg[4]/P0001  , \u2_mast1_adr_reg[5]/P0001  , \u2_mast1_adr_reg[6]/P0001  , \u2_mast1_adr_reg[7]/P0001  , \u2_mast1_adr_reg[8]/P0001  , \u2_mast1_adr_reg[9]/P0001  , \u2_next_ch_reg/P0001  , \u2_read_r_reg/P0001  , \u2_state_reg[0]/NET0131  , \u2_state_reg[10]/NET0131  , \u2_state_reg[1]/NET0131  , \u2_state_reg[2]/NET0131  , \u2_state_reg[3]/NET0131  , \u2_state_reg[4]/NET0131  , \u2_state_reg[5]/NET0131  , \u2_state_reg[6]/NET0131  , \u2_state_reg[7]/NET0131  , \u2_state_reg[8]/NET0131  , \u2_state_reg[9]/NET0131  , \u2_tsz_cnt_is_0_r_reg/P0001  , \u2_tsz_cnt_reg[0]/NET0131  , \u2_tsz_cnt_reg[10]/NET0131  , \u2_tsz_cnt_reg[11]/NET0131  , \u2_tsz_cnt_reg[1]/NET0131  , \u2_tsz_cnt_reg[2]/NET0131  , \u2_tsz_cnt_reg[3]/NET0131  , \u2_tsz_cnt_reg[4]/NET0131  , \u2_tsz_cnt_reg[5]/NET0131  , \u2_tsz_cnt_reg[6]/NET0131  , \u2_tsz_cnt_reg[7]/NET0131  , \u2_tsz_cnt_reg[8]/NET0131  , \u2_tsz_cnt_reg[9]/NET0131  , \u2_u0_out_r_reg[0]/P0001  , \u2_u0_out_r_reg[10]/P0001  , \u2_u0_out_r_reg[11]/P0001  , \u2_u0_out_r_reg[12]/P0001  , \u2_u0_out_r_reg[13]/P0001  , \u2_u0_out_r_reg[14]/P0001  , \u2_u0_out_r_reg[15]/P0001  , \u2_u0_out_r_reg[16]/P0001  , \u2_u0_out_r_reg[1]/P0001  , \u2_u0_out_r_reg[2]/P0001  , \u2_u0_out_r_reg[3]/P0001  , \u2_u0_out_r_reg[4]/P0001  , \u2_u0_out_r_reg[5]/P0001  , \u2_u0_out_r_reg[6]/P0001  , \u2_u0_out_r_reg[7]/P0001  , \u2_u0_out_r_reg[8]/P0001  , \u2_u0_out_r_reg[9]/P0001  , \u2_u1_out_r_reg[0]/P0001  , \u2_u1_out_r_reg[10]/P0001  , \u2_u1_out_r_reg[11]/P0001  , \u2_u1_out_r_reg[12]/P0001  , \u2_u1_out_r_reg[13]/P0001  , \u2_u1_out_r_reg[14]/P0001  , \u2_u1_out_r_reg[15]/P0001  , \u2_u1_out_r_reg[16]/P0001  , \u2_u1_out_r_reg[1]/P0001  , \u2_u1_out_r_reg[2]/P0001  , \u2_u1_out_r_reg[3]/P0001  , \u2_u1_out_r_reg[4]/P0001  , \u2_u1_out_r_reg[5]/P0001  , \u2_u1_out_r_reg[6]/P0001  , \u2_u1_out_r_reg[7]/P0001  , \u2_u1_out_r_reg[8]/P0001  , \u2_u1_out_r_reg[9]/P0001  , \u2_write_hold_r_reg/P0001  , \u2_write_r_reg/P0001  , \u3_u0_mast_cyc_reg/P0001  , \u3_u0_mast_dout_reg[0]/P0001  , \u3_u0_mast_dout_reg[10]/P0001  , \u3_u0_mast_dout_reg[11]/P0001  , \u3_u0_mast_dout_reg[12]/P0001  , \u3_u0_mast_dout_reg[13]/P0001  , \u3_u0_mast_dout_reg[14]/P0001  , \u3_u0_mast_dout_reg[15]/P0001  , \u3_u0_mast_dout_reg[16]/P0001  , \u3_u0_mast_dout_reg[17]/P0001  , \u3_u0_mast_dout_reg[18]/P0001  , \u3_u0_mast_dout_reg[19]/P0001  , \u3_u0_mast_dout_reg[1]/P0001  , \u3_u0_mast_dout_reg[20]/P0001  , \u3_u0_mast_dout_reg[21]/P0001  , \u3_u0_mast_dout_reg[22]/P0001  , \u3_u0_mast_dout_reg[23]/P0001  , \u3_u0_mast_dout_reg[24]/P0001  , \u3_u0_mast_dout_reg[25]/P0001  , \u3_u0_mast_dout_reg[26]/P0001  , \u3_u0_mast_dout_reg[27]/P0001  , \u3_u0_mast_dout_reg[28]/P0001  , \u3_u0_mast_dout_reg[29]/P0001  , \u3_u0_mast_dout_reg[2]/P0001  , \u3_u0_mast_dout_reg[30]/P0001  , \u3_u0_mast_dout_reg[31]/P0001  , \u3_u0_mast_dout_reg[3]/P0001  , \u3_u0_mast_dout_reg[4]/P0001  , \u3_u0_mast_dout_reg[5]/P0001  , \u3_u0_mast_dout_reg[6]/P0001  , \u3_u0_mast_dout_reg[7]/P0001  , \u3_u0_mast_dout_reg[8]/P0001  , \u3_u0_mast_dout_reg[9]/P0001  , \u3_u0_mast_stb_reg/P0001  , \u3_u0_mast_we_r_reg/P0002  , \u3_u1_rf_ack_reg/P0001  , \u3_u1_slv_adr_reg[2]/NET0131  , \u3_u1_slv_adr_reg[3]/P0001  , \u3_u1_slv_adr_reg[4]/NET0131  , \u3_u1_slv_adr_reg[5]/P0001  , \u3_u1_slv_adr_reg[6]/NET0131  , \u3_u1_slv_adr_reg[7]/NET0131  , \u3_u1_slv_adr_reg[8]/NET0131  , \u3_u1_slv_adr_reg[9]/NET0131  , \u3_u1_slv_dout_reg[0]/P0001  , \u3_u1_slv_dout_reg[10]/P0001  , \u3_u1_slv_dout_reg[11]/P0001  , \u3_u1_slv_dout_reg[12]/P0001  , \u3_u1_slv_dout_reg[13]/P0001  , \u3_u1_slv_dout_reg[14]/P0001  , \u3_u1_slv_dout_reg[15]/P0001  , \u3_u1_slv_dout_reg[16]/P0001  , \u3_u1_slv_dout_reg[17]/P0001  , \u3_u1_slv_dout_reg[18]/P0001  , \u3_u1_slv_dout_reg[19]/P0001  , \u3_u1_slv_dout_reg[1]/P0001  , \u3_u1_slv_dout_reg[20]/P0001  , \u3_u1_slv_dout_reg[21]/P0001  , \u3_u1_slv_dout_reg[22]/P0001  , \u3_u1_slv_dout_reg[23]/P0001  , \u3_u1_slv_dout_reg[24]/P0001  , \u3_u1_slv_dout_reg[25]/P0001  , \u3_u1_slv_dout_reg[26]/P0001  , \u3_u1_slv_dout_reg[27]/P0001  , \u3_u1_slv_dout_reg[28]/P0001  , \u3_u1_slv_dout_reg[29]/P0001  , \u3_u1_slv_dout_reg[2]/P0001  , \u3_u1_slv_dout_reg[30]/P0001  , \u3_u1_slv_dout_reg[31]/P0001  , \u3_u1_slv_dout_reg[3]/P0001  , \u3_u1_slv_dout_reg[4]/P0001  , \u3_u1_slv_dout_reg[5]/P0001  , \u3_u1_slv_dout_reg[6]/P0001  , \u3_u1_slv_dout_reg[7]/P0001  , \u3_u1_slv_dout_reg[8]/P0001  , \u3_u1_slv_dout_reg[9]/P0001  , \u3_u1_slv_re_reg/P0001  , \u3_u1_slv_we_reg/P0001  , \u4_u0_mast_cyc_reg/P0001  , \u4_u0_mast_dout_reg[0]/P0001  , \u4_u0_mast_dout_reg[10]/P0001  , \u4_u0_mast_dout_reg[11]/P0001  , \u4_u0_mast_dout_reg[12]/P0001  , \u4_u0_mast_dout_reg[13]/P0001  , \u4_u0_mast_dout_reg[14]/P0001  , \u4_u0_mast_dout_reg[15]/P0001  , \u4_u0_mast_dout_reg[16]/P0001  , \u4_u0_mast_dout_reg[17]/P0001  , \u4_u0_mast_dout_reg[18]/P0001  , \u4_u0_mast_dout_reg[19]/P0001  , \u4_u0_mast_dout_reg[1]/P0001  , \u4_u0_mast_dout_reg[20]/P0001  , \u4_u0_mast_dout_reg[21]/P0001  , \u4_u0_mast_dout_reg[22]/P0001  , \u4_u0_mast_dout_reg[23]/P0001  , \u4_u0_mast_dout_reg[24]/P0001  , \u4_u0_mast_dout_reg[25]/P0001  , \u4_u0_mast_dout_reg[26]/P0001  , \u4_u0_mast_dout_reg[27]/P0001  , \u4_u0_mast_dout_reg[28]/P0001  , \u4_u0_mast_dout_reg[29]/P0001  , \u4_u0_mast_dout_reg[2]/P0001  , \u4_u0_mast_dout_reg[30]/P0001  , \u4_u0_mast_dout_reg[31]/P0001  , \u4_u0_mast_dout_reg[3]/P0001  , \u4_u0_mast_dout_reg[4]/P0001  , \u4_u0_mast_dout_reg[5]/P0001  , \u4_u0_mast_dout_reg[6]/P0001  , \u4_u0_mast_dout_reg[7]/P0001  , \u4_u0_mast_dout_reg[8]/P0001  , \u4_u0_mast_dout_reg[9]/P0001  , \u4_u0_mast_stb_reg/P0001  , \u4_u0_mast_we_r_reg/P0001  , \u4_u1_rf_ack_reg/P0001  , \u4_u1_slv_re_reg/P0001  , \u4_u1_slv_we_reg/P0001  , \wb0_ack_i_pad  , \wb0_addr_i[0]_pad  , \wb0_addr_i[10]_pad  , \wb0_addr_i[11]_pad  , \wb0_addr_i[12]_pad  , \wb0_addr_i[13]_pad  , \wb0_addr_i[14]_pad  , \wb0_addr_i[15]_pad  , \wb0_addr_i[16]_pad  , \wb0_addr_i[17]_pad  , \wb0_addr_i[18]_pad  , \wb0_addr_i[19]_pad  , \wb0_addr_i[1]_pad  , \wb0_addr_i[20]_pad  , \wb0_addr_i[21]_pad  , \wb0_addr_i[22]_pad  , \wb0_addr_i[23]_pad  , \wb0_addr_i[24]_pad  , \wb0_addr_i[25]_pad  , \wb0_addr_i[26]_pad  , \wb0_addr_i[27]_pad  , \wb0_addr_i[28]_pad  , \wb0_addr_i[29]_pad  , \wb0_addr_i[2]_pad  , \wb0_addr_i[30]_pad  , \wb0_addr_i[31]_pad  , \wb0_addr_i[3]_pad  , \wb0_addr_i[4]_pad  , \wb0_addr_i[5]_pad  , \wb0_addr_i[6]_pad  , \wb0_addr_i[7]_pad  , \wb0_addr_i[8]_pad  , \wb0_addr_i[9]_pad  , \wb0_cyc_i_pad  , \wb0_err_i_pad  , \wb0_rty_i_pad  , \wb0_sel_i[0]_pad  , \wb0_sel_i[1]_pad  , \wb0_sel_i[2]_pad  , \wb0_sel_i[3]_pad  , \wb0_stb_i_pad  , \wb0_we_i_pad  , \wb0m_data_i[0]_pad  , \wb0m_data_i[10]_pad  , \wb0m_data_i[11]_pad  , \wb0m_data_i[12]_pad  , \wb0m_data_i[13]_pad  , \wb0m_data_i[14]_pad  , \wb0m_data_i[15]_pad  , \wb0m_data_i[16]_pad  , \wb0m_data_i[17]_pad  , \wb0m_data_i[18]_pad  , \wb0m_data_i[19]_pad  , \wb0m_data_i[1]_pad  , \wb0m_data_i[20]_pad  , \wb0m_data_i[21]_pad  , \wb0m_data_i[22]_pad  , \wb0m_data_i[23]_pad  , \wb0m_data_i[24]_pad  , \wb0m_data_i[25]_pad  , \wb0m_data_i[26]_pad  , \wb0m_data_i[27]_pad  , \wb0m_data_i[28]_pad  , \wb0m_data_i[29]_pad  , \wb0m_data_i[2]_pad  , \wb0m_data_i[30]_pad  , \wb0m_data_i[31]_pad  , \wb0m_data_i[3]_pad  , \wb0m_data_i[4]_pad  , \wb0m_data_i[5]_pad  , \wb0m_data_i[6]_pad  , \wb0m_data_i[7]_pad  , \wb0m_data_i[8]_pad  , \wb0m_data_i[9]_pad  , \wb0s_data_i[0]_pad  , \wb0s_data_i[10]_pad  , \wb0s_data_i[11]_pad  , \wb0s_data_i[12]_pad  , \wb0s_data_i[13]_pad  , \wb0s_data_i[14]_pad  , \wb0s_data_i[15]_pad  , \wb0s_data_i[16]_pad  , \wb0s_data_i[17]_pad  , \wb0s_data_i[18]_pad  , \wb0s_data_i[19]_pad  , \wb0s_data_i[1]_pad  , \wb0s_data_i[20]_pad  , \wb0s_data_i[21]_pad  , \wb0s_data_i[22]_pad  , \wb0s_data_i[23]_pad  , \wb0s_data_i[24]_pad  , \wb0s_data_i[25]_pad  , \wb0s_data_i[26]_pad  , \wb0s_data_i[27]_pad  , \wb0s_data_i[28]_pad  , \wb0s_data_i[29]_pad  , \wb0s_data_i[2]_pad  , \wb0s_data_i[30]_pad  , \wb0s_data_i[31]_pad  , \wb0s_data_i[3]_pad  , \wb0s_data_i[4]_pad  , \wb0s_data_i[5]_pad  , \wb0s_data_i[6]_pad  , \wb0s_data_i[7]_pad  , \wb0s_data_i[8]_pad  , \wb0s_data_i[9]_pad  , \wb1_ack_i_pad  , \wb1_addr_i[0]_pad  , \wb1_addr_i[10]_pad  , \wb1_addr_i[11]_pad  , \wb1_addr_i[12]_pad  , \wb1_addr_i[13]_pad  , \wb1_addr_i[14]_pad  , \wb1_addr_i[15]_pad  , \wb1_addr_i[16]_pad  , \wb1_addr_i[17]_pad  , \wb1_addr_i[18]_pad  , \wb1_addr_i[19]_pad  , \wb1_addr_i[1]_pad  , \wb1_addr_i[20]_pad  , \wb1_addr_i[21]_pad  , \wb1_addr_i[22]_pad  , \wb1_addr_i[23]_pad  , \wb1_addr_i[24]_pad  , \wb1_addr_i[25]_pad  , \wb1_addr_i[26]_pad  , \wb1_addr_i[27]_pad  , \wb1_addr_i[28]_pad  , \wb1_addr_i[29]_pad  , \wb1_addr_i[2]_pad  , \wb1_addr_i[30]_pad  , \wb1_addr_i[31]_pad  , \wb1_addr_i[3]_pad  , \wb1_addr_i[4]_pad  , \wb1_addr_i[5]_pad  , \wb1_addr_i[6]_pad  , \wb1_addr_i[7]_pad  , \wb1_addr_i[8]_pad  , \wb1_addr_i[9]_pad  , \wb1_cyc_i_pad  , \wb1_err_i_pad  , \wb1_rty_i_pad  , \wb1_sel_i[0]_pad  , \wb1_sel_i[1]_pad  , \wb1_sel_i[2]_pad  , \wb1_sel_i[3]_pad  , \wb1_stb_i_pad  , \wb1_we_i_pad  , \wb1m_data_i[0]_pad  , \wb1m_data_i[10]_pad  , \wb1m_data_i[11]_pad  , \wb1m_data_i[12]_pad  , \wb1m_data_i[13]_pad  , \wb1m_data_i[14]_pad  , \wb1m_data_i[15]_pad  , \wb1m_data_i[16]_pad  , \wb1m_data_i[17]_pad  , \wb1m_data_i[18]_pad  , \wb1m_data_i[19]_pad  , \wb1m_data_i[1]_pad  , \wb1m_data_i[20]_pad  , \wb1m_data_i[21]_pad  , \wb1m_data_i[22]_pad  , \wb1m_data_i[23]_pad  , \wb1m_data_i[24]_pad  , \wb1m_data_i[25]_pad  , \wb1m_data_i[26]_pad  , \wb1m_data_i[27]_pad  , \wb1m_data_i[28]_pad  , \wb1m_data_i[29]_pad  , \wb1m_data_i[2]_pad  , \wb1m_data_i[30]_pad  , \wb1m_data_i[31]_pad  , \wb1m_data_i[3]_pad  , \wb1m_data_i[4]_pad  , \wb1m_data_i[5]_pad  , \wb1m_data_i[6]_pad  , \wb1m_data_i[7]_pad  , \wb1m_data_i[8]_pad  , \wb1m_data_i[9]_pad  , \wb1s_data_i[0]_pad  , \wb1s_data_i[10]_pad  , \wb1s_data_i[11]_pad  , \wb1s_data_i[12]_pad  , \wb1s_data_i[13]_pad  , \wb1s_data_i[14]_pad  , \wb1s_data_i[15]_pad  , \wb1s_data_i[16]_pad  , \wb1s_data_i[17]_pad  , \wb1s_data_i[18]_pad  , \wb1s_data_i[19]_pad  , \wb1s_data_i[1]_pad  , \wb1s_data_i[20]_pad  , \wb1s_data_i[21]_pad  , \wb1s_data_i[22]_pad  , \wb1s_data_i[23]_pad  , \wb1s_data_i[24]_pad  , \wb1s_data_i[25]_pad  , \wb1s_data_i[26]_pad  , \wb1s_data_i[27]_pad  , \wb1s_data_i[28]_pad  , \wb1s_data_i[29]_pad  , \wb1s_data_i[2]_pad  , \wb1s_data_i[30]_pad  , \wb1s_data_i[31]_pad  , \wb1s_data_i[3]_pad  , \wb1s_data_i[4]_pad  , \wb1s_data_i[5]_pad  , \wb1s_data_i[6]_pad  , \wb1s_data_i[7]_pad  , \wb1s_data_i[8]_pad  , \wb1s_data_i[9]_pad  , \_al_n0  , \_al_n1  , \g22594/_0_  , \g22595/_0_  , \g22599/_0_  , \g22600/_0_  , \g22606/_0_  , \g22607/_0_  , \g22610/_0_  , \g22614/_0_  , \g22615/_0_  , \g22616/_0_  , \g22619/_0_  , \g22620/_0_  , \g22626/_0_  , \g22635/_0_  , \g22650/_0_  , \g22651/_0_  , \g22692/_0_  , \g22727/_0_  , \g22729/_3_  , \g22774/_0_  , \g22775/_0_  , \g22776/_0_  , \g22777/_0_  , \g22779/_3_  , \g22780/_0_  , \g22781/_0_  , \g22782/_0_  , \g22784/_0_  , \g22785/_0_  , \g22786/_0_  , \g22787/_0_  , \g22789/_3_  , \g22790/_0_  , \g22791/_0_  , \g22792/_0_  , \g22793/_0_  , \g22794/_0_  , \g22795/_0_  , \g22796/_0_  , \g22797/_0_  , \g22798/_0_  , \g22799/_0_  , \g22838/_0_  , \g22839/_0_  , \g22841/_0_  , \g22842/_0_  , \g22847/_0_  , \g22848/_0_  , \g22849/_0_  , \g22850/_0_  , \g22851/_0_  , \g22852/_0_  , \g22853/_0_  , \g22854/_0_  , \g22855/_0_  , \g22856/_0_  , \g22857/_0_  , \g22858/_0_  , \g22859/_0_  , \g22860/_0_  , \g22861/_0_  , \g22862/_0_  , \g22863/_0_  , \g22864/_0_  , \g22865/_0_  , \g22867/_0_  , \g22868/_0_  , \g22869/_0_  , \g22871/_0_  , \g22872/_0_  , \g22873/_0_  , \g22874/_0_  , \g22875/_0_  , \g22876/_0_  , \g22878/_0_  , \g22882/_2_  , \g22995/_0_  , \g23030/_0_  , \g23046/_0_  , \g23077/_0_  , \g23111/_0_  , \g23115/_1_  , \g23124/_2_  , \g23126/_2_  , \g23128/_2_  , \g23130/_2_  , \g23132/_2_  , \g23134/_2_  , \g23136/_2_  , \g23137/_0_  , \g23140/_2_  , \g23142/_2_  , \g23144/_2_  , \g23146/_2_  , \g23148/_2_  , \g23150/_2_  , \g23152/_2_  , \g23154/_2_  , \g23156/_2_  , \g23158/_2_  , \g23160/_2_  , \g23162/_2_  , \g23163/_3_  , \g23164/_0_  , \g23166/_0_  , \g23168/_0_  , \g23170/_2_  , \g23172/_2_  , \g23174/_2_  , \g23175/_0_  , \g23177/_0_  , \g23180/_2_  , \g23220/_0_  , \g23238/_0_  , \g23239/_0_  , \g23240/_0_  , \g23241/_0_  , \g23242/_0_  , \g23243/_0_  , \g23244/_0_  , \g23245/_0_  , \g23247/_3_  , \g23248/_0_  , \g23249/_0_  , \g23250/_0_  , \g23251/_0_  , \g23252/_0_  , \g23253/_0_  , \g23255/_3_  , \g23260/_0_  , \g23284/_3_  , \g23285/_0_  , \g23334/_0_  , \g23343/_0_  , \g23366/_0_  , \g23402/_0_  , \g23403/_0_  , \g23404/_0_  , \g23405/_0_  , \g23407/_0_  , \g23408/_0_  , \g23409/_0_  , \g23410/_0_  , \g23411/_0_  , \g23413/_2_  , \g23415/_2_  , \g23417/_2_  , \g23542/_0_  , \g23607/_0_  , \g23608/_0_  , \g23609/_3_  , \g23707/_0_  , \g23708/_0_  , \g23709/_0_  , \g23710/_0_  , \g23711/_0_  , \g23712/_0_  , \g23713/_0_  , \g23714/_0_  , \g23715/_0_  , \g23716/_0_  , \g23754/_0_  , \g23755/_0_  , \g23756/_0_  , \g23757/_0_  , \g23758/_0_  , \g23759/_0_  , \g23760/_0_  , \g23761/_0_  , \g23763/_3_  , \g23767/_0_  , \g23768/_0_  , \g23833/_0_  , \g23837/_0_  , \g23838/_0_  , \g23839/_0_  , \g23840/_0_  , \g23841/_0_  , \g23842/_0_  , \g23843/_0_  , \g23844/_0_  , \g23845/_0_  , \g23849/_3_  , \g23851/_3_  , \g23858/_0_  , \g23870/_0_  , \g23871/_0_  , \g23872/_3_  , \g23873/_3_  , \g23874/_3_  , \g23875/_3_  , \g23876/_3_  , \g23877/_3_  , \g23878/_3_  , \g23879/_3_  , \g23880/_3_  , \g23881/_3_  , \g23882/_3_  , \g23883/_3_  , \g23884/_3_  , \g23885/_3_  , \g23886/_3_  , \g23887/_3_  , \g23888/_3_  , \g23889/_3_  , \g23890/_3_  , \g23891/_3_  , \g23892/_3_  , \g23893/_3_  , \g23894/_3_  , \g23895/_3_  , \g23896/_3_  , \g23897/_3_  , \g23898/_3_  , \g23899/_3_  , \g23900/_3_  , \g23901/_3_  , \g23902/_3_  , \g23903/_3_  , \g23904/_3_  , \g23905/_3_  , \g23906/_3_  , \g23907/_3_  , \g23908/_3_  , \g23909/_3_  , \g23910/_3_  , \g23911/_3_  , \g23912/_3_  , \g23913/_3_  , \g23914/_3_  , \g23915/_3_  , \g23959/_0_  , \g23961/_0_  , \g23962/_0_  , \g23966/_0_  , \g23967/_0_  , \g23969/_0_  , \g23970/_0_  , \g23971/_0_  , \g23972/_0_  , \g23979/_0_  , \g23987/_0_  , \g23988/_0_  , \g23989/_0_  , \g23990/_0_  , \g24005/_0_  , \g24010/_0_  , \g24012/_0_  , \g24013/_0_  , \g24014/_0_  , \g24015/_0_  , \g24016/_0_  , \g24017/_0_  , \g24018/_0_  , \g24019/_0_  , \g24020/_0_  , \g24026/_0_  , \g24027/_0_  , \g24028/_0_  , \g24029/_0_  , \g24030/_0_  , \g24031/_0_  , \g24032/_0_  , \g24033/_0_  , \g24034/_0_  , \g24035/_0_  , \g24036/_0_  , \g24037/_0_  , \g24038/_0_  , \g24039/_0_  , \g24042/_0_  , \g24049/_0_  , \g24063/_0_  , \g24119/_0_  , \g24120/_0_  , \g24357/_0_  , \g24432/_0_  , \g24433/_0_  , \g24437/_0_  , \g24438/_0_  , \g24477/_0_  , \g24491/_0_  , \g24530/_2_  , \g24532/_0_  , \g24534/_0_  , \g24537/_0_  , \g24538/_0_  , \g24539/_0_  , \g24540/_0_  , \g24606/_2_  , \g24612/_0_  , \g24677/_0_  , \g24678/_0_  , \g24679/_0_  , \g24688/_0_  , \g24743/_0_  , \g24847/_0_  , \g24849/_0_  , \g24850/_0_  , \g24854/_0_  , \g24862/_0_  , \g24872/_0_  , \g24873/_0_  , \g24874/_0_  , \g24876/_0_  , \g24879/_0_  , \g24880/_0_  , \g24881/_0_  , \g24882/_0_  , \g24952/_2_  , \g24976/_1_  , \g25003/_0_  , \g25004/_0_  , \g25005/_0_  , \g25006/_0_  , \g25011/_0_  , \g25012/_0_  , \g25013/_0_  , \g25031/_0_  , \g25032/_0_  , \g25033/_0_  , \g25034/_0_  , \g25035/_0_  , \g25153/_2_  , \g25183/_0_  , \g25184/_0_  , \g25224/_0_  , \g25232/_0_  , \g25237/_0_  , \g25241/_2_  , \g25243/_2_  , \g25248/_3_  , \g25261/_0_  , \g25262/_0_  , \g25266/_3_  , \g25267/_0_  , \g25269/_0_  , \g25543/_1_  , \g25602/_3_  , \g25610/_0_  , \g25611/_0_  , \g25841/_0_  , \g25843/_0_  , \g25893/_0_  , \g27013/_0_  , \g27060/_0_  , \g27073/_0_  , \g27184/_0_  , \g27186/_0_  , \g27189/_2_  , \g47/_0_  , \u0_u0_ch_done_reg/_05_  , \u2_adr0_cnt_reg[0]/P0000  , \u2_adr1_cnt_reg[0]/P0000  , \u3_u0_mast_we_r_reg/_05_  , \wb0_ack_o_pad  , \wb0_addr_o[0]_pad  , \wb0_addr_o[10]_pad  , \wb0_addr_o[11]_pad  , \wb0_addr_o[12]_pad  , \wb0_addr_o[13]_pad  , \wb0_addr_o[14]_pad  , \wb0_addr_o[15]_pad  , \wb0_addr_o[16]_pad  , \wb0_addr_o[17]_pad  , \wb0_addr_o[18]_pad  , \wb0_addr_o[19]_pad  , \wb0_addr_o[1]_pad  , \wb0_addr_o[20]_pad  , \wb0_addr_o[21]_pad  , \wb0_addr_o[22]_pad  , \wb0_addr_o[23]_pad  , \wb0_addr_o[24]_pad  , \wb0_addr_o[25]_pad  , \wb0_addr_o[26]_pad  , \wb0_addr_o[27]_pad  , \wb0_addr_o[28]_pad  , \wb0_addr_o[29]_pad  , \wb0_addr_o[2]_pad  , \wb0_addr_o[30]_pad  , \wb0_addr_o[31]_pad  , \wb0_addr_o[3]_pad  , \wb0_addr_o[4]_pad  , \wb0_addr_o[5]_pad  , \wb0_addr_o[6]_pad  , \wb0_addr_o[7]_pad  , \wb0_addr_o[8]_pad  , \wb0_addr_o[9]_pad  , \wb0_cyc_o_pad  , \wb0_err_o_pad  , \wb0_rty_o_pad  , \wb0_sel_o[0]_pad  , \wb0_sel_o[1]_pad  , \wb0_sel_o[2]_pad  , \wb0_sel_o[3]_pad  , \wb0_stb_o_pad  , \wb0_we_o_pad  , \wb0m_data_o[0]_pad  , \wb0m_data_o[10]_pad  , \wb0m_data_o[11]_pad  , \wb0m_data_o[12]_pad  , \wb0m_data_o[13]_pad  , \wb0m_data_o[14]_pad  , \wb0m_data_o[15]_pad  , \wb0m_data_o[16]_pad  , \wb0m_data_o[17]_pad  , \wb0m_data_o[18]_pad  , \wb0m_data_o[19]_pad  , \wb0m_data_o[1]_pad  , \wb0m_data_o[20]_pad  , \wb0m_data_o[21]_pad  , \wb0m_data_o[22]_pad  , \wb0m_data_o[23]_pad  , \wb0m_data_o[24]_pad  , \wb0m_data_o[25]_pad  , \wb0m_data_o[26]_pad  , \wb0m_data_o[27]_pad  , \wb0m_data_o[28]_pad  , \wb0m_data_o[29]_pad  , \wb0m_data_o[2]_pad  , \wb0m_data_o[30]_pad  , \wb0m_data_o[31]_pad  , \wb0m_data_o[3]_pad  , \wb0m_data_o[4]_pad  , \wb0m_data_o[5]_pad  , \wb0m_data_o[6]_pad  , \wb0m_data_o[7]_pad  , \wb0m_data_o[8]_pad  , \wb0m_data_o[9]_pad  , \wb0s_data_o[0]_pad  , \wb0s_data_o[10]_pad  , \wb0s_data_o[11]_pad  , \wb0s_data_o[12]_pad  , \wb0s_data_o[13]_pad  , \wb0s_data_o[14]_pad  , \wb0s_data_o[15]_pad  , \wb0s_data_o[16]_pad  , \wb0s_data_o[17]_pad  , \wb0s_data_o[18]_pad  , \wb0s_data_o[19]_pad  , \wb0s_data_o[1]_pad  , \wb0s_data_o[20]_pad  , \wb0s_data_o[21]_pad  , \wb0s_data_o[22]_pad  , \wb0s_data_o[23]_pad  , \wb0s_data_o[24]_pad  , \wb0s_data_o[25]_pad  , \wb0s_data_o[26]_pad  , \wb0s_data_o[27]_pad  , \wb0s_data_o[28]_pad  , \wb0s_data_o[29]_pad  , \wb0s_data_o[2]_pad  , \wb0s_data_o[30]_pad  , \wb0s_data_o[31]_pad  , \wb0s_data_o[3]_pad  , \wb0s_data_o[4]_pad  , \wb0s_data_o[5]_pad  , \wb0s_data_o[6]_pad  , \wb0s_data_o[7]_pad  , \wb0s_data_o[8]_pad  , \wb0s_data_o[9]_pad  , \wb1_ack_o_pad  , \wb1_addr_o[0]_pad  , \wb1_addr_o[10]_pad  , \wb1_addr_o[11]_pad  , \wb1_addr_o[12]_pad  , \wb1_addr_o[13]_pad  , \wb1_addr_o[14]_pad  , \wb1_addr_o[15]_pad  , \wb1_addr_o[16]_pad  , \wb1_addr_o[17]_pad  , \wb1_addr_o[18]_pad  , \wb1_addr_o[19]_pad  , \wb1_addr_o[1]_pad  , \wb1_addr_o[20]_pad  , \wb1_addr_o[21]_pad  , \wb1_addr_o[22]_pad  , \wb1_addr_o[23]_pad  , \wb1_addr_o[24]_pad  , \wb1_addr_o[25]_pad  , \wb1_addr_o[26]_pad  , \wb1_addr_o[27]_pad  , \wb1_addr_o[28]_pad  , \wb1_addr_o[29]_pad  , \wb1_addr_o[2]_pad  , \wb1_addr_o[30]_pad  , \wb1_addr_o[31]_pad  , \wb1_addr_o[3]_pad  , \wb1_addr_o[4]_pad  , \wb1_addr_o[5]_pad  , \wb1_addr_o[6]_pad  , \wb1_addr_o[7]_pad  , \wb1_addr_o[8]_pad  , \wb1_addr_o[9]_pad  , \wb1_cyc_o_pad  , \wb1_err_o_pad  , \wb1_rty_o_pad  , \wb1_sel_o[0]_pad  , \wb1_sel_o[1]_pad  , \wb1_sel_o[2]_pad  , \wb1_sel_o[3]_pad  , \wb1_stb_o_pad  , \wb1_we_o_pad  , \wb1m_data_o[0]_pad  , \wb1m_data_o[10]_pad  , \wb1m_data_o[11]_pad  , \wb1m_data_o[12]_pad  , \wb1m_data_o[13]_pad  , \wb1m_data_o[14]_pad  , \wb1m_data_o[15]_pad  , \wb1m_data_o[16]_pad  , \wb1m_data_o[17]_pad  , \wb1m_data_o[18]_pad  , \wb1m_data_o[19]_pad  , \wb1m_data_o[1]_pad  , \wb1m_data_o[20]_pad  , \wb1m_data_o[21]_pad  , \wb1m_data_o[22]_pad  , \wb1m_data_o[23]_pad  , \wb1m_data_o[24]_pad  , \wb1m_data_o[25]_pad  , \wb1m_data_o[26]_pad  , \wb1m_data_o[27]_pad  , \wb1m_data_o[28]_pad  , \wb1m_data_o[29]_pad  , \wb1m_data_o[2]_pad  , \wb1m_data_o[30]_pad  , \wb1m_data_o[31]_pad  , \wb1m_data_o[3]_pad  , \wb1m_data_o[4]_pad  , \wb1m_data_o[5]_pad  , \wb1m_data_o[6]_pad  , \wb1m_data_o[7]_pad  , \wb1m_data_o[8]_pad  , \wb1m_data_o[9]_pad  , \wb1s_data_o[0]_pad  , \wb1s_data_o[10]_pad  , \wb1s_data_o[11]_pad  , \wb1s_data_o[12]_pad  , \wb1s_data_o[13]_pad  , \wb1s_data_o[14]_pad  , \wb1s_data_o[15]_pad  , \wb1s_data_o[16]_pad  , \wb1s_data_o[17]_pad  , \wb1s_data_o[18]_pad  , \wb1s_data_o[19]_pad  , \wb1s_data_o[1]_pad  , \wb1s_data_o[20]_pad  , \wb1s_data_o[21]_pad  , \wb1s_data_o[22]_pad  , \wb1s_data_o[23]_pad  , \wb1s_data_o[24]_pad  , \wb1s_data_o[25]_pad  , \wb1s_data_o[26]_pad  , \wb1s_data_o[27]_pad  , \wb1s_data_o[28]_pad  , \wb1s_data_o[29]_pad  , \wb1s_data_o[2]_pad  , \wb1s_data_o[30]_pad  , \wb1s_data_o[31]_pad  , \wb1s_data_o[3]_pad  , \wb1s_data_o[4]_pad  , \wb1s_data_o[5]_pad  , \wb1s_data_o[6]_pad  , \wb1s_data_o[7]_pad  , \wb1s_data_o[8]_pad  , \wb1s_data_o[9]_pad  );
  input dma_ack_o_pad ;
  input dma_nd_i_pad ;
  input dma_req_i_pad ;
  input \u0_csr_r_reg[0]/NET0131  ;
  input \u0_int_maska_r_reg[0]/NET0131  ;
  input \u0_int_maska_r_reg[10]/NET0131  ;
  input \u0_int_maska_r_reg[11]/NET0131  ;
  input \u0_int_maska_r_reg[12]/NET0131  ;
  input \u0_int_maska_r_reg[13]/NET0131  ;
  input \u0_int_maska_r_reg[14]/NET0131  ;
  input \u0_int_maska_r_reg[15]/NET0131  ;
  input \u0_int_maska_r_reg[16]/NET0131  ;
  input \u0_int_maska_r_reg[17]/NET0131  ;
  input \u0_int_maska_r_reg[18]/NET0131  ;
  input \u0_int_maska_r_reg[19]/NET0131  ;
  input \u0_int_maska_r_reg[1]/NET0131  ;
  input \u0_int_maska_r_reg[20]/NET0131  ;
  input \u0_int_maska_r_reg[21]/NET0131  ;
  input \u0_int_maska_r_reg[22]/NET0131  ;
  input \u0_int_maska_r_reg[23]/NET0131  ;
  input \u0_int_maska_r_reg[24]/NET0131  ;
  input \u0_int_maska_r_reg[25]/NET0131  ;
  input \u0_int_maska_r_reg[26]/NET0131  ;
  input \u0_int_maska_r_reg[27]/NET0131  ;
  input \u0_int_maska_r_reg[28]/NET0131  ;
  input \u0_int_maska_r_reg[29]/NET0131  ;
  input \u0_int_maska_r_reg[2]/NET0131  ;
  input \u0_int_maska_r_reg[30]/NET0131  ;
  input \u0_int_maska_r_reg[3]/NET0131  ;
  input \u0_int_maska_r_reg[4]/NET0131  ;
  input \u0_int_maska_r_reg[5]/NET0131  ;
  input \u0_int_maska_r_reg[6]/NET0131  ;
  input \u0_int_maska_r_reg[7]/NET0131  ;
  input \u0_int_maska_r_reg[8]/NET0131  ;
  input \u0_int_maska_r_reg[9]/NET0131  ;
  input \u0_int_maskb_r_reg[0]/NET0131  ;
  input \u0_int_maskb_r_reg[10]/NET0131  ;
  input \u0_int_maskb_r_reg[11]/NET0131  ;
  input \u0_int_maskb_r_reg[12]/NET0131  ;
  input \u0_int_maskb_r_reg[13]/NET0131  ;
  input \u0_int_maskb_r_reg[14]/NET0131  ;
  input \u0_int_maskb_r_reg[15]/NET0131  ;
  input \u0_int_maskb_r_reg[16]/NET0131  ;
  input \u0_int_maskb_r_reg[17]/NET0131  ;
  input \u0_int_maskb_r_reg[18]/NET0131  ;
  input \u0_int_maskb_r_reg[19]/NET0131  ;
  input \u0_int_maskb_r_reg[1]/NET0131  ;
  input \u0_int_maskb_r_reg[20]/NET0131  ;
  input \u0_int_maskb_r_reg[21]/NET0131  ;
  input \u0_int_maskb_r_reg[22]/NET0131  ;
  input \u0_int_maskb_r_reg[23]/NET0131  ;
  input \u0_int_maskb_r_reg[24]/NET0131  ;
  input \u0_int_maskb_r_reg[25]/NET0131  ;
  input \u0_int_maskb_r_reg[26]/NET0131  ;
  input \u0_int_maskb_r_reg[27]/NET0131  ;
  input \u0_int_maskb_r_reg[28]/NET0131  ;
  input \u0_int_maskb_r_reg[29]/NET0131  ;
  input \u0_int_maskb_r_reg[2]/NET0131  ;
  input \u0_int_maskb_r_reg[30]/NET0131  ;
  input \u0_int_maskb_r_reg[3]/NET0131  ;
  input \u0_int_maskb_r_reg[4]/NET0131  ;
  input \u0_int_maskb_r_reg[5]/NET0131  ;
  input \u0_int_maskb_r_reg[6]/NET0131  ;
  input \u0_int_maskb_r_reg[7]/NET0131  ;
  input \u0_int_maskb_r_reg[8]/NET0131  ;
  input \u0_int_maskb_r_reg[9]/NET0131  ;
  input \u0_u0_ch_adr0_r_reg[0]/P0001  ;
  input \u0_u0_ch_adr0_r_reg[10]/P0001  ;
  input \u0_u0_ch_adr0_r_reg[11]/P0001  ;
  input \u0_u0_ch_adr0_r_reg[12]/P0001  ;
  input \u0_u0_ch_adr0_r_reg[13]/P0001  ;
  input \u0_u0_ch_adr0_r_reg[14]/P0001  ;
  input \u0_u0_ch_adr0_r_reg[15]/P0001  ;
  input \u0_u0_ch_adr0_r_reg[16]/P0001  ;
  input \u0_u0_ch_adr0_r_reg[17]/P0001  ;
  input \u0_u0_ch_adr0_r_reg[18]/P0001  ;
  input \u0_u0_ch_adr0_r_reg[19]/P0001  ;
  input \u0_u0_ch_adr0_r_reg[1]/P0001  ;
  input \u0_u0_ch_adr0_r_reg[20]/P0001  ;
  input \u0_u0_ch_adr0_r_reg[21]/P0001  ;
  input \u0_u0_ch_adr0_r_reg[22]/P0001  ;
  input \u0_u0_ch_adr0_r_reg[23]/P0001  ;
  input \u0_u0_ch_adr0_r_reg[24]/P0001  ;
  input \u0_u0_ch_adr0_r_reg[25]/P0001  ;
  input \u0_u0_ch_adr0_r_reg[26]/P0001  ;
  input \u0_u0_ch_adr0_r_reg[27]/P0001  ;
  input \u0_u0_ch_adr0_r_reg[28]/P0001  ;
  input \u0_u0_ch_adr0_r_reg[29]/P0001  ;
  input \u0_u0_ch_adr0_r_reg[2]/P0001  ;
  input \u0_u0_ch_adr0_r_reg[3]/P0001  ;
  input \u0_u0_ch_adr0_r_reg[4]/P0001  ;
  input \u0_u0_ch_adr0_r_reg[5]/P0001  ;
  input \u0_u0_ch_adr0_r_reg[6]/P0001  ;
  input \u0_u0_ch_adr0_r_reg[7]/P0001  ;
  input \u0_u0_ch_adr0_r_reg[8]/P0001  ;
  input \u0_u0_ch_adr0_r_reg[9]/P0001  ;
  input \u0_u0_ch_adr1_r_reg[0]/P0001  ;
  input \u0_u0_ch_adr1_r_reg[10]/P0001  ;
  input \u0_u0_ch_adr1_r_reg[11]/P0001  ;
  input \u0_u0_ch_adr1_r_reg[12]/P0001  ;
  input \u0_u0_ch_adr1_r_reg[13]/P0001  ;
  input \u0_u0_ch_adr1_r_reg[14]/P0001  ;
  input \u0_u0_ch_adr1_r_reg[15]/P0001  ;
  input \u0_u0_ch_adr1_r_reg[16]/P0001  ;
  input \u0_u0_ch_adr1_r_reg[17]/P0001  ;
  input \u0_u0_ch_adr1_r_reg[18]/P0001  ;
  input \u0_u0_ch_adr1_r_reg[19]/P0001  ;
  input \u0_u0_ch_adr1_r_reg[1]/P0001  ;
  input \u0_u0_ch_adr1_r_reg[20]/P0001  ;
  input \u0_u0_ch_adr1_r_reg[21]/P0001  ;
  input \u0_u0_ch_adr1_r_reg[22]/P0001  ;
  input \u0_u0_ch_adr1_r_reg[23]/P0001  ;
  input \u0_u0_ch_adr1_r_reg[24]/P0001  ;
  input \u0_u0_ch_adr1_r_reg[25]/P0001  ;
  input \u0_u0_ch_adr1_r_reg[26]/P0001  ;
  input \u0_u0_ch_adr1_r_reg[27]/P0001  ;
  input \u0_u0_ch_adr1_r_reg[28]/P0001  ;
  input \u0_u0_ch_adr1_r_reg[29]/P0001  ;
  input \u0_u0_ch_adr1_r_reg[2]/P0001  ;
  input \u0_u0_ch_adr1_r_reg[3]/P0001  ;
  input \u0_u0_ch_adr1_r_reg[4]/P0001  ;
  input \u0_u0_ch_adr1_r_reg[5]/P0001  ;
  input \u0_u0_ch_adr1_r_reg[6]/P0001  ;
  input \u0_u0_ch_adr1_r_reg[7]/P0001  ;
  input \u0_u0_ch_adr1_r_reg[8]/P0001  ;
  input \u0_u0_ch_adr1_r_reg[9]/P0001  ;
  input \u0_u0_ch_busy_reg/P0001  ;
  input \u0_u0_ch_chk_sz_r_reg[0]/P0001  ;
  input \u0_u0_ch_chk_sz_r_reg[10]/P0001  ;
  input \u0_u0_ch_chk_sz_r_reg[1]/P0001  ;
  input \u0_u0_ch_chk_sz_r_reg[2]/P0001  ;
  input \u0_u0_ch_chk_sz_r_reg[3]/P0001  ;
  input \u0_u0_ch_chk_sz_r_reg[4]/P0001  ;
  input \u0_u0_ch_chk_sz_r_reg[5]/P0001  ;
  input \u0_u0_ch_chk_sz_r_reg[6]/P0001  ;
  input \u0_u0_ch_chk_sz_r_reg[7]/P0001  ;
  input \u0_u0_ch_chk_sz_r_reg[8]/P0001  ;
  input \u0_u0_ch_chk_sz_r_reg[9]/P0001  ;
  input \u0_u0_ch_csr_r2_reg[0]/NET0131  ;
  input \u0_u0_ch_csr_r2_reg[1]/NET0131  ;
  input \u0_u0_ch_csr_r2_reg[2]/NET0131  ;
  input \u0_u0_ch_csr_r3_reg[0]/NET0131  ;
  input \u0_u0_ch_csr_r3_reg[1]/NET0131  ;
  input \u0_u0_ch_csr_r3_reg[2]/NET0131  ;
  input \u0_u0_ch_csr_r_reg[0]/NET0131  ;
  input \u0_u0_ch_csr_r_reg[1]/NET0131  ;
  input \u0_u0_ch_csr_r_reg[2]/NET0131  ;
  input \u0_u0_ch_csr_r_reg[3]/NET0131  ;
  input \u0_u0_ch_csr_r_reg[4]/NET0131  ;
  input \u0_u0_ch_csr_r_reg[5]/NET0131  ;
  input \u0_u0_ch_csr_r_reg[6]/NET0131  ;
  input \u0_u0_ch_csr_r_reg[7]/NET0131  ;
  input \u0_u0_ch_csr_r_reg[8]/NET0131  ;
  input \u0_u0_ch_done_reg/P0002  ;
  input \u0_u0_ch_err_reg/NET0131  ;
  input \u0_u0_ch_stop_reg/P0001  ;
  input \u0_u0_ch_sz_inf_reg/NET0131  ;
  input \u0_u0_ch_tot_sz_r_reg[0]/P0001  ;
  input \u0_u0_ch_tot_sz_r_reg[10]/P0001  ;
  input \u0_u0_ch_tot_sz_r_reg[11]/P0001  ;
  input \u0_u0_ch_tot_sz_r_reg[1]/P0001  ;
  input \u0_u0_ch_tot_sz_r_reg[2]/P0001  ;
  input \u0_u0_ch_tot_sz_r_reg[3]/P0001  ;
  input \u0_u0_ch_tot_sz_r_reg[4]/P0001  ;
  input \u0_u0_ch_tot_sz_r_reg[5]/P0001  ;
  input \u0_u0_ch_tot_sz_r_reg[6]/P0001  ;
  input \u0_u0_ch_tot_sz_r_reg[7]/P0001  ;
  input \u0_u0_ch_tot_sz_r_reg[8]/P0001  ;
  input \u0_u0_ch_tot_sz_r_reg[9]/P0001  ;
  input \u0_u0_int_src_r_reg[1]/NET0131  ;
  input \u0_u0_int_src_r_reg[2]/NET0131  ;
  input \u0_u0_rest_en_reg/NET0131  ;
  input \u0_wb_rf_dout_reg[0]/P0001  ;
  input \u0_wb_rf_dout_reg[10]/P0001  ;
  input \u0_wb_rf_dout_reg[11]/P0001  ;
  input \u0_wb_rf_dout_reg[12]/P0001  ;
  input \u0_wb_rf_dout_reg[13]/P0001  ;
  input \u0_wb_rf_dout_reg[14]/P0001  ;
  input \u0_wb_rf_dout_reg[15]/P0001  ;
  input \u0_wb_rf_dout_reg[16]/P0001  ;
  input \u0_wb_rf_dout_reg[17]/P0001  ;
  input \u0_wb_rf_dout_reg[18]/P0001  ;
  input \u0_wb_rf_dout_reg[19]/P0001  ;
  input \u0_wb_rf_dout_reg[1]/P0001  ;
  input \u0_wb_rf_dout_reg[20]/P0001  ;
  input \u0_wb_rf_dout_reg[21]/P0001  ;
  input \u0_wb_rf_dout_reg[22]/P0001  ;
  input \u0_wb_rf_dout_reg[23]/P0001  ;
  input \u0_wb_rf_dout_reg[24]/P0001  ;
  input \u0_wb_rf_dout_reg[25]/P0001  ;
  input \u0_wb_rf_dout_reg[26]/P0001  ;
  input \u0_wb_rf_dout_reg[27]/P0001  ;
  input \u0_wb_rf_dout_reg[28]/P0001  ;
  input \u0_wb_rf_dout_reg[29]/P0001  ;
  input \u0_wb_rf_dout_reg[2]/P0001  ;
  input \u0_wb_rf_dout_reg[30]/P0001  ;
  input \u0_wb_rf_dout_reg[31]/P0001  ;
  input \u0_wb_rf_dout_reg[3]/P0001  ;
  input \u0_wb_rf_dout_reg[4]/P0001  ;
  input \u0_wb_rf_dout_reg[5]/P0001  ;
  input \u0_wb_rf_dout_reg[6]/P0001  ;
  input \u0_wb_rf_dout_reg[7]/P0001  ;
  input \u0_wb_rf_dout_reg[8]/P0001  ;
  input \u0_wb_rf_dout_reg[9]/P0001  ;
  input \u1_de_start_r_reg/P0001  ;
  input \u1_ndnr_reg[0]/P0001  ;
  input \u1_ndr_r_reg[0]/NET0131  ;
  input \u1_next_start_reg/P0001  ;
  input \u1_req_r_reg[0]/P0001  ;
  input \u2_adr0_cnt_reg[0]/P0001  ;
  input \u2_adr0_cnt_reg[10]/P0001  ;
  input \u2_adr0_cnt_reg[11]/P0001  ;
  input \u2_adr0_cnt_reg[12]/P0001  ;
  input \u2_adr0_cnt_reg[13]/P0001  ;
  input \u2_adr0_cnt_reg[14]/P0001  ;
  input \u2_adr0_cnt_reg[15]/P0001  ;
  input \u2_adr0_cnt_reg[16]/NET0131  ;
  input \u2_adr0_cnt_reg[17]/P0001  ;
  input \u2_adr0_cnt_reg[18]/P0001  ;
  input \u2_adr0_cnt_reg[19]/P0001  ;
  input \u2_adr0_cnt_reg[1]/P0001  ;
  input \u2_adr0_cnt_reg[20]/P0001  ;
  input \u2_adr0_cnt_reg[21]/P0001  ;
  input \u2_adr0_cnt_reg[22]/P0001  ;
  input \u2_adr0_cnt_reg[23]/P0001  ;
  input \u2_adr0_cnt_reg[24]/P0001  ;
  input \u2_adr0_cnt_reg[25]/P0001  ;
  input \u2_adr0_cnt_reg[26]/P0001  ;
  input \u2_adr0_cnt_reg[27]/P0001  ;
  input \u2_adr0_cnt_reg[28]/P0001  ;
  input \u2_adr0_cnt_reg[29]/P0001  ;
  input \u2_adr0_cnt_reg[2]/P0001  ;
  input \u2_adr0_cnt_reg[3]/P0001  ;
  input \u2_adr0_cnt_reg[4]/P0001  ;
  input \u2_adr0_cnt_reg[5]/P0001  ;
  input \u2_adr0_cnt_reg[6]/P0001  ;
  input \u2_adr0_cnt_reg[7]/P0001  ;
  input \u2_adr0_cnt_reg[8]/P0001  ;
  input \u2_adr0_cnt_reg[9]/P0001  ;
  input \u2_adr1_cnt_reg[0]/P0001  ;
  input \u2_adr1_cnt_reg[10]/P0001  ;
  input \u2_adr1_cnt_reg[11]/P0001  ;
  input \u2_adr1_cnt_reg[12]/P0001  ;
  input \u2_adr1_cnt_reg[13]/P0001  ;
  input \u2_adr1_cnt_reg[14]/P0001  ;
  input \u2_adr1_cnt_reg[15]/P0001  ;
  input \u2_adr1_cnt_reg[16]/NET0131  ;
  input \u2_adr1_cnt_reg[17]/P0001  ;
  input \u2_adr1_cnt_reg[18]/P0001  ;
  input \u2_adr1_cnt_reg[19]/P0001  ;
  input \u2_adr1_cnt_reg[1]/P0001  ;
  input \u2_adr1_cnt_reg[20]/P0001  ;
  input \u2_adr1_cnt_reg[21]/P0001  ;
  input \u2_adr1_cnt_reg[22]/P0001  ;
  input \u2_adr1_cnt_reg[23]/P0001  ;
  input \u2_adr1_cnt_reg[24]/P0001  ;
  input \u2_adr1_cnt_reg[25]/P0001  ;
  input \u2_adr1_cnt_reg[26]/P0001  ;
  input \u2_adr1_cnt_reg[27]/P0001  ;
  input \u2_adr1_cnt_reg[28]/P0001  ;
  input \u2_adr1_cnt_reg[29]/P0001  ;
  input \u2_adr1_cnt_reg[2]/P0001  ;
  input \u2_adr1_cnt_reg[3]/P0001  ;
  input \u2_adr1_cnt_reg[4]/P0001  ;
  input \u2_adr1_cnt_reg[5]/P0001  ;
  input \u2_adr1_cnt_reg[6]/P0001  ;
  input \u2_adr1_cnt_reg[7]/P0001  ;
  input \u2_adr1_cnt_reg[8]/P0001  ;
  input \u2_adr1_cnt_reg[9]/P0001  ;
  input \u2_chunk_0_reg/P0001  ;
  input \u2_chunk_cnt_is_0_r_reg/P0001  ;
  input \u2_chunk_cnt_reg[0]/NET0131  ;
  input \u2_chunk_cnt_reg[1]/NET0131  ;
  input \u2_chunk_cnt_reg[2]/NET0131  ;
  input \u2_chunk_cnt_reg[3]/NET0131  ;
  input \u2_chunk_cnt_reg[4]/NET0131  ;
  input \u2_chunk_cnt_reg[5]/NET0131  ;
  input \u2_chunk_cnt_reg[6]/NET0131  ;
  input \u2_chunk_cnt_reg[7]/NET0131  ;
  input \u2_chunk_cnt_reg[8]/NET0131  ;
  input \u2_chunk_dec_reg/P0001  ;
  input \u2_dma_abort_r_reg/NET0131  ;
  input \u2_mast0_adr_reg[10]/P0001  ;
  input \u2_mast0_adr_reg[11]/P0001  ;
  input \u2_mast0_adr_reg[12]/P0001  ;
  input \u2_mast0_adr_reg[13]/P0001  ;
  input \u2_mast0_adr_reg[14]/P0001  ;
  input \u2_mast0_adr_reg[15]/P0001  ;
  input \u2_mast0_adr_reg[16]/P0001  ;
  input \u2_mast0_adr_reg[17]/P0001  ;
  input \u2_mast0_adr_reg[18]/P0001  ;
  input \u2_mast0_adr_reg[19]/P0001  ;
  input \u2_mast0_adr_reg[20]/P0001  ;
  input \u2_mast0_adr_reg[21]/P0001  ;
  input \u2_mast0_adr_reg[22]/P0001  ;
  input \u2_mast0_adr_reg[23]/P0001  ;
  input \u2_mast0_adr_reg[24]/P0001  ;
  input \u2_mast0_adr_reg[25]/P0001  ;
  input \u2_mast0_adr_reg[26]/P0001  ;
  input \u2_mast0_adr_reg[27]/P0001  ;
  input \u2_mast0_adr_reg[28]/P0001  ;
  input \u2_mast0_adr_reg[29]/P0001  ;
  input \u2_mast0_adr_reg[2]/P0001  ;
  input \u2_mast0_adr_reg[30]/P0001  ;
  input \u2_mast0_adr_reg[31]/P0001  ;
  input \u2_mast0_adr_reg[3]/NET0131  ;
  input \u2_mast0_adr_reg[4]/P0001  ;
  input \u2_mast0_adr_reg[5]/P0001  ;
  input \u2_mast0_adr_reg[6]/P0001  ;
  input \u2_mast0_adr_reg[7]/P0001  ;
  input \u2_mast0_adr_reg[8]/P0001  ;
  input \u2_mast0_adr_reg[9]/P0001  ;
  input \u2_mast0_drdy_r_reg/P0001  ;
  input \u2_mast1_adr_reg[10]/P0001  ;
  input \u2_mast1_adr_reg[11]/P0001  ;
  input \u2_mast1_adr_reg[12]/P0001  ;
  input \u2_mast1_adr_reg[13]/P0001  ;
  input \u2_mast1_adr_reg[14]/P0001  ;
  input \u2_mast1_adr_reg[15]/P0001  ;
  input \u2_mast1_adr_reg[16]/P0001  ;
  input \u2_mast1_adr_reg[17]/P0001  ;
  input \u2_mast1_adr_reg[18]/P0001  ;
  input \u2_mast1_adr_reg[19]/P0001  ;
  input \u2_mast1_adr_reg[20]/P0001  ;
  input \u2_mast1_adr_reg[21]/P0001  ;
  input \u2_mast1_adr_reg[22]/P0001  ;
  input \u2_mast1_adr_reg[23]/P0001  ;
  input \u2_mast1_adr_reg[24]/P0001  ;
  input \u2_mast1_adr_reg[25]/P0001  ;
  input \u2_mast1_adr_reg[26]/P0001  ;
  input \u2_mast1_adr_reg[27]/P0001  ;
  input \u2_mast1_adr_reg[28]/P0001  ;
  input \u2_mast1_adr_reg[29]/P0001  ;
  input \u2_mast1_adr_reg[2]/P0001  ;
  input \u2_mast1_adr_reg[30]/P0001  ;
  input \u2_mast1_adr_reg[31]/P0001  ;
  input \u2_mast1_adr_reg[3]/P0001  ;
  input \u2_mast1_adr_reg[4]/P0001  ;
  input \u2_mast1_adr_reg[5]/P0001  ;
  input \u2_mast1_adr_reg[6]/P0001  ;
  input \u2_mast1_adr_reg[7]/P0001  ;
  input \u2_mast1_adr_reg[8]/P0001  ;
  input \u2_mast1_adr_reg[9]/P0001  ;
  input \u2_next_ch_reg/P0001  ;
  input \u2_read_r_reg/P0001  ;
  input \u2_state_reg[0]/NET0131  ;
  input \u2_state_reg[10]/NET0131  ;
  input \u2_state_reg[1]/NET0131  ;
  input \u2_state_reg[2]/NET0131  ;
  input \u2_state_reg[3]/NET0131  ;
  input \u2_state_reg[4]/NET0131  ;
  input \u2_state_reg[5]/NET0131  ;
  input \u2_state_reg[6]/NET0131  ;
  input \u2_state_reg[7]/NET0131  ;
  input \u2_state_reg[8]/NET0131  ;
  input \u2_state_reg[9]/NET0131  ;
  input \u2_tsz_cnt_is_0_r_reg/P0001  ;
  input \u2_tsz_cnt_reg[0]/NET0131  ;
  input \u2_tsz_cnt_reg[10]/NET0131  ;
  input \u2_tsz_cnt_reg[11]/NET0131  ;
  input \u2_tsz_cnt_reg[1]/NET0131  ;
  input \u2_tsz_cnt_reg[2]/NET0131  ;
  input \u2_tsz_cnt_reg[3]/NET0131  ;
  input \u2_tsz_cnt_reg[4]/NET0131  ;
  input \u2_tsz_cnt_reg[5]/NET0131  ;
  input \u2_tsz_cnt_reg[6]/NET0131  ;
  input \u2_tsz_cnt_reg[7]/NET0131  ;
  input \u2_tsz_cnt_reg[8]/NET0131  ;
  input \u2_tsz_cnt_reg[9]/NET0131  ;
  input \u2_u0_out_r_reg[0]/P0001  ;
  input \u2_u0_out_r_reg[10]/P0001  ;
  input \u2_u0_out_r_reg[11]/P0001  ;
  input \u2_u0_out_r_reg[12]/P0001  ;
  input \u2_u0_out_r_reg[13]/P0001  ;
  input \u2_u0_out_r_reg[14]/P0001  ;
  input \u2_u0_out_r_reg[15]/P0001  ;
  input \u2_u0_out_r_reg[16]/P0001  ;
  input \u2_u0_out_r_reg[1]/P0001  ;
  input \u2_u0_out_r_reg[2]/P0001  ;
  input \u2_u0_out_r_reg[3]/P0001  ;
  input \u2_u0_out_r_reg[4]/P0001  ;
  input \u2_u0_out_r_reg[5]/P0001  ;
  input \u2_u0_out_r_reg[6]/P0001  ;
  input \u2_u0_out_r_reg[7]/P0001  ;
  input \u2_u0_out_r_reg[8]/P0001  ;
  input \u2_u0_out_r_reg[9]/P0001  ;
  input \u2_u1_out_r_reg[0]/P0001  ;
  input \u2_u1_out_r_reg[10]/P0001  ;
  input \u2_u1_out_r_reg[11]/P0001  ;
  input \u2_u1_out_r_reg[12]/P0001  ;
  input \u2_u1_out_r_reg[13]/P0001  ;
  input \u2_u1_out_r_reg[14]/P0001  ;
  input \u2_u1_out_r_reg[15]/P0001  ;
  input \u2_u1_out_r_reg[16]/P0001  ;
  input \u2_u1_out_r_reg[1]/P0001  ;
  input \u2_u1_out_r_reg[2]/P0001  ;
  input \u2_u1_out_r_reg[3]/P0001  ;
  input \u2_u1_out_r_reg[4]/P0001  ;
  input \u2_u1_out_r_reg[5]/P0001  ;
  input \u2_u1_out_r_reg[6]/P0001  ;
  input \u2_u1_out_r_reg[7]/P0001  ;
  input \u2_u1_out_r_reg[8]/P0001  ;
  input \u2_u1_out_r_reg[9]/P0001  ;
  input \u2_write_hold_r_reg/P0001  ;
  input \u2_write_r_reg/P0001  ;
  input \u3_u0_mast_cyc_reg/P0001  ;
  input \u3_u0_mast_dout_reg[0]/P0001  ;
  input \u3_u0_mast_dout_reg[10]/P0001  ;
  input \u3_u0_mast_dout_reg[11]/P0001  ;
  input \u3_u0_mast_dout_reg[12]/P0001  ;
  input \u3_u0_mast_dout_reg[13]/P0001  ;
  input \u3_u0_mast_dout_reg[14]/P0001  ;
  input \u3_u0_mast_dout_reg[15]/P0001  ;
  input \u3_u0_mast_dout_reg[16]/P0001  ;
  input \u3_u0_mast_dout_reg[17]/P0001  ;
  input \u3_u0_mast_dout_reg[18]/P0001  ;
  input \u3_u0_mast_dout_reg[19]/P0001  ;
  input \u3_u0_mast_dout_reg[1]/P0001  ;
  input \u3_u0_mast_dout_reg[20]/P0001  ;
  input \u3_u0_mast_dout_reg[21]/P0001  ;
  input \u3_u0_mast_dout_reg[22]/P0001  ;
  input \u3_u0_mast_dout_reg[23]/P0001  ;
  input \u3_u0_mast_dout_reg[24]/P0001  ;
  input \u3_u0_mast_dout_reg[25]/P0001  ;
  input \u3_u0_mast_dout_reg[26]/P0001  ;
  input \u3_u0_mast_dout_reg[27]/P0001  ;
  input \u3_u0_mast_dout_reg[28]/P0001  ;
  input \u3_u0_mast_dout_reg[29]/P0001  ;
  input \u3_u0_mast_dout_reg[2]/P0001  ;
  input \u3_u0_mast_dout_reg[30]/P0001  ;
  input \u3_u0_mast_dout_reg[31]/P0001  ;
  input \u3_u0_mast_dout_reg[3]/P0001  ;
  input \u3_u0_mast_dout_reg[4]/P0001  ;
  input \u3_u0_mast_dout_reg[5]/P0001  ;
  input \u3_u0_mast_dout_reg[6]/P0001  ;
  input \u3_u0_mast_dout_reg[7]/P0001  ;
  input \u3_u0_mast_dout_reg[8]/P0001  ;
  input \u3_u0_mast_dout_reg[9]/P0001  ;
  input \u3_u0_mast_stb_reg/P0001  ;
  input \u3_u0_mast_we_r_reg/P0002  ;
  input \u3_u1_rf_ack_reg/P0001  ;
  input \u3_u1_slv_adr_reg[2]/NET0131  ;
  input \u3_u1_slv_adr_reg[3]/P0001  ;
  input \u3_u1_slv_adr_reg[4]/NET0131  ;
  input \u3_u1_slv_adr_reg[5]/P0001  ;
  input \u3_u1_slv_adr_reg[6]/NET0131  ;
  input \u3_u1_slv_adr_reg[7]/NET0131  ;
  input \u3_u1_slv_adr_reg[8]/NET0131  ;
  input \u3_u1_slv_adr_reg[9]/NET0131  ;
  input \u3_u1_slv_dout_reg[0]/P0001  ;
  input \u3_u1_slv_dout_reg[10]/P0001  ;
  input \u3_u1_slv_dout_reg[11]/P0001  ;
  input \u3_u1_slv_dout_reg[12]/P0001  ;
  input \u3_u1_slv_dout_reg[13]/P0001  ;
  input \u3_u1_slv_dout_reg[14]/P0001  ;
  input \u3_u1_slv_dout_reg[15]/P0001  ;
  input \u3_u1_slv_dout_reg[16]/P0001  ;
  input \u3_u1_slv_dout_reg[17]/P0001  ;
  input \u3_u1_slv_dout_reg[18]/P0001  ;
  input \u3_u1_slv_dout_reg[19]/P0001  ;
  input \u3_u1_slv_dout_reg[1]/P0001  ;
  input \u3_u1_slv_dout_reg[20]/P0001  ;
  input \u3_u1_slv_dout_reg[21]/P0001  ;
  input \u3_u1_slv_dout_reg[22]/P0001  ;
  input \u3_u1_slv_dout_reg[23]/P0001  ;
  input \u3_u1_slv_dout_reg[24]/P0001  ;
  input \u3_u1_slv_dout_reg[25]/P0001  ;
  input \u3_u1_slv_dout_reg[26]/P0001  ;
  input \u3_u1_slv_dout_reg[27]/P0001  ;
  input \u3_u1_slv_dout_reg[28]/P0001  ;
  input \u3_u1_slv_dout_reg[29]/P0001  ;
  input \u3_u1_slv_dout_reg[2]/P0001  ;
  input \u3_u1_slv_dout_reg[30]/P0001  ;
  input \u3_u1_slv_dout_reg[31]/P0001  ;
  input \u3_u1_slv_dout_reg[3]/P0001  ;
  input \u3_u1_slv_dout_reg[4]/P0001  ;
  input \u3_u1_slv_dout_reg[5]/P0001  ;
  input \u3_u1_slv_dout_reg[6]/P0001  ;
  input \u3_u1_slv_dout_reg[7]/P0001  ;
  input \u3_u1_slv_dout_reg[8]/P0001  ;
  input \u3_u1_slv_dout_reg[9]/P0001  ;
  input \u3_u1_slv_re_reg/P0001  ;
  input \u3_u1_slv_we_reg/P0001  ;
  input \u4_u0_mast_cyc_reg/P0001  ;
  input \u4_u0_mast_dout_reg[0]/P0001  ;
  input \u4_u0_mast_dout_reg[10]/P0001  ;
  input \u4_u0_mast_dout_reg[11]/P0001  ;
  input \u4_u0_mast_dout_reg[12]/P0001  ;
  input \u4_u0_mast_dout_reg[13]/P0001  ;
  input \u4_u0_mast_dout_reg[14]/P0001  ;
  input \u4_u0_mast_dout_reg[15]/P0001  ;
  input \u4_u0_mast_dout_reg[16]/P0001  ;
  input \u4_u0_mast_dout_reg[17]/P0001  ;
  input \u4_u0_mast_dout_reg[18]/P0001  ;
  input \u4_u0_mast_dout_reg[19]/P0001  ;
  input \u4_u0_mast_dout_reg[1]/P0001  ;
  input \u4_u0_mast_dout_reg[20]/P0001  ;
  input \u4_u0_mast_dout_reg[21]/P0001  ;
  input \u4_u0_mast_dout_reg[22]/P0001  ;
  input \u4_u0_mast_dout_reg[23]/P0001  ;
  input \u4_u0_mast_dout_reg[24]/P0001  ;
  input \u4_u0_mast_dout_reg[25]/P0001  ;
  input \u4_u0_mast_dout_reg[26]/P0001  ;
  input \u4_u0_mast_dout_reg[27]/P0001  ;
  input \u4_u0_mast_dout_reg[28]/P0001  ;
  input \u4_u0_mast_dout_reg[29]/P0001  ;
  input \u4_u0_mast_dout_reg[2]/P0001  ;
  input \u4_u0_mast_dout_reg[30]/P0001  ;
  input \u4_u0_mast_dout_reg[31]/P0001  ;
  input \u4_u0_mast_dout_reg[3]/P0001  ;
  input \u4_u0_mast_dout_reg[4]/P0001  ;
  input \u4_u0_mast_dout_reg[5]/P0001  ;
  input \u4_u0_mast_dout_reg[6]/P0001  ;
  input \u4_u0_mast_dout_reg[7]/P0001  ;
  input \u4_u0_mast_dout_reg[8]/P0001  ;
  input \u4_u0_mast_dout_reg[9]/P0001  ;
  input \u4_u0_mast_stb_reg/P0001  ;
  input \u4_u0_mast_we_r_reg/P0001  ;
  input \u4_u1_rf_ack_reg/P0001  ;
  input \u4_u1_slv_re_reg/P0001  ;
  input \u4_u1_slv_we_reg/P0001  ;
  input \wb0_ack_i_pad  ;
  input \wb0_addr_i[0]_pad  ;
  input \wb0_addr_i[10]_pad  ;
  input \wb0_addr_i[11]_pad  ;
  input \wb0_addr_i[12]_pad  ;
  input \wb0_addr_i[13]_pad  ;
  input \wb0_addr_i[14]_pad  ;
  input \wb0_addr_i[15]_pad  ;
  input \wb0_addr_i[16]_pad  ;
  input \wb0_addr_i[17]_pad  ;
  input \wb0_addr_i[18]_pad  ;
  input \wb0_addr_i[19]_pad  ;
  input \wb0_addr_i[1]_pad  ;
  input \wb0_addr_i[20]_pad  ;
  input \wb0_addr_i[21]_pad  ;
  input \wb0_addr_i[22]_pad  ;
  input \wb0_addr_i[23]_pad  ;
  input \wb0_addr_i[24]_pad  ;
  input \wb0_addr_i[25]_pad  ;
  input \wb0_addr_i[26]_pad  ;
  input \wb0_addr_i[27]_pad  ;
  input \wb0_addr_i[28]_pad  ;
  input \wb0_addr_i[29]_pad  ;
  input \wb0_addr_i[2]_pad  ;
  input \wb0_addr_i[30]_pad  ;
  input \wb0_addr_i[31]_pad  ;
  input \wb0_addr_i[3]_pad  ;
  input \wb0_addr_i[4]_pad  ;
  input \wb0_addr_i[5]_pad  ;
  input \wb0_addr_i[6]_pad  ;
  input \wb0_addr_i[7]_pad  ;
  input \wb0_addr_i[8]_pad  ;
  input \wb0_addr_i[9]_pad  ;
  input \wb0_cyc_i_pad  ;
  input \wb0_err_i_pad  ;
  input \wb0_rty_i_pad  ;
  input \wb0_sel_i[0]_pad  ;
  input \wb0_sel_i[1]_pad  ;
  input \wb0_sel_i[2]_pad  ;
  input \wb0_sel_i[3]_pad  ;
  input \wb0_stb_i_pad  ;
  input \wb0_we_i_pad  ;
  input \wb0m_data_i[0]_pad  ;
  input \wb0m_data_i[10]_pad  ;
  input \wb0m_data_i[11]_pad  ;
  input \wb0m_data_i[12]_pad  ;
  input \wb0m_data_i[13]_pad  ;
  input \wb0m_data_i[14]_pad  ;
  input \wb0m_data_i[15]_pad  ;
  input \wb0m_data_i[16]_pad  ;
  input \wb0m_data_i[17]_pad  ;
  input \wb0m_data_i[18]_pad  ;
  input \wb0m_data_i[19]_pad  ;
  input \wb0m_data_i[1]_pad  ;
  input \wb0m_data_i[20]_pad  ;
  input \wb0m_data_i[21]_pad  ;
  input \wb0m_data_i[22]_pad  ;
  input \wb0m_data_i[23]_pad  ;
  input \wb0m_data_i[24]_pad  ;
  input \wb0m_data_i[25]_pad  ;
  input \wb0m_data_i[26]_pad  ;
  input \wb0m_data_i[27]_pad  ;
  input \wb0m_data_i[28]_pad  ;
  input \wb0m_data_i[29]_pad  ;
  input \wb0m_data_i[2]_pad  ;
  input \wb0m_data_i[30]_pad  ;
  input \wb0m_data_i[31]_pad  ;
  input \wb0m_data_i[3]_pad  ;
  input \wb0m_data_i[4]_pad  ;
  input \wb0m_data_i[5]_pad  ;
  input \wb0m_data_i[6]_pad  ;
  input \wb0m_data_i[7]_pad  ;
  input \wb0m_data_i[8]_pad  ;
  input \wb0m_data_i[9]_pad  ;
  input \wb0s_data_i[0]_pad  ;
  input \wb0s_data_i[10]_pad  ;
  input \wb0s_data_i[11]_pad  ;
  input \wb0s_data_i[12]_pad  ;
  input \wb0s_data_i[13]_pad  ;
  input \wb0s_data_i[14]_pad  ;
  input \wb0s_data_i[15]_pad  ;
  input \wb0s_data_i[16]_pad  ;
  input \wb0s_data_i[17]_pad  ;
  input \wb0s_data_i[18]_pad  ;
  input \wb0s_data_i[19]_pad  ;
  input \wb0s_data_i[1]_pad  ;
  input \wb0s_data_i[20]_pad  ;
  input \wb0s_data_i[21]_pad  ;
  input \wb0s_data_i[22]_pad  ;
  input \wb0s_data_i[23]_pad  ;
  input \wb0s_data_i[24]_pad  ;
  input \wb0s_data_i[25]_pad  ;
  input \wb0s_data_i[26]_pad  ;
  input \wb0s_data_i[27]_pad  ;
  input \wb0s_data_i[28]_pad  ;
  input \wb0s_data_i[29]_pad  ;
  input \wb0s_data_i[2]_pad  ;
  input \wb0s_data_i[30]_pad  ;
  input \wb0s_data_i[31]_pad  ;
  input \wb0s_data_i[3]_pad  ;
  input \wb0s_data_i[4]_pad  ;
  input \wb0s_data_i[5]_pad  ;
  input \wb0s_data_i[6]_pad  ;
  input \wb0s_data_i[7]_pad  ;
  input \wb0s_data_i[8]_pad  ;
  input \wb0s_data_i[9]_pad  ;
  input \wb1_ack_i_pad  ;
  input \wb1_addr_i[0]_pad  ;
  input \wb1_addr_i[10]_pad  ;
  input \wb1_addr_i[11]_pad  ;
  input \wb1_addr_i[12]_pad  ;
  input \wb1_addr_i[13]_pad  ;
  input \wb1_addr_i[14]_pad  ;
  input \wb1_addr_i[15]_pad  ;
  input \wb1_addr_i[16]_pad  ;
  input \wb1_addr_i[17]_pad  ;
  input \wb1_addr_i[18]_pad  ;
  input \wb1_addr_i[19]_pad  ;
  input \wb1_addr_i[1]_pad  ;
  input \wb1_addr_i[20]_pad  ;
  input \wb1_addr_i[21]_pad  ;
  input \wb1_addr_i[22]_pad  ;
  input \wb1_addr_i[23]_pad  ;
  input \wb1_addr_i[24]_pad  ;
  input \wb1_addr_i[25]_pad  ;
  input \wb1_addr_i[26]_pad  ;
  input \wb1_addr_i[27]_pad  ;
  input \wb1_addr_i[28]_pad  ;
  input \wb1_addr_i[29]_pad  ;
  input \wb1_addr_i[2]_pad  ;
  input \wb1_addr_i[30]_pad  ;
  input \wb1_addr_i[31]_pad  ;
  input \wb1_addr_i[3]_pad  ;
  input \wb1_addr_i[4]_pad  ;
  input \wb1_addr_i[5]_pad  ;
  input \wb1_addr_i[6]_pad  ;
  input \wb1_addr_i[7]_pad  ;
  input \wb1_addr_i[8]_pad  ;
  input \wb1_addr_i[9]_pad  ;
  input \wb1_cyc_i_pad  ;
  input \wb1_err_i_pad  ;
  input \wb1_rty_i_pad  ;
  input \wb1_sel_i[0]_pad  ;
  input \wb1_sel_i[1]_pad  ;
  input \wb1_sel_i[2]_pad  ;
  input \wb1_sel_i[3]_pad  ;
  input \wb1_stb_i_pad  ;
  input \wb1_we_i_pad  ;
  input \wb1m_data_i[0]_pad  ;
  input \wb1m_data_i[10]_pad  ;
  input \wb1m_data_i[11]_pad  ;
  input \wb1m_data_i[12]_pad  ;
  input \wb1m_data_i[13]_pad  ;
  input \wb1m_data_i[14]_pad  ;
  input \wb1m_data_i[15]_pad  ;
  input \wb1m_data_i[16]_pad  ;
  input \wb1m_data_i[17]_pad  ;
  input \wb1m_data_i[18]_pad  ;
  input \wb1m_data_i[19]_pad  ;
  input \wb1m_data_i[1]_pad  ;
  input \wb1m_data_i[20]_pad  ;
  input \wb1m_data_i[21]_pad  ;
  input \wb1m_data_i[22]_pad  ;
  input \wb1m_data_i[23]_pad  ;
  input \wb1m_data_i[24]_pad  ;
  input \wb1m_data_i[25]_pad  ;
  input \wb1m_data_i[26]_pad  ;
  input \wb1m_data_i[27]_pad  ;
  input \wb1m_data_i[28]_pad  ;
  input \wb1m_data_i[29]_pad  ;
  input \wb1m_data_i[2]_pad  ;
  input \wb1m_data_i[30]_pad  ;
  input \wb1m_data_i[31]_pad  ;
  input \wb1m_data_i[3]_pad  ;
  input \wb1m_data_i[4]_pad  ;
  input \wb1m_data_i[5]_pad  ;
  input \wb1m_data_i[6]_pad  ;
  input \wb1m_data_i[7]_pad  ;
  input \wb1m_data_i[8]_pad  ;
  input \wb1m_data_i[9]_pad  ;
  input \wb1s_data_i[0]_pad  ;
  input \wb1s_data_i[10]_pad  ;
  input \wb1s_data_i[11]_pad  ;
  input \wb1s_data_i[12]_pad  ;
  input \wb1s_data_i[13]_pad  ;
  input \wb1s_data_i[14]_pad  ;
  input \wb1s_data_i[15]_pad  ;
  input \wb1s_data_i[16]_pad  ;
  input \wb1s_data_i[17]_pad  ;
  input \wb1s_data_i[18]_pad  ;
  input \wb1s_data_i[19]_pad  ;
  input \wb1s_data_i[1]_pad  ;
  input \wb1s_data_i[20]_pad  ;
  input \wb1s_data_i[21]_pad  ;
  input \wb1s_data_i[22]_pad  ;
  input \wb1s_data_i[23]_pad  ;
  input \wb1s_data_i[24]_pad  ;
  input \wb1s_data_i[25]_pad  ;
  input \wb1s_data_i[26]_pad  ;
  input \wb1s_data_i[27]_pad  ;
  input \wb1s_data_i[28]_pad  ;
  input \wb1s_data_i[29]_pad  ;
  input \wb1s_data_i[2]_pad  ;
  input \wb1s_data_i[30]_pad  ;
  input \wb1s_data_i[31]_pad  ;
  input \wb1s_data_i[3]_pad  ;
  input \wb1s_data_i[4]_pad  ;
  input \wb1s_data_i[5]_pad  ;
  input \wb1s_data_i[6]_pad  ;
  input \wb1s_data_i[7]_pad  ;
  input \wb1s_data_i[8]_pad  ;
  input \wb1s_data_i[9]_pad  ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g22594/_0_  ;
  output \g22595/_0_  ;
  output \g22599/_0_  ;
  output \g22600/_0_  ;
  output \g22606/_0_  ;
  output \g22607/_0_  ;
  output \g22610/_0_  ;
  output \g22614/_0_  ;
  output \g22615/_0_  ;
  output \g22616/_0_  ;
  output \g22619/_0_  ;
  output \g22620/_0_  ;
  output \g22626/_0_  ;
  output \g22635/_0_  ;
  output \g22650/_0_  ;
  output \g22651/_0_  ;
  output \g22692/_0_  ;
  output \g22727/_0_  ;
  output \g22729/_3_  ;
  output \g22774/_0_  ;
  output \g22775/_0_  ;
  output \g22776/_0_  ;
  output \g22777/_0_  ;
  output \g22779/_3_  ;
  output \g22780/_0_  ;
  output \g22781/_0_  ;
  output \g22782/_0_  ;
  output \g22784/_0_  ;
  output \g22785/_0_  ;
  output \g22786/_0_  ;
  output \g22787/_0_  ;
  output \g22789/_3_  ;
  output \g22790/_0_  ;
  output \g22791/_0_  ;
  output \g22792/_0_  ;
  output \g22793/_0_  ;
  output \g22794/_0_  ;
  output \g22795/_0_  ;
  output \g22796/_0_  ;
  output \g22797/_0_  ;
  output \g22798/_0_  ;
  output \g22799/_0_  ;
  output \g22838/_0_  ;
  output \g22839/_0_  ;
  output \g22841/_0_  ;
  output \g22842/_0_  ;
  output \g22847/_0_  ;
  output \g22848/_0_  ;
  output \g22849/_0_  ;
  output \g22850/_0_  ;
  output \g22851/_0_  ;
  output \g22852/_0_  ;
  output \g22853/_0_  ;
  output \g22854/_0_  ;
  output \g22855/_0_  ;
  output \g22856/_0_  ;
  output \g22857/_0_  ;
  output \g22858/_0_  ;
  output \g22859/_0_  ;
  output \g22860/_0_  ;
  output \g22861/_0_  ;
  output \g22862/_0_  ;
  output \g22863/_0_  ;
  output \g22864/_0_  ;
  output \g22865/_0_  ;
  output \g22867/_0_  ;
  output \g22868/_0_  ;
  output \g22869/_0_  ;
  output \g22871/_0_  ;
  output \g22872/_0_  ;
  output \g22873/_0_  ;
  output \g22874/_0_  ;
  output \g22875/_0_  ;
  output \g22876/_0_  ;
  output \g22878/_0_  ;
  output \g22882/_2_  ;
  output \g22995/_0_  ;
  output \g23030/_0_  ;
  output \g23046/_0_  ;
  output \g23077/_0_  ;
  output \g23111/_0_  ;
  output \g23115/_1_  ;
  output \g23124/_2_  ;
  output \g23126/_2_  ;
  output \g23128/_2_  ;
  output \g23130/_2_  ;
  output \g23132/_2_  ;
  output \g23134/_2_  ;
  output \g23136/_2_  ;
  output \g23137/_0_  ;
  output \g23140/_2_  ;
  output \g23142/_2_  ;
  output \g23144/_2_  ;
  output \g23146/_2_  ;
  output \g23148/_2_  ;
  output \g23150/_2_  ;
  output \g23152/_2_  ;
  output \g23154/_2_  ;
  output \g23156/_2_  ;
  output \g23158/_2_  ;
  output \g23160/_2_  ;
  output \g23162/_2_  ;
  output \g23163/_3_  ;
  output \g23164/_0_  ;
  output \g23166/_0_  ;
  output \g23168/_0_  ;
  output \g23170/_2_  ;
  output \g23172/_2_  ;
  output \g23174/_2_  ;
  output \g23175/_0_  ;
  output \g23177/_0_  ;
  output \g23180/_2_  ;
  output \g23220/_0_  ;
  output \g23238/_0_  ;
  output \g23239/_0_  ;
  output \g23240/_0_  ;
  output \g23241/_0_  ;
  output \g23242/_0_  ;
  output \g23243/_0_  ;
  output \g23244/_0_  ;
  output \g23245/_0_  ;
  output \g23247/_3_  ;
  output \g23248/_0_  ;
  output \g23249/_0_  ;
  output \g23250/_0_  ;
  output \g23251/_0_  ;
  output \g23252/_0_  ;
  output \g23253/_0_  ;
  output \g23255/_3_  ;
  output \g23260/_0_  ;
  output \g23284/_3_  ;
  output \g23285/_0_  ;
  output \g23334/_0_  ;
  output \g23343/_0_  ;
  output \g23366/_0_  ;
  output \g23402/_0_  ;
  output \g23403/_0_  ;
  output \g23404/_0_  ;
  output \g23405/_0_  ;
  output \g23407/_0_  ;
  output \g23408/_0_  ;
  output \g23409/_0_  ;
  output \g23410/_0_  ;
  output \g23411/_0_  ;
  output \g23413/_2_  ;
  output \g23415/_2_  ;
  output \g23417/_2_  ;
  output \g23542/_0_  ;
  output \g23607/_0_  ;
  output \g23608/_0_  ;
  output \g23609/_3_  ;
  output \g23707/_0_  ;
  output \g23708/_0_  ;
  output \g23709/_0_  ;
  output \g23710/_0_  ;
  output \g23711/_0_  ;
  output \g23712/_0_  ;
  output \g23713/_0_  ;
  output \g23714/_0_  ;
  output \g23715/_0_  ;
  output \g23716/_0_  ;
  output \g23754/_0_  ;
  output \g23755/_0_  ;
  output \g23756/_0_  ;
  output \g23757/_0_  ;
  output \g23758/_0_  ;
  output \g23759/_0_  ;
  output \g23760/_0_  ;
  output \g23761/_0_  ;
  output \g23763/_3_  ;
  output \g23767/_0_  ;
  output \g23768/_0_  ;
  output \g23833/_0_  ;
  output \g23837/_0_  ;
  output \g23838/_0_  ;
  output \g23839/_0_  ;
  output \g23840/_0_  ;
  output \g23841/_0_  ;
  output \g23842/_0_  ;
  output \g23843/_0_  ;
  output \g23844/_0_  ;
  output \g23845/_0_  ;
  output \g23849/_3_  ;
  output \g23851/_3_  ;
  output \g23858/_0_  ;
  output \g23870/_0_  ;
  output \g23871/_0_  ;
  output \g23872/_3_  ;
  output \g23873/_3_  ;
  output \g23874/_3_  ;
  output \g23875/_3_  ;
  output \g23876/_3_  ;
  output \g23877/_3_  ;
  output \g23878/_3_  ;
  output \g23879/_3_  ;
  output \g23880/_3_  ;
  output \g23881/_3_  ;
  output \g23882/_3_  ;
  output \g23883/_3_  ;
  output \g23884/_3_  ;
  output \g23885/_3_  ;
  output \g23886/_3_  ;
  output \g23887/_3_  ;
  output \g23888/_3_  ;
  output \g23889/_3_  ;
  output \g23890/_3_  ;
  output \g23891/_3_  ;
  output \g23892/_3_  ;
  output \g23893/_3_  ;
  output \g23894/_3_  ;
  output \g23895/_3_  ;
  output \g23896/_3_  ;
  output \g23897/_3_  ;
  output \g23898/_3_  ;
  output \g23899/_3_  ;
  output \g23900/_3_  ;
  output \g23901/_3_  ;
  output \g23902/_3_  ;
  output \g23903/_3_  ;
  output \g23904/_3_  ;
  output \g23905/_3_  ;
  output \g23906/_3_  ;
  output \g23907/_3_  ;
  output \g23908/_3_  ;
  output \g23909/_3_  ;
  output \g23910/_3_  ;
  output \g23911/_3_  ;
  output \g23912/_3_  ;
  output \g23913/_3_  ;
  output \g23914/_3_  ;
  output \g23915/_3_  ;
  output \g23959/_0_  ;
  output \g23961/_0_  ;
  output \g23962/_0_  ;
  output \g23966/_0_  ;
  output \g23967/_0_  ;
  output \g23969/_0_  ;
  output \g23970/_0_  ;
  output \g23971/_0_  ;
  output \g23972/_0_  ;
  output \g23979/_0_  ;
  output \g23987/_0_  ;
  output \g23988/_0_  ;
  output \g23989/_0_  ;
  output \g23990/_0_  ;
  output \g24005/_0_  ;
  output \g24010/_0_  ;
  output \g24012/_0_  ;
  output \g24013/_0_  ;
  output \g24014/_0_  ;
  output \g24015/_0_  ;
  output \g24016/_0_  ;
  output \g24017/_0_  ;
  output \g24018/_0_  ;
  output \g24019/_0_  ;
  output \g24020/_0_  ;
  output \g24026/_0_  ;
  output \g24027/_0_  ;
  output \g24028/_0_  ;
  output \g24029/_0_  ;
  output \g24030/_0_  ;
  output \g24031/_0_  ;
  output \g24032/_0_  ;
  output \g24033/_0_  ;
  output \g24034/_0_  ;
  output \g24035/_0_  ;
  output \g24036/_0_  ;
  output \g24037/_0_  ;
  output \g24038/_0_  ;
  output \g24039/_0_  ;
  output \g24042/_0_  ;
  output \g24049/_0_  ;
  output \g24063/_0_  ;
  output \g24119/_0_  ;
  output \g24120/_0_  ;
  output \g24357/_0_  ;
  output \g24432/_0_  ;
  output \g24433/_0_  ;
  output \g24437/_0_  ;
  output \g24438/_0_  ;
  output \g24477/_0_  ;
  output \g24491/_0_  ;
  output \g24530/_2_  ;
  output \g24532/_0_  ;
  output \g24534/_0_  ;
  output \g24537/_0_  ;
  output \g24538/_0_  ;
  output \g24539/_0_  ;
  output \g24540/_0_  ;
  output \g24606/_2_  ;
  output \g24612/_0_  ;
  output \g24677/_0_  ;
  output \g24678/_0_  ;
  output \g24679/_0_  ;
  output \g24688/_0_  ;
  output \g24743/_0_  ;
  output \g24847/_0_  ;
  output \g24849/_0_  ;
  output \g24850/_0_  ;
  output \g24854/_0_  ;
  output \g24862/_0_  ;
  output \g24872/_0_  ;
  output \g24873/_0_  ;
  output \g24874/_0_  ;
  output \g24876/_0_  ;
  output \g24879/_0_  ;
  output \g24880/_0_  ;
  output \g24881/_0_  ;
  output \g24882/_0_  ;
  output \g24952/_2_  ;
  output \g24976/_1_  ;
  output \g25003/_0_  ;
  output \g25004/_0_  ;
  output \g25005/_0_  ;
  output \g25006/_0_  ;
  output \g25011/_0_  ;
  output \g25012/_0_  ;
  output \g25013/_0_  ;
  output \g25031/_0_  ;
  output \g25032/_0_  ;
  output \g25033/_0_  ;
  output \g25034/_0_  ;
  output \g25035/_0_  ;
  output \g25153/_2_  ;
  output \g25183/_0_  ;
  output \g25184/_0_  ;
  output \g25224/_0_  ;
  output \g25232/_0_  ;
  output \g25237/_0_  ;
  output \g25241/_2_  ;
  output \g25243/_2_  ;
  output \g25248/_3_  ;
  output \g25261/_0_  ;
  output \g25262/_0_  ;
  output \g25266/_3_  ;
  output \g25267/_0_  ;
  output \g25269/_0_  ;
  output \g25543/_1_  ;
  output \g25602/_3_  ;
  output \g25610/_0_  ;
  output \g25611/_0_  ;
  output \g25841/_0_  ;
  output \g25843/_0_  ;
  output \g25893/_0_  ;
  output \g27013/_0_  ;
  output \g27060/_0_  ;
  output \g27073/_0_  ;
  output \g27184/_0_  ;
  output \g27186/_0_  ;
  output \g27189/_2_  ;
  output \g47/_0_  ;
  output \u0_u0_ch_done_reg/_05_  ;
  output \u2_adr0_cnt_reg[0]/P0000  ;
  output \u2_adr1_cnt_reg[0]/P0000  ;
  output \u3_u0_mast_we_r_reg/_05_  ;
  output \wb0_ack_o_pad  ;
  output \wb0_addr_o[0]_pad  ;
  output \wb0_addr_o[10]_pad  ;
  output \wb0_addr_o[11]_pad  ;
  output \wb0_addr_o[12]_pad  ;
  output \wb0_addr_o[13]_pad  ;
  output \wb0_addr_o[14]_pad  ;
  output \wb0_addr_o[15]_pad  ;
  output \wb0_addr_o[16]_pad  ;
  output \wb0_addr_o[17]_pad  ;
  output \wb0_addr_o[18]_pad  ;
  output \wb0_addr_o[19]_pad  ;
  output \wb0_addr_o[1]_pad  ;
  output \wb0_addr_o[20]_pad  ;
  output \wb0_addr_o[21]_pad  ;
  output \wb0_addr_o[22]_pad  ;
  output \wb0_addr_o[23]_pad  ;
  output \wb0_addr_o[24]_pad  ;
  output \wb0_addr_o[25]_pad  ;
  output \wb0_addr_o[26]_pad  ;
  output \wb0_addr_o[27]_pad  ;
  output \wb0_addr_o[28]_pad  ;
  output \wb0_addr_o[29]_pad  ;
  output \wb0_addr_o[2]_pad  ;
  output \wb0_addr_o[30]_pad  ;
  output \wb0_addr_o[31]_pad  ;
  output \wb0_addr_o[3]_pad  ;
  output \wb0_addr_o[4]_pad  ;
  output \wb0_addr_o[5]_pad  ;
  output \wb0_addr_o[6]_pad  ;
  output \wb0_addr_o[7]_pad  ;
  output \wb0_addr_o[8]_pad  ;
  output \wb0_addr_o[9]_pad  ;
  output \wb0_cyc_o_pad  ;
  output \wb0_err_o_pad  ;
  output \wb0_rty_o_pad  ;
  output \wb0_sel_o[0]_pad  ;
  output \wb0_sel_o[1]_pad  ;
  output \wb0_sel_o[2]_pad  ;
  output \wb0_sel_o[3]_pad  ;
  output \wb0_stb_o_pad  ;
  output \wb0_we_o_pad  ;
  output \wb0m_data_o[0]_pad  ;
  output \wb0m_data_o[10]_pad  ;
  output \wb0m_data_o[11]_pad  ;
  output \wb0m_data_o[12]_pad  ;
  output \wb0m_data_o[13]_pad  ;
  output \wb0m_data_o[14]_pad  ;
  output \wb0m_data_o[15]_pad  ;
  output \wb0m_data_o[16]_pad  ;
  output \wb0m_data_o[17]_pad  ;
  output \wb0m_data_o[18]_pad  ;
  output \wb0m_data_o[19]_pad  ;
  output \wb0m_data_o[1]_pad  ;
  output \wb0m_data_o[20]_pad  ;
  output \wb0m_data_o[21]_pad  ;
  output \wb0m_data_o[22]_pad  ;
  output \wb0m_data_o[23]_pad  ;
  output \wb0m_data_o[24]_pad  ;
  output \wb0m_data_o[25]_pad  ;
  output \wb0m_data_o[26]_pad  ;
  output \wb0m_data_o[27]_pad  ;
  output \wb0m_data_o[28]_pad  ;
  output \wb0m_data_o[29]_pad  ;
  output \wb0m_data_o[2]_pad  ;
  output \wb0m_data_o[30]_pad  ;
  output \wb0m_data_o[31]_pad  ;
  output \wb0m_data_o[3]_pad  ;
  output \wb0m_data_o[4]_pad  ;
  output \wb0m_data_o[5]_pad  ;
  output \wb0m_data_o[6]_pad  ;
  output \wb0m_data_o[7]_pad  ;
  output \wb0m_data_o[8]_pad  ;
  output \wb0m_data_o[9]_pad  ;
  output \wb0s_data_o[0]_pad  ;
  output \wb0s_data_o[10]_pad  ;
  output \wb0s_data_o[11]_pad  ;
  output \wb0s_data_o[12]_pad  ;
  output \wb0s_data_o[13]_pad  ;
  output \wb0s_data_o[14]_pad  ;
  output \wb0s_data_o[15]_pad  ;
  output \wb0s_data_o[16]_pad  ;
  output \wb0s_data_o[17]_pad  ;
  output \wb0s_data_o[18]_pad  ;
  output \wb0s_data_o[19]_pad  ;
  output \wb0s_data_o[1]_pad  ;
  output \wb0s_data_o[20]_pad  ;
  output \wb0s_data_o[21]_pad  ;
  output \wb0s_data_o[22]_pad  ;
  output \wb0s_data_o[23]_pad  ;
  output \wb0s_data_o[24]_pad  ;
  output \wb0s_data_o[25]_pad  ;
  output \wb0s_data_o[26]_pad  ;
  output \wb0s_data_o[27]_pad  ;
  output \wb0s_data_o[28]_pad  ;
  output \wb0s_data_o[29]_pad  ;
  output \wb0s_data_o[2]_pad  ;
  output \wb0s_data_o[30]_pad  ;
  output \wb0s_data_o[31]_pad  ;
  output \wb0s_data_o[3]_pad  ;
  output \wb0s_data_o[4]_pad  ;
  output \wb0s_data_o[5]_pad  ;
  output \wb0s_data_o[6]_pad  ;
  output \wb0s_data_o[7]_pad  ;
  output \wb0s_data_o[8]_pad  ;
  output \wb0s_data_o[9]_pad  ;
  output \wb1_ack_o_pad  ;
  output \wb1_addr_o[0]_pad  ;
  output \wb1_addr_o[10]_pad  ;
  output \wb1_addr_o[11]_pad  ;
  output \wb1_addr_o[12]_pad  ;
  output \wb1_addr_o[13]_pad  ;
  output \wb1_addr_o[14]_pad  ;
  output \wb1_addr_o[15]_pad  ;
  output \wb1_addr_o[16]_pad  ;
  output \wb1_addr_o[17]_pad  ;
  output \wb1_addr_o[18]_pad  ;
  output \wb1_addr_o[19]_pad  ;
  output \wb1_addr_o[1]_pad  ;
  output \wb1_addr_o[20]_pad  ;
  output \wb1_addr_o[21]_pad  ;
  output \wb1_addr_o[22]_pad  ;
  output \wb1_addr_o[23]_pad  ;
  output \wb1_addr_o[24]_pad  ;
  output \wb1_addr_o[25]_pad  ;
  output \wb1_addr_o[26]_pad  ;
  output \wb1_addr_o[27]_pad  ;
  output \wb1_addr_o[28]_pad  ;
  output \wb1_addr_o[29]_pad  ;
  output \wb1_addr_o[2]_pad  ;
  output \wb1_addr_o[30]_pad  ;
  output \wb1_addr_o[31]_pad  ;
  output \wb1_addr_o[3]_pad  ;
  output \wb1_addr_o[4]_pad  ;
  output \wb1_addr_o[5]_pad  ;
  output \wb1_addr_o[6]_pad  ;
  output \wb1_addr_o[7]_pad  ;
  output \wb1_addr_o[8]_pad  ;
  output \wb1_addr_o[9]_pad  ;
  output \wb1_cyc_o_pad  ;
  output \wb1_err_o_pad  ;
  output \wb1_rty_o_pad  ;
  output \wb1_sel_o[0]_pad  ;
  output \wb1_sel_o[1]_pad  ;
  output \wb1_sel_o[2]_pad  ;
  output \wb1_sel_o[3]_pad  ;
  output \wb1_stb_o_pad  ;
  output \wb1_we_o_pad  ;
  output \wb1m_data_o[0]_pad  ;
  output \wb1m_data_o[10]_pad  ;
  output \wb1m_data_o[11]_pad  ;
  output \wb1m_data_o[12]_pad  ;
  output \wb1m_data_o[13]_pad  ;
  output \wb1m_data_o[14]_pad  ;
  output \wb1m_data_o[15]_pad  ;
  output \wb1m_data_o[16]_pad  ;
  output \wb1m_data_o[17]_pad  ;
  output \wb1m_data_o[18]_pad  ;
  output \wb1m_data_o[19]_pad  ;
  output \wb1m_data_o[1]_pad  ;
  output \wb1m_data_o[20]_pad  ;
  output \wb1m_data_o[21]_pad  ;
  output \wb1m_data_o[22]_pad  ;
  output \wb1m_data_o[23]_pad  ;
  output \wb1m_data_o[24]_pad  ;
  output \wb1m_data_o[25]_pad  ;
  output \wb1m_data_o[26]_pad  ;
  output \wb1m_data_o[27]_pad  ;
  output \wb1m_data_o[28]_pad  ;
  output \wb1m_data_o[29]_pad  ;
  output \wb1m_data_o[2]_pad  ;
  output \wb1m_data_o[30]_pad  ;
  output \wb1m_data_o[31]_pad  ;
  output \wb1m_data_o[3]_pad  ;
  output \wb1m_data_o[4]_pad  ;
  output \wb1m_data_o[5]_pad  ;
  output \wb1m_data_o[6]_pad  ;
  output \wb1m_data_o[7]_pad  ;
  output \wb1m_data_o[8]_pad  ;
  output \wb1m_data_o[9]_pad  ;
  output \wb1s_data_o[0]_pad  ;
  output \wb1s_data_o[10]_pad  ;
  output \wb1s_data_o[11]_pad  ;
  output \wb1s_data_o[12]_pad  ;
  output \wb1s_data_o[13]_pad  ;
  output \wb1s_data_o[14]_pad  ;
  output \wb1s_data_o[15]_pad  ;
  output \wb1s_data_o[16]_pad  ;
  output \wb1s_data_o[17]_pad  ;
  output \wb1s_data_o[18]_pad  ;
  output \wb1s_data_o[19]_pad  ;
  output \wb1s_data_o[1]_pad  ;
  output \wb1s_data_o[20]_pad  ;
  output \wb1s_data_o[21]_pad  ;
  output \wb1s_data_o[22]_pad  ;
  output \wb1s_data_o[23]_pad  ;
  output \wb1s_data_o[24]_pad  ;
  output \wb1s_data_o[25]_pad  ;
  output \wb1s_data_o[26]_pad  ;
  output \wb1s_data_o[27]_pad  ;
  output \wb1s_data_o[28]_pad  ;
  output \wb1s_data_o[29]_pad  ;
  output \wb1s_data_o[2]_pad  ;
  output \wb1s_data_o[30]_pad  ;
  output \wb1s_data_o[31]_pad  ;
  output \wb1s_data_o[3]_pad  ;
  output \wb1s_data_o[4]_pad  ;
  output \wb1s_data_o[5]_pad  ;
  output \wb1s_data_o[6]_pad  ;
  output \wb1s_data_o[7]_pad  ;
  output \wb1s_data_o[8]_pad  ;
  output \wb1s_data_o[9]_pad  ;
  wire n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 ;
  assign n734 = ~\u0_u0_ch_csr_r_reg[1]/NET0131  & \wb0_ack_i_pad  ;
  assign n735 = \u0_u0_ch_csr_r_reg[1]/NET0131  & \wb1_ack_i_pad  ;
  assign n736 = ~n734 & ~n735 ;
  assign n737 = \u0_u0_ch_csr_r_reg[3]/NET0131  & \u2_write_r_reg/P0001  ;
  assign n738 = ~n736 & n737 ;
  assign n739 = \u2_adr1_cnt_reg[16]/NET0131  & \u2_u1_out_r_reg[16]/P0001  ;
  assign n740 = \u2_adr1_cnt_reg[17]/P0001  & n739 ;
  assign n741 = \u2_adr1_cnt_reg[19]/P0001  & \u2_adr1_cnt_reg[20]/P0001  ;
  assign n742 = \u2_adr1_cnt_reg[18]/P0001  & n741 ;
  assign n743 = n740 & n742 ;
  assign n744 = n738 & n743 ;
  assign n745 = \u2_adr1_cnt_reg[23]/P0001  & \u2_adr1_cnt_reg[24]/P0001  ;
  assign n746 = \u2_adr1_cnt_reg[25]/P0001  & n745 ;
  assign n747 = \u2_adr1_cnt_reg[21]/P0001  & \u2_adr1_cnt_reg[22]/P0001  ;
  assign n748 = \u2_adr1_cnt_reg[26]/P0001  & n747 ;
  assign n749 = n746 & n748 ;
  assign n750 = n744 & n749 ;
  assign n751 = \u2_adr1_cnt_reg[27]/P0001  & n750 ;
  assign n752 = ~dma_ack_o_pad & \u1_req_r_reg[0]/P0001  ;
  assign n753 = \u0_u0_ch_csr_r_reg[5]/NET0131  & ~n752 ;
  assign n754 = \u0_u0_ch_csr_r_reg[0]/NET0131  & ~\u1_de_start_r_reg/P0001  ;
  assign n755 = ~n753 & n754 ;
  assign n756 = ~\u1_next_start_reg/P0001  & ~\u2_state_reg[8]/NET0131  ;
  assign n757 = ~n755 & n756 ;
  assign n758 = \u2_adr1_cnt_reg[28]/P0001  & n757 ;
  assign n759 = ~n751 & n758 ;
  assign n760 = ~\u2_adr1_cnt_reg[28]/P0001  & n757 ;
  assign n761 = n751 & n760 ;
  assign n762 = ~n759 & ~n761 ;
  assign n763 = \u0_u0_ch_adr1_r_reg[28]/P0001  & ~n757 ;
  assign n764 = n762 & ~n763 ;
  assign n765 = \u0_u0_ch_csr_r_reg[2]/NET0131  & \wb1_ack_i_pad  ;
  assign n766 = ~\u0_u0_ch_csr_r_reg[2]/NET0131  & \wb0_ack_i_pad  ;
  assign n767 = ~n765 & ~n766 ;
  assign n768 = \u0_u0_ch_csr_r_reg[4]/NET0131  & \u2_read_r_reg/P0001  ;
  assign n769 = \u2_u0_out_r_reg[16]/P0001  & n768 ;
  assign n770 = ~n767 & n769 ;
  assign n771 = \u2_adr0_cnt_reg[16]/NET0131  & \u2_adr0_cnt_reg[17]/P0001  ;
  assign n772 = \u2_adr0_cnt_reg[18]/P0001  & \u2_adr0_cnt_reg[19]/P0001  ;
  assign n773 = n771 & n772 ;
  assign n774 = \u2_adr0_cnt_reg[20]/P0001  & n773 ;
  assign n775 = n770 & n774 ;
  assign n776 = \u2_adr0_cnt_reg[21]/P0001  & \u2_adr0_cnt_reg[22]/P0001  ;
  assign n777 = \u2_adr0_cnt_reg[23]/P0001  & n776 ;
  assign n778 = \u2_adr0_cnt_reg[24]/P0001  & \u2_adr0_cnt_reg[25]/P0001  ;
  assign n779 = \u2_adr0_cnt_reg[26]/P0001  & \u2_adr0_cnt_reg[27]/P0001  ;
  assign n780 = n778 & n779 ;
  assign n781 = n777 & n780 ;
  assign n782 = n775 & n781 ;
  assign n783 = \u2_adr0_cnt_reg[28]/P0001  & n757 ;
  assign n784 = ~n782 & n783 ;
  assign n785 = ~\u2_adr0_cnt_reg[28]/P0001  & n757 ;
  assign n786 = n782 & n785 ;
  assign n787 = ~n784 & ~n786 ;
  assign n788 = \u0_u0_ch_adr0_r_reg[28]/P0001  & ~n757 ;
  assign n789 = n787 & ~n788 ;
  assign n790 = \u2_adr1_cnt_reg[27]/P0001  & n757 ;
  assign n791 = ~n750 & n790 ;
  assign n792 = ~\u2_adr1_cnt_reg[27]/P0001  & n757 ;
  assign n793 = n750 & n792 ;
  assign n794 = ~n791 & ~n793 ;
  assign n795 = \u0_u0_ch_adr1_r_reg[27]/P0001  & ~n757 ;
  assign n796 = n794 & ~n795 ;
  assign n797 = \u0_u0_ch_adr0_r_reg[27]/P0001  & ~n757 ;
  assign n798 = \u2_adr0_cnt_reg[26]/P0001  & n778 ;
  assign n799 = n777 & n798 ;
  assign n800 = n775 & n799 ;
  assign n801 = ~\u2_adr0_cnt_reg[27]/P0001  & ~n800 ;
  assign n802 = n757 & ~n782 ;
  assign n803 = ~n801 & n802 ;
  assign n804 = ~n797 & ~n803 ;
  assign n805 = n746 & n747 ;
  assign n806 = n744 & n805 ;
  assign n807 = ~\u2_adr1_cnt_reg[26]/P0001  & ~n806 ;
  assign n808 = ~n750 & n757 ;
  assign n809 = ~n807 & n808 ;
  assign n810 = \u0_u0_ch_adr1_r_reg[26]/P0001  & ~n757 ;
  assign n811 = ~n809 & ~n810 ;
  assign n812 = n777 & n778 ;
  assign n813 = n775 & n812 ;
  assign n814 = ~\u2_adr0_cnt_reg[26]/P0001  & ~n813 ;
  assign n815 = n757 & ~n800 ;
  assign n816 = ~n814 & n815 ;
  assign n817 = \u0_u0_ch_adr0_r_reg[26]/P0001  & ~n757 ;
  assign n818 = ~n816 & ~n817 ;
  assign n819 = n775 & n777 ;
  assign n820 = ~\u2_adr0_cnt_reg[24]/P0001  & ~n819 ;
  assign n821 = \u2_adr0_cnt_reg[24]/P0001  & n777 ;
  assign n822 = n775 & n821 ;
  assign n823 = n757 & ~n822 ;
  assign n824 = ~n820 & n823 ;
  assign n825 = \u0_u0_ch_adr0_r_reg[24]/P0001  & ~n757 ;
  assign n826 = ~n824 & ~n825 ;
  assign n827 = \u2_adr1_cnt_reg[23]/P0001  & n747 ;
  assign n828 = n744 & n827 ;
  assign n829 = ~\u2_adr1_cnt_reg[24]/P0001  & ~n828 ;
  assign n830 = n745 & n747 ;
  assign n831 = n744 & n830 ;
  assign n832 = n757 & ~n831 ;
  assign n833 = ~n829 & n832 ;
  assign n834 = \u0_u0_ch_adr1_r_reg[24]/P0001  & ~n757 ;
  assign n835 = ~n833 & ~n834 ;
  assign n836 = \u0_u0_ch_adr0_r_reg[23]/P0001  & ~n757 ;
  assign n837 = \u2_adr0_cnt_reg[20]/P0001  & \u2_adr0_cnt_reg[21]/P0001  ;
  assign n838 = n773 & n837 ;
  assign n839 = n770 & n838 ;
  assign n840 = \u2_adr0_cnt_reg[22]/P0001  & n839 ;
  assign n841 = ~\u2_adr0_cnt_reg[23]/P0001  & ~n840 ;
  assign n842 = n757 & ~n819 ;
  assign n843 = ~n841 & n842 ;
  assign n844 = ~n836 & ~n843 ;
  assign n845 = n744 & n747 ;
  assign n846 = ~\u2_adr1_cnt_reg[23]/P0001  & ~n845 ;
  assign n847 = n757 & ~n828 ;
  assign n848 = ~n846 & n847 ;
  assign n849 = \u0_u0_ch_adr1_r_reg[23]/P0001  & ~n757 ;
  assign n850 = ~n848 & ~n849 ;
  assign n851 = ~\u2_adr0_cnt_reg[22]/P0001  & ~n839 ;
  assign n852 = n757 & ~n840 ;
  assign n853 = ~n851 & n852 ;
  assign n854 = \u0_u0_ch_adr0_r_reg[22]/P0001  & ~n757 ;
  assign n855 = ~n853 & ~n854 ;
  assign n856 = \u0_u0_ch_adr1_r_reg[22]/P0001  & ~n757 ;
  assign n857 = \u2_adr1_cnt_reg[21]/P0001  & n744 ;
  assign n858 = ~\u2_adr1_cnt_reg[22]/P0001  & ~n857 ;
  assign n859 = n757 & ~n845 ;
  assign n860 = ~n858 & n859 ;
  assign n861 = ~n856 & ~n860 ;
  assign n862 = n770 & n773 ;
  assign n863 = ~\u2_adr0_cnt_reg[20]/P0001  & ~n862 ;
  assign n864 = n757 & ~n775 ;
  assign n865 = ~n863 & n864 ;
  assign n866 = \u0_u0_ch_adr0_r_reg[20]/P0001  & ~n757 ;
  assign n867 = ~n865 & ~n866 ;
  assign n868 = \u0_u0_ch_adr1_r_reg[20]/P0001  & ~n757 ;
  assign n869 = \u2_adr1_cnt_reg[18]/P0001  & \u2_adr1_cnt_reg[19]/P0001  ;
  assign n870 = n740 & n869 ;
  assign n871 = n738 & n870 ;
  assign n872 = ~\u2_adr1_cnt_reg[20]/P0001  & ~n871 ;
  assign n873 = ~n744 & n757 ;
  assign n874 = ~n872 & n873 ;
  assign n875 = ~n868 & ~n874 ;
  assign n876 = \u0_u0_ch_adr0_r_reg[19]/P0001  & ~n757 ;
  assign n877 = \u2_adr0_cnt_reg[16]/NET0131  & \u2_u0_out_r_reg[16]/P0001  ;
  assign n878 = n768 & n877 ;
  assign n879 = ~n767 & n878 ;
  assign n880 = \u2_adr0_cnt_reg[17]/P0001  & \u2_adr0_cnt_reg[18]/P0001  ;
  assign n881 = n879 & n880 ;
  assign n882 = ~\u2_adr0_cnt_reg[19]/P0001  & ~n881 ;
  assign n883 = n757 & ~n862 ;
  assign n884 = ~n882 & n883 ;
  assign n885 = ~n876 & ~n884 ;
  assign n886 = \u2_adr1_cnt_reg[18]/P0001  & n740 ;
  assign n887 = n738 & n886 ;
  assign n888 = ~\u2_adr1_cnt_reg[19]/P0001  & ~n887 ;
  assign n889 = n757 & ~n871 ;
  assign n890 = ~n888 & n889 ;
  assign n891 = \u0_u0_ch_adr1_r_reg[19]/P0001  & ~n757 ;
  assign n892 = ~n890 & ~n891 ;
  assign n893 = \u2_adr0_cnt_reg[17]/P0001  & n879 ;
  assign n894 = ~\u2_adr0_cnt_reg[18]/P0001  & ~n893 ;
  assign n895 = n757 & ~n881 ;
  assign n896 = ~n894 & n895 ;
  assign n897 = \u0_u0_ch_adr0_r_reg[18]/P0001  & ~n757 ;
  assign n898 = ~n896 & ~n897 ;
  assign n899 = n738 & n740 ;
  assign n900 = ~\u2_adr1_cnt_reg[18]/P0001  & ~n899 ;
  assign n901 = n757 & ~n887 ;
  assign n902 = ~n900 & n901 ;
  assign n903 = \u0_u0_ch_adr1_r_reg[18]/P0001  & ~n757 ;
  assign n904 = ~n902 & ~n903 ;
  assign n905 = \u2_adr0_cnt_reg[28]/P0001  & n782 ;
  assign n906 = ~\u2_adr0_cnt_reg[29]/P0001  & n757 ;
  assign n907 = ~n905 & n906 ;
  assign n908 = \u2_adr0_cnt_reg[29]/P0001  & n757 ;
  assign n909 = n905 & n908 ;
  assign n910 = ~n907 & ~n909 ;
  assign n911 = ~\u0_u0_ch_adr0_r_reg[29]/P0001  & ~n757 ;
  assign n912 = n910 & ~n911 ;
  assign n913 = ~\u2_chunk_cnt_reg[6]/NET0131  & ~\u2_chunk_cnt_reg[7]/NET0131  ;
  assign n914 = ~\u2_chunk_cnt_reg[0]/NET0131  & ~\u2_chunk_cnt_reg[1]/NET0131  ;
  assign n915 = ~\u2_chunk_cnt_reg[2]/NET0131  & ~\u2_chunk_cnt_reg[3]/NET0131  ;
  assign n916 = n914 & n915 ;
  assign n917 = n913 & n916 ;
  assign n918 = ~\u2_chunk_cnt_reg[4]/NET0131  & ~\u2_chunk_cnt_reg[5]/NET0131  ;
  assign n919 = ~\u2_chunk_cnt_reg[8]/NET0131  & n918 ;
  assign n920 = ~\u2_chunk_0_reg/P0001  & n919 ;
  assign n921 = n917 & n920 ;
  assign n922 = ~\u0_u0_ch_sz_inf_reg/NET0131  & ~\u2_tsz_cnt_reg[0]/NET0131  ;
  assign n923 = ~\u2_tsz_cnt_reg[10]/NET0131  & ~\u2_tsz_cnt_reg[11]/NET0131  ;
  assign n924 = ~\u2_tsz_cnt_reg[1]/NET0131  & ~\u2_tsz_cnt_reg[2]/NET0131  ;
  assign n925 = n923 & n924 ;
  assign n926 = n922 & n925 ;
  assign n927 = ~\u2_tsz_cnt_reg[7]/NET0131  & ~\u2_tsz_cnt_reg[8]/NET0131  ;
  assign n928 = ~\u2_tsz_cnt_reg[9]/NET0131  & n927 ;
  assign n929 = ~\u2_tsz_cnt_reg[3]/NET0131  & ~\u2_tsz_cnt_reg[4]/NET0131  ;
  assign n930 = ~\u2_tsz_cnt_reg[5]/NET0131  & ~\u2_tsz_cnt_reg[6]/NET0131  ;
  assign n931 = n929 & n930 ;
  assign n932 = n928 & n931 ;
  assign n933 = n926 & n932 ;
  assign n934 = ~n921 & ~n933 ;
  assign n935 = ~\u2_state_reg[1]/NET0131  & \u2_state_reg[2]/NET0131  ;
  assign n936 = ~\u2_dma_abort_r_reg/NET0131  & n935 ;
  assign n937 = ~n736 & n936 ;
  assign n938 = n934 & n937 ;
  assign n939 = \u2_state_reg[1]/NET0131  & ~\u2_state_reg[2]/NET0131  ;
  assign n940 = ~\u2_dma_abort_r_reg/NET0131  & n939 ;
  assign n941 = n767 & n940 ;
  assign n942 = ~n938 & ~n941 ;
  assign n943 = ~\u0_u0_ch_csr_r_reg[2]/NET0131  & ~n942 ;
  assign n944 = n736 & n936 ;
  assign n945 = ~n767 & n940 ;
  assign n946 = ~n944 & ~n945 ;
  assign n947 = ~\u0_u0_ch_csr_r_reg[1]/NET0131  & ~n946 ;
  assign n948 = ~\u2_state_reg[10]/NET0131  & ~\u2_state_reg[8]/NET0131  ;
  assign n949 = ~\u2_state_reg[3]/NET0131  & ~\u2_state_reg[9]/NET0131  ;
  assign n950 = n948 & n949 ;
  assign n951 = ~\u2_state_reg[7]/NET0131  & n950 ;
  assign n952 = ~\u2_state_reg[0]/NET0131  & ~\u2_state_reg[1]/NET0131  ;
  assign n953 = ~\u2_state_reg[2]/NET0131  & n952 ;
  assign n954 = \u2_state_reg[4]/NET0131  & \u2_state_reg[6]/NET0131  ;
  assign n955 = n953 & ~n954 ;
  assign n956 = ~\u2_state_reg[4]/NET0131  & ~\u2_state_reg[6]/NET0131  ;
  assign n957 = ~\u2_state_reg[5]/NET0131  & n956 ;
  assign n958 = \u2_state_reg[5]/NET0131  & ~n956 ;
  assign n959 = ~n957 & ~n958 ;
  assign n960 = n955 & n959 ;
  assign n961 = n951 & n960 ;
  assign n962 = ~\u2_state_reg[7]/NET0131  & ~\u2_state_reg[9]/NET0131  ;
  assign n963 = \u0_u0_ch_csr_r_reg[7]/NET0131  & \u0_u0_ch_csr_r_reg[8]/NET0131  ;
  assign n964 = \u1_ndr_r_reg[0]/NET0131  & \u2_state_reg[3]/NET0131  ;
  assign n965 = n963 & n964 ;
  assign n966 = n962 & n965 ;
  assign n967 = ~\wb0_ack_i_pad  & ~n962 ;
  assign n968 = ~n966 & ~n967 ;
  assign n969 = ~n961 & n968 ;
  assign n970 = ~n947 & n969 ;
  assign n971 = ~n943 & n970 ;
  assign n972 = ~n941 & n946 ;
  assign n973 = ~n938 & n972 ;
  assign n974 = ~\u0_u0_ch_csr_r_reg[1]/NET0131  & \u2_write_hold_r_reg/P0001  ;
  assign n975 = ~n973 & n974 ;
  assign n976 = \u0_u0_ch_csr_r_reg[2]/NET0131  & n969 ;
  assign n977 = n934 & ~n946 ;
  assign n978 = n969 & ~n977 ;
  assign n979 = n942 & n978 ;
  assign n980 = ~n976 & ~n979 ;
  assign n981 = ~n975 & ~n980 ;
  assign n982 = ~n971 & ~n981 ;
  assign n983 = \u2_adr1_cnt_reg[25]/P0001  & \u2_adr1_cnt_reg[26]/P0001  ;
  assign n984 = \u2_adr1_cnt_reg[27]/P0001  & \u2_adr1_cnt_reg[28]/P0001  ;
  assign n985 = n983 & n984 ;
  assign n986 = n831 & n985 ;
  assign n987 = ~\u2_adr1_cnt_reg[29]/P0001  & n757 ;
  assign n988 = ~n986 & n987 ;
  assign n989 = \u2_adr1_cnt_reg[29]/P0001  & n757 ;
  assign n990 = n986 & n989 ;
  assign n991 = ~n988 & ~n990 ;
  assign n992 = ~\u0_u0_ch_adr1_r_reg[29]/P0001  & ~n757 ;
  assign n993 = n991 & ~n992 ;
  assign n994 = \u2_adr1_cnt_reg[0]/P0001  & ~n941 ;
  assign n995 = ~n938 & n994 ;
  assign n996 = n969 & n995 ;
  assign n997 = \u2_adr0_cnt_reg[0]/P0001  & n969 ;
  assign n998 = ~n942 & n997 ;
  assign n999 = ~n996 & ~n998 ;
  assign n1000 = ~n961 & ~n967 ;
  assign n1001 = ~\u2_state_reg[2]/NET0131  & ~\u2_state_reg[3]/NET0131  ;
  assign n1002 = n952 & n1001 ;
  assign n1003 = ~\u2_state_reg[5]/NET0131  & ~\u2_state_reg[7]/NET0131  ;
  assign n1004 = n956 & n1003 ;
  assign n1005 = \u2_state_reg[9]/NET0131  & n948 ;
  assign n1006 = n1004 & n1005 ;
  assign n1007 = n1002 & n1006 ;
  assign n1008 = ~n965 & ~n1007 ;
  assign n1009 = ~\u2_state_reg[1]/NET0131  & ~\u2_state_reg[2]/NET0131  ;
  assign n1010 = n950 & n1009 ;
  assign n1011 = ~\u2_state_reg[0]/NET0131  & ~\u2_state_reg[5]/NET0131  ;
  assign n1012 = \u2_state_reg[7]/NET0131  & n956 ;
  assign n1013 = n1011 & n1012 ;
  assign n1014 = n1010 & n1013 ;
  assign n1015 = \wb0_ack_i_pad  & ~n956 ;
  assign n1016 = \u2_state_reg[5]/NET0131  & ~\wb0_ack_i_pad  ;
  assign n1017 = n956 & n1016 ;
  assign n1018 = ~n1015 & ~n1017 ;
  assign n1019 = ~n1014 & n1018 ;
  assign n1020 = n1008 & ~n1019 ;
  assign n1021 = ~n1000 & n1020 ;
  assign n1022 = n999 & ~n1021 ;
  assign n1023 = \u2_adr1_cnt_reg[1]/P0001  & ~n941 ;
  assign n1024 = ~n938 & n1023 ;
  assign n1025 = n969 & n1024 ;
  assign n1026 = \u2_adr0_cnt_reg[1]/P0001  & n969 ;
  assign n1027 = ~n942 & n1026 ;
  assign n1028 = ~n1025 & ~n1027 ;
  assign n1029 = ~\u2_state_reg[5]/NET0131  & ~\u2_state_reg[6]/NET0131  ;
  assign n1030 = ~\wb0_ack_i_pad  & n956 ;
  assign n1031 = ~n1029 & ~n1030 ;
  assign n1032 = ~n1014 & ~n1031 ;
  assign n1033 = n1008 & ~n1032 ;
  assign n1034 = ~n1000 & n1033 ;
  assign n1035 = n1028 & ~n1034 ;
  assign n1036 = ~n767 & n768 ;
  assign n1037 = \u2_adr0_cnt_reg[0]/P0001  & ~n1036 ;
  assign n1038 = \u2_u0_out_r_reg[0]/P0001  & n768 ;
  assign n1039 = ~n767 & n1038 ;
  assign n1040 = ~n1037 & ~n1039 ;
  assign n1041 = n757 & ~n1040 ;
  assign n1042 = \u0_u0_ch_adr0_r_reg[0]/P0001  & ~n757 ;
  assign n1043 = ~n1041 & ~n1042 ;
  assign n1044 = \u2_adr0_cnt_reg[10]/P0001  & ~n1036 ;
  assign n1045 = \u2_u0_out_r_reg[10]/P0001  & n768 ;
  assign n1046 = ~n767 & n1045 ;
  assign n1047 = ~n1044 & ~n1046 ;
  assign n1048 = n757 & ~n1047 ;
  assign n1049 = \u0_u0_ch_adr0_r_reg[10]/P0001  & ~n757 ;
  assign n1050 = ~n1048 & ~n1049 ;
  assign n1051 = \u2_adr0_cnt_reg[11]/P0001  & ~n1036 ;
  assign n1052 = \u2_u0_out_r_reg[11]/P0001  & n768 ;
  assign n1053 = ~n767 & n1052 ;
  assign n1054 = ~n1051 & ~n1053 ;
  assign n1055 = n757 & ~n1054 ;
  assign n1056 = \u0_u0_ch_adr0_r_reg[11]/P0001  & ~n757 ;
  assign n1057 = ~n1055 & ~n1056 ;
  assign n1058 = \u2_adr0_cnt_reg[12]/P0001  & ~n1036 ;
  assign n1059 = \u2_u0_out_r_reg[12]/P0001  & n768 ;
  assign n1060 = ~n767 & n1059 ;
  assign n1061 = ~n1058 & ~n1060 ;
  assign n1062 = n757 & ~n1061 ;
  assign n1063 = \u0_u0_ch_adr0_r_reg[12]/P0001  & ~n757 ;
  assign n1064 = ~n1062 & ~n1063 ;
  assign n1065 = \u2_adr0_cnt_reg[14]/P0001  & ~n1036 ;
  assign n1066 = \u2_u0_out_r_reg[14]/P0001  & n768 ;
  assign n1067 = ~n767 & n1066 ;
  assign n1068 = ~n1065 & ~n1067 ;
  assign n1069 = n757 & ~n1068 ;
  assign n1070 = \u0_u0_ch_adr0_r_reg[14]/P0001  & ~n757 ;
  assign n1071 = ~n1069 & ~n1070 ;
  assign n1072 = \u2_adr0_cnt_reg[15]/P0001  & ~n1036 ;
  assign n1073 = \u2_u0_out_r_reg[15]/P0001  & n768 ;
  assign n1074 = ~n767 & n1073 ;
  assign n1075 = ~n1072 & ~n1074 ;
  assign n1076 = n757 & ~n1075 ;
  assign n1077 = \u0_u0_ch_adr0_r_reg[15]/P0001  & ~n757 ;
  assign n1078 = ~n1076 & ~n1077 ;
  assign n1079 = ~\u2_adr0_cnt_reg[16]/NET0131  & ~n770 ;
  assign n1080 = ~n879 & ~n1079 ;
  assign n1081 = n757 & n1080 ;
  assign n1082 = \u0_u0_ch_adr0_r_reg[16]/P0001  & ~n757 ;
  assign n1083 = ~n1081 & ~n1082 ;
  assign n1084 = ~\u2_adr0_cnt_reg[17]/P0001  & ~n879 ;
  assign n1085 = n757 & ~n893 ;
  assign n1086 = ~n1084 & n1085 ;
  assign n1087 = \u0_u0_ch_adr0_r_reg[17]/P0001  & ~n757 ;
  assign n1088 = ~n1086 & ~n1087 ;
  assign n1089 = \u2_adr0_cnt_reg[1]/P0001  & ~n1036 ;
  assign n1090 = \u2_u0_out_r_reg[1]/P0001  & n768 ;
  assign n1091 = ~n767 & n1090 ;
  assign n1092 = ~n1089 & ~n1091 ;
  assign n1093 = n757 & ~n1092 ;
  assign n1094 = \u0_u0_ch_adr0_r_reg[1]/P0001  & ~n757 ;
  assign n1095 = ~n1093 & ~n1094 ;
  assign n1096 = ~\u2_adr0_cnt_reg[21]/P0001  & ~n775 ;
  assign n1097 = n757 & ~n839 ;
  assign n1098 = ~n1096 & n1097 ;
  assign n1099 = \u0_u0_ch_adr0_r_reg[21]/P0001  & ~n757 ;
  assign n1100 = ~n1098 & ~n1099 ;
  assign n1101 = \u0_u0_ch_adr0_r_reg[25]/P0001  & ~n757 ;
  assign n1102 = ~\u2_adr0_cnt_reg[25]/P0001  & ~n822 ;
  assign n1103 = n757 & ~n813 ;
  assign n1104 = ~n1102 & n1103 ;
  assign n1105 = ~n1101 & ~n1104 ;
  assign n1106 = \u2_adr0_cnt_reg[2]/P0001  & ~n1036 ;
  assign n1107 = \u2_u0_out_r_reg[2]/P0001  & n768 ;
  assign n1108 = ~n767 & n1107 ;
  assign n1109 = ~n1106 & ~n1108 ;
  assign n1110 = n757 & ~n1109 ;
  assign n1111 = \u0_u0_ch_adr0_r_reg[2]/P0001  & ~n757 ;
  assign n1112 = ~n1110 & ~n1111 ;
  assign n1113 = \u2_adr0_cnt_reg[3]/P0001  & ~n1036 ;
  assign n1114 = \u2_u0_out_r_reg[3]/P0001  & n768 ;
  assign n1115 = ~n767 & n1114 ;
  assign n1116 = ~n1113 & ~n1115 ;
  assign n1117 = n757 & ~n1116 ;
  assign n1118 = \u0_u0_ch_adr0_r_reg[3]/P0001  & ~n757 ;
  assign n1119 = ~n1117 & ~n1118 ;
  assign n1120 = \u2_adr0_cnt_reg[4]/P0001  & ~n1036 ;
  assign n1121 = \u2_u0_out_r_reg[4]/P0001  & n768 ;
  assign n1122 = ~n767 & n1121 ;
  assign n1123 = ~n1120 & ~n1122 ;
  assign n1124 = n757 & ~n1123 ;
  assign n1125 = \u0_u0_ch_adr0_r_reg[4]/P0001  & ~n757 ;
  assign n1126 = ~n1124 & ~n1125 ;
  assign n1127 = \u2_adr0_cnt_reg[5]/P0001  & ~n1036 ;
  assign n1128 = \u2_u0_out_r_reg[5]/P0001  & n768 ;
  assign n1129 = ~n767 & n1128 ;
  assign n1130 = ~n1127 & ~n1129 ;
  assign n1131 = n757 & ~n1130 ;
  assign n1132 = \u0_u0_ch_adr0_r_reg[5]/P0001  & ~n757 ;
  assign n1133 = ~n1131 & ~n1132 ;
  assign n1134 = \u2_adr0_cnt_reg[6]/P0001  & ~n1036 ;
  assign n1135 = \u2_u0_out_r_reg[6]/P0001  & n768 ;
  assign n1136 = ~n767 & n1135 ;
  assign n1137 = ~n1134 & ~n1136 ;
  assign n1138 = n757 & ~n1137 ;
  assign n1139 = \u0_u0_ch_adr0_r_reg[6]/P0001  & ~n757 ;
  assign n1140 = ~n1138 & ~n1139 ;
  assign n1141 = \u2_adr0_cnt_reg[7]/P0001  & ~n1036 ;
  assign n1142 = \u2_u0_out_r_reg[7]/P0001  & n768 ;
  assign n1143 = ~n767 & n1142 ;
  assign n1144 = ~n1141 & ~n1143 ;
  assign n1145 = n757 & ~n1144 ;
  assign n1146 = \u0_u0_ch_adr0_r_reg[7]/P0001  & ~n757 ;
  assign n1147 = ~n1145 & ~n1146 ;
  assign n1148 = \u2_adr0_cnt_reg[8]/P0001  & ~n1036 ;
  assign n1149 = \u2_u0_out_r_reg[8]/P0001  & n768 ;
  assign n1150 = ~n767 & n1149 ;
  assign n1151 = ~n1148 & ~n1150 ;
  assign n1152 = n757 & ~n1151 ;
  assign n1153 = \u0_u0_ch_adr0_r_reg[8]/P0001  & ~n757 ;
  assign n1154 = ~n1152 & ~n1153 ;
  assign n1155 = \u2_adr0_cnt_reg[9]/P0001  & ~n1036 ;
  assign n1156 = \u2_u0_out_r_reg[9]/P0001  & n768 ;
  assign n1157 = ~n767 & n1156 ;
  assign n1158 = ~n1155 & ~n1157 ;
  assign n1159 = n757 & ~n1158 ;
  assign n1160 = \u0_u0_ch_adr0_r_reg[9]/P0001  & ~n757 ;
  assign n1161 = ~n1159 & ~n1160 ;
  assign n1162 = \u0_u0_ch_csr_r_reg[1]/NET0131  & ~n946 ;
  assign n1163 = ~\u0_u0_ch_csr_r_reg[2]/NET0131  & ~n1162 ;
  assign n1164 = ~n941 & ~n1162 ;
  assign n1165 = ~n938 & n1164 ;
  assign n1166 = ~n1163 & ~n1165 ;
  assign n1167 = n942 & ~n977 ;
  assign n1168 = \u0_u0_ch_csr_r_reg[2]/NET0131  & ~n1167 ;
  assign n1169 = \u0_u0_ch_csr_r_reg[1]/NET0131  & \u2_write_hold_r_reg/P0001  ;
  assign n1170 = ~n973 & n1169 ;
  assign n1171 = ~n1168 & ~n1170 ;
  assign n1172 = n1166 & ~n1171 ;
  assign n1173 = \u0_u0_ch_adr1_r_reg[17]/P0001  & ~n757 ;
  assign n1174 = n737 & n739 ;
  assign n1175 = ~n736 & n1174 ;
  assign n1176 = ~\u2_adr1_cnt_reg[17]/P0001  & ~n1175 ;
  assign n1177 = ~n899 & ~n1176 ;
  assign n1178 = n757 & n1177 ;
  assign n1179 = ~n1173 & ~n1178 ;
  assign n1180 = ~\u2_adr1_cnt_reg[21]/P0001  & ~n744 ;
  assign n1181 = n757 & ~n857 ;
  assign n1182 = ~n1180 & n1181 ;
  assign n1183 = \u0_u0_ch_adr1_r_reg[21]/P0001  & ~n757 ;
  assign n1184 = ~n1182 & ~n1183 ;
  assign n1185 = \u2_adr1_cnt_reg[9]/P0001  & ~n941 ;
  assign n1186 = ~n938 & n1185 ;
  assign n1187 = n969 & n1186 ;
  assign n1188 = \u2_adr0_cnt_reg[9]/P0001  & n969 ;
  assign n1189 = ~n942 & n1188 ;
  assign n1190 = ~n1187 & ~n1189 ;
  assign n1191 = \u2_adr1_cnt_reg[10]/P0001  & ~n941 ;
  assign n1192 = ~n938 & n1191 ;
  assign n1193 = n969 & n1192 ;
  assign n1194 = \u2_adr0_cnt_reg[10]/P0001  & n969 ;
  assign n1195 = ~n942 & n1194 ;
  assign n1196 = ~n1193 & ~n1195 ;
  assign n1197 = \u2_adr1_cnt_reg[11]/P0001  & ~n941 ;
  assign n1198 = ~n938 & n1197 ;
  assign n1199 = n969 & n1198 ;
  assign n1200 = \u2_adr0_cnt_reg[11]/P0001  & n969 ;
  assign n1201 = ~n942 & n1200 ;
  assign n1202 = ~n1199 & ~n1201 ;
  assign n1203 = \u2_adr1_cnt_reg[12]/P0001  & ~n941 ;
  assign n1204 = ~n938 & n1203 ;
  assign n1205 = n969 & n1204 ;
  assign n1206 = \u2_adr0_cnt_reg[12]/P0001  & n969 ;
  assign n1207 = ~n942 & n1206 ;
  assign n1208 = ~n1205 & ~n1207 ;
  assign n1209 = \u2_adr1_cnt_reg[13]/P0001  & ~n941 ;
  assign n1210 = ~n938 & n1209 ;
  assign n1211 = n969 & n1210 ;
  assign n1212 = \u2_adr0_cnt_reg[13]/P0001  & n969 ;
  assign n1213 = ~n942 & n1212 ;
  assign n1214 = ~n1211 & ~n1213 ;
  assign n1215 = \u2_adr1_cnt_reg[14]/P0001  & ~n941 ;
  assign n1216 = ~n938 & n1215 ;
  assign n1217 = n969 & n1216 ;
  assign n1218 = \u2_adr0_cnt_reg[14]/P0001  & n969 ;
  assign n1219 = ~n942 & n1218 ;
  assign n1220 = ~n1217 & ~n1219 ;
  assign n1221 = \u2_adr1_cnt_reg[15]/P0001  & ~n941 ;
  assign n1222 = ~n938 & n1221 ;
  assign n1223 = n969 & n1222 ;
  assign n1224 = \u2_adr0_cnt_reg[15]/P0001  & n969 ;
  assign n1225 = ~n942 & n1224 ;
  assign n1226 = ~n1223 & ~n1225 ;
  assign n1227 = \u2_adr1_cnt_reg[16]/NET0131  & ~n941 ;
  assign n1228 = ~n938 & n1227 ;
  assign n1229 = n969 & n1228 ;
  assign n1230 = \u2_adr0_cnt_reg[16]/NET0131  & n969 ;
  assign n1231 = ~n942 & n1230 ;
  assign n1232 = ~n1229 & ~n1231 ;
  assign n1233 = \u2_adr1_cnt_reg[17]/P0001  & ~n941 ;
  assign n1234 = ~n938 & n1233 ;
  assign n1235 = n969 & n1234 ;
  assign n1236 = \u2_adr0_cnt_reg[17]/P0001  & n969 ;
  assign n1237 = ~n942 & n1236 ;
  assign n1238 = ~n1235 & ~n1237 ;
  assign n1239 = \u2_adr1_cnt_reg[18]/P0001  & ~n941 ;
  assign n1240 = ~n938 & n1239 ;
  assign n1241 = n969 & n1240 ;
  assign n1242 = \u2_adr0_cnt_reg[18]/P0001  & n969 ;
  assign n1243 = ~n942 & n1242 ;
  assign n1244 = ~n1241 & ~n1243 ;
  assign n1245 = \u2_adr1_cnt_reg[19]/P0001  & ~n941 ;
  assign n1246 = ~n938 & n1245 ;
  assign n1247 = n969 & n1246 ;
  assign n1248 = \u2_adr0_cnt_reg[19]/P0001  & n969 ;
  assign n1249 = ~n942 & n1248 ;
  assign n1250 = ~n1247 & ~n1249 ;
  assign n1251 = \u2_adr1_cnt_reg[20]/P0001  & ~n941 ;
  assign n1252 = ~n938 & n1251 ;
  assign n1253 = n969 & n1252 ;
  assign n1254 = \u2_adr0_cnt_reg[20]/P0001  & n969 ;
  assign n1255 = ~n942 & n1254 ;
  assign n1256 = ~n1253 & ~n1255 ;
  assign n1257 = \u2_adr1_cnt_reg[21]/P0001  & ~n941 ;
  assign n1258 = ~n938 & n1257 ;
  assign n1259 = n969 & n1258 ;
  assign n1260 = \u2_adr0_cnt_reg[21]/P0001  & n969 ;
  assign n1261 = ~n942 & n1260 ;
  assign n1262 = ~n1259 & ~n1261 ;
  assign n1263 = \u2_adr1_cnt_reg[22]/P0001  & ~n941 ;
  assign n1264 = ~n938 & n1263 ;
  assign n1265 = n969 & n1264 ;
  assign n1266 = \u2_adr0_cnt_reg[22]/P0001  & n969 ;
  assign n1267 = ~n942 & n1266 ;
  assign n1268 = ~n1265 & ~n1267 ;
  assign n1269 = \u2_adr1_cnt_reg[23]/P0001  & ~n941 ;
  assign n1270 = ~n938 & n1269 ;
  assign n1271 = n969 & n1270 ;
  assign n1272 = \u2_adr0_cnt_reg[23]/P0001  & n969 ;
  assign n1273 = ~n942 & n1272 ;
  assign n1274 = ~n1271 & ~n1273 ;
  assign n1275 = \u2_adr1_cnt_reg[24]/P0001  & ~n941 ;
  assign n1276 = ~n938 & n1275 ;
  assign n1277 = n969 & n1276 ;
  assign n1278 = \u2_adr0_cnt_reg[24]/P0001  & n969 ;
  assign n1279 = ~n942 & n1278 ;
  assign n1280 = ~n1277 & ~n1279 ;
  assign n1281 = \u2_adr1_cnt_reg[25]/P0001  & ~n941 ;
  assign n1282 = ~n938 & n1281 ;
  assign n1283 = n969 & n1282 ;
  assign n1284 = \u2_adr0_cnt_reg[25]/P0001  & n969 ;
  assign n1285 = ~n942 & n1284 ;
  assign n1286 = ~n1283 & ~n1285 ;
  assign n1287 = \u2_adr1_cnt_reg[26]/P0001  & ~n941 ;
  assign n1288 = ~n938 & n1287 ;
  assign n1289 = n969 & n1288 ;
  assign n1290 = \u2_adr0_cnt_reg[26]/P0001  & n969 ;
  assign n1291 = ~n942 & n1290 ;
  assign n1292 = ~n1289 & ~n1291 ;
  assign n1293 = \u2_adr1_cnt_reg[27]/P0001  & ~n941 ;
  assign n1294 = ~n938 & n1293 ;
  assign n1295 = n969 & n1294 ;
  assign n1296 = \u2_adr0_cnt_reg[27]/P0001  & n969 ;
  assign n1297 = ~n942 & n1296 ;
  assign n1298 = ~n1295 & ~n1297 ;
  assign n1299 = \u2_adr1_cnt_reg[28]/P0001  & ~n941 ;
  assign n1300 = ~n938 & n1299 ;
  assign n1301 = n969 & n1300 ;
  assign n1302 = \u2_adr0_cnt_reg[28]/P0001  & n969 ;
  assign n1303 = ~n942 & n1302 ;
  assign n1304 = ~n1301 & ~n1303 ;
  assign n1305 = \u2_adr1_cnt_reg[29]/P0001  & ~n941 ;
  assign n1306 = ~n938 & n1305 ;
  assign n1307 = n969 & n1306 ;
  assign n1308 = \u2_adr0_cnt_reg[29]/P0001  & n969 ;
  assign n1309 = ~n942 & n1308 ;
  assign n1310 = ~n1307 & ~n1309 ;
  assign n1311 = \u2_adr1_cnt_reg[8]/P0001  & ~n941 ;
  assign n1312 = ~n938 & n1311 ;
  assign n1313 = n969 & n1312 ;
  assign n1314 = \u2_adr0_cnt_reg[8]/P0001  & n969 ;
  assign n1315 = ~n942 & n1314 ;
  assign n1316 = ~n1313 & ~n1315 ;
  assign n1317 = \u2_adr1_cnt_reg[2]/P0001  & ~n941 ;
  assign n1318 = ~n938 & n1317 ;
  assign n1319 = n969 & n1318 ;
  assign n1320 = \u2_adr0_cnt_reg[2]/P0001  & n969 ;
  assign n1321 = ~n942 & n1320 ;
  assign n1322 = ~n1319 & ~n1321 ;
  assign n1323 = \u2_adr1_cnt_reg[3]/P0001  & ~n941 ;
  assign n1324 = ~n938 & n1323 ;
  assign n1325 = n969 & n1324 ;
  assign n1326 = \u2_adr0_cnt_reg[3]/P0001  & n969 ;
  assign n1327 = ~n942 & n1326 ;
  assign n1328 = ~n1325 & ~n1327 ;
  assign n1329 = \u2_adr1_cnt_reg[4]/P0001  & ~n941 ;
  assign n1330 = ~n938 & n1329 ;
  assign n1331 = n969 & n1330 ;
  assign n1332 = \u2_adr0_cnt_reg[4]/P0001  & n969 ;
  assign n1333 = ~n942 & n1332 ;
  assign n1334 = ~n1331 & ~n1333 ;
  assign n1335 = \u2_adr1_cnt_reg[5]/P0001  & ~n941 ;
  assign n1336 = ~n938 & n1335 ;
  assign n1337 = n969 & n1336 ;
  assign n1338 = \u2_adr0_cnt_reg[5]/P0001  & n969 ;
  assign n1339 = ~n942 & n1338 ;
  assign n1340 = ~n1337 & ~n1339 ;
  assign n1341 = \u2_adr1_cnt_reg[6]/P0001  & ~n941 ;
  assign n1342 = ~n938 & n1341 ;
  assign n1343 = n969 & n1342 ;
  assign n1344 = \u2_adr0_cnt_reg[6]/P0001  & n969 ;
  assign n1345 = ~n942 & n1344 ;
  assign n1346 = ~n1343 & ~n1345 ;
  assign n1347 = \u2_adr1_cnt_reg[7]/P0001  & ~n941 ;
  assign n1348 = ~n938 & n1347 ;
  assign n1349 = n969 & n1348 ;
  assign n1350 = \u2_adr0_cnt_reg[7]/P0001  & n969 ;
  assign n1351 = ~n942 & n1350 ;
  assign n1352 = ~n1349 & ~n1351 ;
  assign n1353 = ~\u3_u1_slv_adr_reg[6]/NET0131  & ~\u3_u1_slv_adr_reg[7]/NET0131  ;
  assign n1354 = ~\u3_u1_slv_adr_reg[8]/NET0131  & ~\u3_u1_slv_adr_reg[9]/NET0131  ;
  assign n1355 = n1353 & n1354 ;
  assign n1356 = ~\u3_u1_slv_adr_reg[2]/NET0131  & ~\u3_u1_slv_adr_reg[3]/P0001  ;
  assign n1357 = \u3_u1_slv_adr_reg[5]/P0001  & n1356 ;
  assign n1358 = n1355 & n1357 ;
  assign n1359 = ~\u3_u1_slv_adr_reg[4]/NET0131  & \u3_u1_slv_we_reg/P0001  ;
  assign n1360 = ~\u3_u1_slv_dout_reg[0]/P0001  & n1359 ;
  assign n1361 = n1358 & n1360 ;
  assign n1362 = n1358 & n1359 ;
  assign n1363 = ~\u0_u0_ch_csr_r_reg[0]/NET0131  & ~n1362 ;
  assign n1364 = ~\u1_ndnr_reg[0]/P0001  & ~\u2_state_reg[3]/NET0131  ;
  assign n1365 = \u1_ndr_r_reg[0]/NET0131  & n919 ;
  assign n1366 = n917 & n1365 ;
  assign n1367 = ~\u1_ndnr_reg[0]/P0001  & ~\u2_tsz_cnt_is_0_r_reg/P0001  ;
  assign n1368 = ~n1366 & n1367 ;
  assign n1369 = ~n1364 & ~n1368 ;
  assign n1370 = ~\u0_u0_ch_csr_r_reg[6]/NET0131  & ~\u0_u0_ch_csr_r_reg[7]/NET0131  ;
  assign n1371 = ~n1362 & n1370 ;
  assign n1372 = n1369 & n1371 ;
  assign n1373 = ~n1363 & ~n1372 ;
  assign n1374 = ~n1361 & n1373 ;
  assign n1375 = n948 & n962 ;
  assign n1376 = ~\u2_state_reg[3]/NET0131  & ~\u2_state_reg[4]/NET0131  ;
  assign n1377 = n1029 & n1376 ;
  assign n1378 = n1375 & n1377 ;
  assign n1379 = ~\u2_state_reg[0]/NET0131  & n1378 ;
  assign n1380 = \u2_state_reg[1]/NET0131  & n736 ;
  assign n1381 = n936 & n1380 ;
  assign n1382 = ~n938 & ~n1381 ;
  assign n1383 = ~n941 & n1382 ;
  assign n1384 = n1379 & ~n1383 ;
  assign n1385 = n957 & n1002 ;
  assign n1386 = ~\u2_state_reg[10]/NET0131  & \u2_state_reg[8]/NET0131  ;
  assign n1387 = n962 & n1386 ;
  assign n1388 = n1385 & n1387 ;
  assign n1389 = ~\u1_next_start_reg/P0001  & ~n755 ;
  assign n1390 = \u0_u0_ch_csr_r_reg[7]/NET0131  & ~\u0_u0_ch_err_reg/NET0131  ;
  assign n1391 = ~n1389 & n1390 ;
  assign n1392 = \u2_state_reg[0]/NET0131  & n1009 ;
  assign n1393 = ~\u0_csr_r_reg[0]/NET0131  & n1392 ;
  assign n1394 = n1378 & n1393 ;
  assign n1395 = \u0_u0_ch_err_reg/NET0131  & ~\u2_state_reg[1]/NET0131  ;
  assign n1396 = ~\u1_next_start_reg/P0001  & ~\u2_state_reg[1]/NET0131  ;
  assign n1397 = ~n755 & n1396 ;
  assign n1398 = ~n1395 & ~n1397 ;
  assign n1399 = n1394 & n1398 ;
  assign n1400 = ~n1391 & n1399 ;
  assign n1401 = ~n1388 & ~n1400 ;
  assign n1402 = ~n1384 & n1401 ;
  assign n1403 = ~\u0_u0_ch_err_reg/NET0131  & ~n1389 ;
  assign n1404 = n1394 & ~n1403 ;
  assign n1405 = \u1_ndr_r_reg[0]/NET0131  & n963 ;
  assign n1406 = n1029 & n1375 ;
  assign n1407 = \u2_state_reg[3]/NET0131  & ~\u2_state_reg[4]/NET0131  ;
  assign n1408 = n953 & n1407 ;
  assign n1409 = n1406 & n1408 ;
  assign n1410 = ~n1405 & n1409 ;
  assign n1411 = \wb0_ack_i_pad  & n1002 ;
  assign n1412 = n1006 & n1411 ;
  assign n1413 = \u2_state_reg[10]/NET0131  & ~\u2_state_reg[8]/NET0131  ;
  assign n1414 = \u0_csr_r_reg[0]/NET0131  & ~\u2_state_reg[0]/NET0131  ;
  assign n1415 = n962 & ~n1414 ;
  assign n1416 = n1413 & n1415 ;
  assign n1417 = n1385 & n1416 ;
  assign n1418 = ~n1412 & ~n1417 ;
  assign n1419 = ~n1410 & n1418 ;
  assign n1420 = ~n1404 & n1419 ;
  assign n1421 = n1369 & n1370 ;
  assign n1422 = ~\u3_u1_slv_adr_reg[3]/P0001  & ~\u3_u1_slv_adr_reg[4]/NET0131  ;
  assign n1423 = \u3_u1_slv_adr_reg[5]/P0001  & n1422 ;
  assign n1424 = n1355 & n1423 ;
  assign n1425 = ~\u3_u1_slv_adr_reg[2]/NET0131  & \u3_u1_slv_re_reg/P0001  ;
  assign n1426 = n1424 & n1425 ;
  assign n1427 = \u0_u0_int_src_r_reg[1]/NET0131  & ~n1426 ;
  assign n1428 = ~n1421 & ~n1427 ;
  assign n1429 = \u0_u0_ch_adr1_r_reg[16]/P0001  & ~n757 ;
  assign n1430 = \u2_u1_out_r_reg[16]/P0001  & n737 ;
  assign n1431 = ~n736 & n1430 ;
  assign n1432 = ~\u2_adr1_cnt_reg[16]/NET0131  & ~n1431 ;
  assign n1433 = ~n1175 & ~n1432 ;
  assign n1434 = n757 & n1433 ;
  assign n1435 = ~n1429 & ~n1434 ;
  assign n1436 = ~\u2_read_r_reg/P0001  & ~n942 ;
  assign n1437 = \u2_dma_abort_r_reg/NET0131  & n939 ;
  assign n1438 = \u2_state_reg[3]/NET0131  & n939 ;
  assign n1439 = n767 & n1438 ;
  assign n1440 = ~n1437 & ~n1439 ;
  assign n1441 = n1379 & ~n1440 ;
  assign n1442 = ~\u2_state_reg[3]/NET0131  & n736 ;
  assign n1443 = ~\u2_dma_abort_r_reg/NET0131  & n1442 ;
  assign n1444 = ~\u2_dma_abort_r_reg/NET0131  & ~n736 ;
  assign n1445 = n934 & n1444 ;
  assign n1446 = ~n1443 & ~n1445 ;
  assign n1447 = n935 & n1379 ;
  assign n1448 = n1446 & n1447 ;
  assign n1449 = ~n1441 & ~n1448 ;
  assign n1450 = \u2_adr0_cnt_reg[9]/P0001  & ~n942 ;
  assign n1451 = ~n1186 & ~n1450 ;
  assign n1452 = \u2_adr0_cnt_reg[8]/P0001  & ~n942 ;
  assign n1453 = ~n1312 & ~n1452 ;
  assign n1454 = \u2_adr0_cnt_reg[10]/P0001  & ~n942 ;
  assign n1455 = ~n1192 & ~n1454 ;
  assign n1456 = \u2_adr0_cnt_reg[11]/P0001  & ~n942 ;
  assign n1457 = ~n1198 & ~n1456 ;
  assign n1458 = \u2_adr0_cnt_reg[12]/P0001  & ~n942 ;
  assign n1459 = ~n1204 & ~n1458 ;
  assign n1460 = \u2_adr0_cnt_reg[13]/P0001  & ~n942 ;
  assign n1461 = ~n1210 & ~n1460 ;
  assign n1462 = \u2_adr0_cnt_reg[14]/P0001  & ~n942 ;
  assign n1463 = ~n1216 & ~n1462 ;
  assign n1464 = \u2_adr0_cnt_reg[15]/P0001  & ~n942 ;
  assign n1465 = ~n1222 & ~n1464 ;
  assign n1466 = \u2_adr0_cnt_reg[16]/NET0131  & ~n942 ;
  assign n1467 = ~n1228 & ~n1466 ;
  assign n1468 = \u2_adr0_cnt_reg[17]/P0001  & ~n942 ;
  assign n1469 = ~n1234 & ~n1468 ;
  assign n1470 = \u2_adr0_cnt_reg[18]/P0001  & ~n942 ;
  assign n1471 = ~n1240 & ~n1470 ;
  assign n1472 = \u2_adr0_cnt_reg[19]/P0001  & ~n942 ;
  assign n1473 = ~n1246 & ~n1472 ;
  assign n1474 = \u2_adr0_cnt_reg[20]/P0001  & ~n942 ;
  assign n1475 = ~n1252 & ~n1474 ;
  assign n1476 = \u2_adr0_cnt_reg[21]/P0001  & ~n942 ;
  assign n1477 = ~n1258 & ~n1476 ;
  assign n1478 = \u2_adr0_cnt_reg[22]/P0001  & ~n942 ;
  assign n1479 = ~n1264 & ~n1478 ;
  assign n1480 = \u2_adr0_cnt_reg[23]/P0001  & ~n942 ;
  assign n1481 = ~n1270 & ~n1480 ;
  assign n1482 = \u2_adr0_cnt_reg[24]/P0001  & ~n942 ;
  assign n1483 = ~n1276 & ~n1482 ;
  assign n1484 = \u2_adr0_cnt_reg[25]/P0001  & ~n942 ;
  assign n1485 = ~n1282 & ~n1484 ;
  assign n1486 = \u2_adr0_cnt_reg[26]/P0001  & ~n942 ;
  assign n1487 = ~n1288 & ~n1486 ;
  assign n1488 = \u2_adr0_cnt_reg[27]/P0001  & ~n942 ;
  assign n1489 = ~n1294 & ~n1488 ;
  assign n1490 = \u2_adr0_cnt_reg[0]/P0001  & ~n942 ;
  assign n1491 = ~n995 & ~n1490 ;
  assign n1492 = \u2_adr0_cnt_reg[28]/P0001  & ~n942 ;
  assign n1493 = ~n1300 & ~n1492 ;
  assign n1494 = \u2_adr0_cnt_reg[29]/P0001  & ~n942 ;
  assign n1495 = ~n1306 & ~n1494 ;
  assign n1496 = \u2_adr0_cnt_reg[1]/P0001  & ~n942 ;
  assign n1497 = ~n1024 & ~n1496 ;
  assign n1498 = \u2_adr0_cnt_reg[2]/P0001  & ~n942 ;
  assign n1499 = ~n1318 & ~n1498 ;
  assign n1500 = \u2_adr0_cnt_reg[3]/P0001  & ~n942 ;
  assign n1501 = ~n1324 & ~n1500 ;
  assign n1502 = \u2_adr0_cnt_reg[4]/P0001  & ~n942 ;
  assign n1503 = ~n1330 & ~n1502 ;
  assign n1504 = \u2_adr0_cnt_reg[5]/P0001  & ~n942 ;
  assign n1505 = ~n1336 & ~n1504 ;
  assign n1506 = \u2_adr0_cnt_reg[6]/P0001  & ~n942 ;
  assign n1507 = ~n1342 & ~n1506 ;
  assign n1508 = \u2_adr0_cnt_reg[7]/P0001  & ~n942 ;
  assign n1509 = ~n1348 & ~n1508 ;
  assign n1510 = n1405 & n1409 ;
  assign n1511 = n1009 & n1011 ;
  assign n1512 = \u2_state_reg[6]/NET0131  & n1376 ;
  assign n1513 = n1375 & n1512 ;
  assign n1514 = n1511 & n1513 ;
  assign n1515 = ~n1007 & ~n1514 ;
  assign n1516 = \u2_state_reg[9]/NET0131  & ~\wb0_ack_i_pad  ;
  assign n1517 = ~n1515 & n1516 ;
  assign n1518 = ~n1510 & ~n1517 ;
  assign n1519 = \u2_adr1_cnt_reg[2]/P0001  & ~n738 ;
  assign n1520 = \u2_u1_out_r_reg[2]/P0001  & n737 ;
  assign n1521 = ~n736 & n1520 ;
  assign n1522 = ~n1519 & ~n1521 ;
  assign n1523 = n757 & ~n1522 ;
  assign n1524 = \u0_u0_ch_adr1_r_reg[2]/P0001  & ~n757 ;
  assign n1525 = ~n1523 & ~n1524 ;
  assign n1526 = \u2_adr1_cnt_reg[3]/P0001  & ~n738 ;
  assign n1527 = \u2_u1_out_r_reg[3]/P0001  & n737 ;
  assign n1528 = ~n736 & n1527 ;
  assign n1529 = ~n1526 & ~n1528 ;
  assign n1530 = n757 & ~n1529 ;
  assign n1531 = \u0_u0_ch_adr1_r_reg[3]/P0001  & ~n757 ;
  assign n1532 = ~n1530 & ~n1531 ;
  assign n1533 = \u2_adr1_cnt_reg[4]/P0001  & ~n738 ;
  assign n1534 = \u2_u1_out_r_reg[4]/P0001  & n737 ;
  assign n1535 = ~n736 & n1534 ;
  assign n1536 = ~n1533 & ~n1535 ;
  assign n1537 = n757 & ~n1536 ;
  assign n1538 = \u0_u0_ch_adr1_r_reg[4]/P0001  & ~n757 ;
  assign n1539 = ~n1537 & ~n1538 ;
  assign n1540 = \u2_adr1_cnt_reg[5]/P0001  & ~n738 ;
  assign n1541 = \u2_u1_out_r_reg[5]/P0001  & n737 ;
  assign n1542 = ~n736 & n1541 ;
  assign n1543 = ~n1540 & ~n1542 ;
  assign n1544 = n757 & ~n1543 ;
  assign n1545 = \u0_u0_ch_adr1_r_reg[5]/P0001  & ~n757 ;
  assign n1546 = ~n1544 & ~n1545 ;
  assign n1547 = \u2_adr1_cnt_reg[6]/P0001  & ~n738 ;
  assign n1548 = \u2_u1_out_r_reg[6]/P0001  & n737 ;
  assign n1549 = ~n736 & n1548 ;
  assign n1550 = ~n1547 & ~n1549 ;
  assign n1551 = n757 & ~n1550 ;
  assign n1552 = \u0_u0_ch_adr1_r_reg[6]/P0001  & ~n757 ;
  assign n1553 = ~n1551 & ~n1552 ;
  assign n1554 = \u2_adr1_cnt_reg[7]/P0001  & ~n738 ;
  assign n1555 = \u2_u1_out_r_reg[7]/P0001  & n737 ;
  assign n1556 = ~n736 & n1555 ;
  assign n1557 = ~n1554 & ~n1556 ;
  assign n1558 = n757 & ~n1557 ;
  assign n1559 = \u0_u0_ch_adr1_r_reg[7]/P0001  & ~n757 ;
  assign n1560 = ~n1558 & ~n1559 ;
  assign n1561 = \u2_adr1_cnt_reg[8]/P0001  & ~n738 ;
  assign n1562 = \u2_u1_out_r_reg[8]/P0001  & n737 ;
  assign n1563 = ~n736 & n1562 ;
  assign n1564 = ~n1561 & ~n1563 ;
  assign n1565 = n757 & ~n1564 ;
  assign n1566 = \u0_u0_ch_adr1_r_reg[8]/P0001  & ~n757 ;
  assign n1567 = ~n1565 & ~n1566 ;
  assign n1568 = \u2_adr1_cnt_reg[9]/P0001  & ~n738 ;
  assign n1569 = \u2_u1_out_r_reg[9]/P0001  & n737 ;
  assign n1570 = ~n736 & n1569 ;
  assign n1571 = ~n1568 & ~n1570 ;
  assign n1572 = n757 & ~n1571 ;
  assign n1573 = \u0_u0_ch_adr1_r_reg[9]/P0001  & ~n757 ;
  assign n1574 = ~n1572 & ~n1573 ;
  assign n1575 = \u2_adr1_cnt_reg[0]/P0001  & ~n738 ;
  assign n1576 = \u2_u1_out_r_reg[0]/P0001  & n737 ;
  assign n1577 = ~n736 & n1576 ;
  assign n1578 = ~n1575 & ~n1577 ;
  assign n1579 = n757 & ~n1578 ;
  assign n1580 = \u0_u0_ch_adr1_r_reg[0]/P0001  & ~n757 ;
  assign n1581 = ~n1579 & ~n1580 ;
  assign n1582 = \u2_adr1_cnt_reg[10]/P0001  & ~n738 ;
  assign n1583 = \u2_u1_out_r_reg[10]/P0001  & n737 ;
  assign n1584 = ~n736 & n1583 ;
  assign n1585 = ~n1582 & ~n1584 ;
  assign n1586 = n757 & ~n1585 ;
  assign n1587 = \u0_u0_ch_adr1_r_reg[10]/P0001  & ~n757 ;
  assign n1588 = ~n1586 & ~n1587 ;
  assign n1589 = \u2_adr1_cnt_reg[11]/P0001  & ~n738 ;
  assign n1590 = \u2_u1_out_r_reg[11]/P0001  & n737 ;
  assign n1591 = ~n736 & n1590 ;
  assign n1592 = ~n1589 & ~n1591 ;
  assign n1593 = n757 & ~n1592 ;
  assign n1594 = \u0_u0_ch_adr1_r_reg[11]/P0001  & ~n757 ;
  assign n1595 = ~n1593 & ~n1594 ;
  assign n1596 = \u2_adr1_cnt_reg[12]/P0001  & ~n738 ;
  assign n1597 = \u2_u1_out_r_reg[12]/P0001  & n737 ;
  assign n1598 = ~n736 & n1597 ;
  assign n1599 = ~n1596 & ~n1598 ;
  assign n1600 = n757 & ~n1599 ;
  assign n1601 = \u0_u0_ch_adr1_r_reg[12]/P0001  & ~n757 ;
  assign n1602 = ~n1600 & ~n1601 ;
  assign n1603 = \u2_adr1_cnt_reg[13]/P0001  & ~n738 ;
  assign n1604 = \u2_u1_out_r_reg[13]/P0001  & n737 ;
  assign n1605 = ~n736 & n1604 ;
  assign n1606 = ~n1603 & ~n1605 ;
  assign n1607 = n757 & ~n1606 ;
  assign n1608 = \u0_u0_ch_adr1_r_reg[13]/P0001  & ~n757 ;
  assign n1609 = ~n1607 & ~n1608 ;
  assign n1610 = \u2_adr1_cnt_reg[14]/P0001  & ~n738 ;
  assign n1611 = \u2_u1_out_r_reg[14]/P0001  & n737 ;
  assign n1612 = ~n736 & n1611 ;
  assign n1613 = ~n1610 & ~n1612 ;
  assign n1614 = n757 & ~n1613 ;
  assign n1615 = \u0_u0_ch_adr1_r_reg[14]/P0001  & ~n757 ;
  assign n1616 = ~n1614 & ~n1615 ;
  assign n1617 = \u2_adr1_cnt_reg[15]/P0001  & ~n738 ;
  assign n1618 = \u2_u1_out_r_reg[15]/P0001  & n737 ;
  assign n1619 = ~n736 & n1618 ;
  assign n1620 = ~n1617 & ~n1619 ;
  assign n1621 = n757 & ~n1620 ;
  assign n1622 = \u0_u0_ch_adr1_r_reg[15]/P0001  & ~n757 ;
  assign n1623 = ~n1621 & ~n1622 ;
  assign n1624 = \u2_adr1_cnt_reg[1]/P0001  & ~n738 ;
  assign n1625 = \u2_u1_out_r_reg[1]/P0001  & n737 ;
  assign n1626 = ~n736 & n1625 ;
  assign n1627 = ~n1624 & ~n1626 ;
  assign n1628 = n757 & ~n1627 ;
  assign n1629 = \u0_u0_ch_adr1_r_reg[1]/P0001  & ~n757 ;
  assign n1630 = ~n1628 & ~n1629 ;
  assign n1631 = \u0_u0_ch_csr_r_reg[0]/NET0131  & \u2_next_ch_reg/P0001  ;
  assign n1632 = ~n753 & n1631 ;
  assign n1633 = \u0_u0_ch_csr_r_reg[5]/NET0131  & \u2_state_reg[3]/NET0131  ;
  assign n1634 = ~n934 & n1633 ;
  assign n1635 = \u2_state_reg[3]/NET0131  & ~n934 ;
  assign n1636 = \u0_u0_int_src_r_reg[2]/NET0131  & ~n1426 ;
  assign n1637 = ~n1635 & ~n1636 ;
  assign n1638 = n1378 & n1392 ;
  assign n1639 = n962 & n1413 ;
  assign n1640 = n1385 & n1639 ;
  assign n1641 = ~n1638 & ~n1640 ;
  assign n1642 = \u0_csr_r_reg[0]/NET0131  & ~n1641 ;
  assign n1643 = \u2_state_reg[10]/NET0131  & n1392 ;
  assign n1644 = n1378 & n1643 ;
  assign n1645 = ~n1403 & n1644 ;
  assign n1646 = ~n1642 & ~n1645 ;
  assign n1647 = \u0_u0_ch_err_reg/NET0131  & \u2_state_reg[4]/NET0131  ;
  assign n1648 = ~\u1_next_start_reg/P0001  & \u2_state_reg[4]/NET0131  ;
  assign n1649 = ~n755 & n1648 ;
  assign n1650 = ~n1647 & ~n1649 ;
  assign n1651 = ~n1391 & n1650 ;
  assign n1652 = n1394 & ~n1651 ;
  assign n1653 = ~\u2_state_reg[3]/NET0131  & \u2_state_reg[4]/NET0131  ;
  assign n1654 = n953 & n1653 ;
  assign n1655 = n1406 & n1654 ;
  assign n1656 = n1515 & ~n1655 ;
  assign n1657 = \u2_state_reg[4]/NET0131  & ~\wb0_ack_i_pad  ;
  assign n1658 = ~n1656 & n1657 ;
  assign n1659 = ~n1652 & ~n1658 ;
  assign n1660 = ~n946 & n1379 ;
  assign n1661 = \u0_u0_ch_tot_sz_r_reg[10]/P0001  & ~n757 ;
  assign n1662 = \u2_chunk_dec_reg/P0001  & ~\u2_tsz_cnt_is_0_r_reg/P0001  ;
  assign n1663 = ~\u2_tsz_cnt_reg[0]/NET0131  & ~\u2_tsz_cnt_reg[1]/NET0131  ;
  assign n1664 = n1662 & n1663 ;
  assign n1665 = ~\u2_tsz_cnt_reg[2]/NET0131  & ~\u2_tsz_cnt_reg[4]/NET0131  ;
  assign n1666 = ~\u2_tsz_cnt_reg[3]/NET0131  & n1665 ;
  assign n1667 = n1664 & n1666 ;
  assign n1668 = n928 & n930 ;
  assign n1669 = n1667 & n1668 ;
  assign n1670 = ~\u2_tsz_cnt_reg[10]/NET0131  & n1669 ;
  assign n1671 = \u2_tsz_cnt_reg[10]/NET0131  & ~n1669 ;
  assign n1672 = ~n1670 & ~n1671 ;
  assign n1673 = n757 & ~n1672 ;
  assign n1674 = ~n1661 & ~n1673 ;
  assign n1675 = ~\u2_tsz_cnt_reg[11]/NET0131  & n757 ;
  assign n1676 = ~n1670 & n1675 ;
  assign n1677 = \u2_tsz_cnt_reg[11]/NET0131  & n757 ;
  assign n1678 = n1670 & n1677 ;
  assign n1679 = ~n1676 & ~n1678 ;
  assign n1680 = ~\u0_u0_ch_tot_sz_r_reg[11]/P0001  & ~n757 ;
  assign n1681 = n1679 & ~n1680 ;
  assign n1682 = ~\u2_tsz_cnt_reg[0]/NET0131  & n1662 ;
  assign n1683 = \u2_tsz_cnt_reg[1]/NET0131  & ~n1682 ;
  assign n1684 = ~n1664 & ~n1683 ;
  assign n1685 = n757 & ~n1684 ;
  assign n1686 = \u0_u0_ch_tot_sz_r_reg[1]/P0001  & ~n757 ;
  assign n1687 = ~n1685 & ~n1686 ;
  assign n1688 = \u0_u0_ch_tot_sz_r_reg[3]/P0001  & ~n757 ;
  assign n1689 = ~\u2_tsz_cnt_reg[2]/NET0131  & ~\u2_tsz_cnt_reg[3]/NET0131  ;
  assign n1690 = n1664 & n1689 ;
  assign n1691 = ~\u2_tsz_cnt_reg[2]/NET0131  & n1664 ;
  assign n1692 = \u2_tsz_cnt_reg[3]/NET0131  & ~n1691 ;
  assign n1693 = ~n1690 & ~n1692 ;
  assign n1694 = n757 & ~n1693 ;
  assign n1695 = ~n1688 & ~n1694 ;
  assign n1696 = ~\u0_u0_ch_tot_sz_r_reg[9]/P0001  & ~n757 ;
  assign n1697 = n927 & n930 ;
  assign n1698 = n1667 & n1697 ;
  assign n1699 = \u2_tsz_cnt_reg[9]/NET0131  & ~n1698 ;
  assign n1700 = n757 & ~n1669 ;
  assign n1701 = ~n1699 & n1700 ;
  assign n1702 = ~n1696 & ~n1701 ;
  assign n1703 = ~\u2_tsz_cnt_reg[5]/NET0131  & n1667 ;
  assign n1704 = \u2_tsz_cnt_reg[5]/NET0131  & ~n1667 ;
  assign n1705 = ~n1703 & ~n1704 ;
  assign n1706 = n757 & ~n1705 ;
  assign n1707 = \u0_u0_ch_tot_sz_r_reg[5]/P0001  & ~n757 ;
  assign n1708 = ~n1706 & ~n1707 ;
  assign n1709 = \u0_u0_ch_tot_sz_r_reg[6]/P0001  & ~n757 ;
  assign n1710 = n930 & n1667 ;
  assign n1711 = \u2_tsz_cnt_reg[6]/NET0131  & ~n1703 ;
  assign n1712 = ~n1710 & ~n1711 ;
  assign n1713 = n757 & ~n1712 ;
  assign n1714 = ~n1709 & ~n1713 ;
  assign n1715 = ~\u2_tsz_cnt_reg[5]/NET0131  & ~\u2_tsz_cnt_reg[7]/NET0131  ;
  assign n1716 = ~\u2_tsz_cnt_reg[6]/NET0131  & n1715 ;
  assign n1717 = n1667 & n1716 ;
  assign n1718 = \u2_tsz_cnt_reg[7]/NET0131  & ~n1710 ;
  assign n1719 = ~n1717 & ~n1718 ;
  assign n1720 = n757 & ~n1719 ;
  assign n1721 = \u0_u0_ch_tot_sz_r_reg[7]/P0001  & ~n757 ;
  assign n1722 = ~n1720 & ~n1721 ;
  assign n1723 = \u0_u0_ch_tot_sz_r_reg[0]/P0001  & ~n757 ;
  assign n1724 = \u2_tsz_cnt_reg[0]/NET0131  & ~n1662 ;
  assign n1725 = ~n1682 & ~n1724 ;
  assign n1726 = n757 & ~n1725 ;
  assign n1727 = ~n1723 & ~n1726 ;
  assign n1728 = \u0_u0_ch_tot_sz_r_reg[4]/P0001  & ~n757 ;
  assign n1729 = \u2_tsz_cnt_reg[4]/NET0131  & ~n1690 ;
  assign n1730 = ~n1667 & ~n1729 ;
  assign n1731 = n757 & ~n1730 ;
  assign n1732 = ~n1728 & ~n1731 ;
  assign n1733 = ~\u0_u0_ch_tot_sz_r_reg[8]/P0001  & ~n757 ;
  assign n1734 = \u2_tsz_cnt_reg[8]/NET0131  & ~n1717 ;
  assign n1735 = n757 & ~n1698 ;
  assign n1736 = ~n1734 & n1735 ;
  assign n1737 = ~n1733 & ~n1736 ;
  assign n1738 = ~\u2_chunk_cnt_is_0_r_reg/P0001  & \u2_chunk_dec_reg/P0001  ;
  assign n1739 = n914 & n1738 ;
  assign n1740 = ~\u2_chunk_cnt_reg[2]/NET0131  & ~\u2_chunk_cnt_reg[4]/NET0131  ;
  assign n1741 = ~\u2_chunk_cnt_reg[3]/NET0131  & n1740 ;
  assign n1742 = n1739 & n1741 ;
  assign n1743 = ~\u2_chunk_cnt_reg[5]/NET0131  & n913 ;
  assign n1744 = n1742 & n1743 ;
  assign n1745 = ~\u1_next_start_reg/P0001  & \u2_chunk_cnt_reg[8]/NET0131  ;
  assign n1746 = ~n755 & n1745 ;
  assign n1747 = ~n1744 & n1746 ;
  assign n1748 = ~\u1_next_start_reg/P0001  & ~\u2_chunk_cnt_reg[8]/NET0131  ;
  assign n1749 = ~n755 & n1748 ;
  assign n1750 = n1744 & n1749 ;
  assign n1751 = ~n1747 & ~n1750 ;
  assign n1752 = \u0_u0_ch_chk_sz_r_reg[8]/P0001  & ~n1389 ;
  assign n1753 = n1751 & ~n1752 ;
  assign n1754 = \u3_u1_slv_adr_reg[5]/P0001  & n1359 ;
  assign n1755 = n1355 & n1754 ;
  assign n1756 = \u3_u1_slv_adr_reg[2]/NET0131  & ~\u3_u1_slv_adr_reg[3]/P0001  ;
  assign n1757 = n1755 & n1756 ;
  assign n1758 = ~n1407 & ~n1653 ;
  assign n1759 = n1511 & ~n1758 ;
  assign n1760 = n1406 & n1759 ;
  assign n1761 = \u2_mast0_drdy_r_reg/P0001  & \u2_state_reg[5]/NET0131  ;
  assign n1762 = \u0_u0_ch_tot_sz_r_reg[0]/P0001  & ~n1761 ;
  assign n1763 = ~n1760 & n1762 ;
  assign n1764 = ~n1757 & n1763 ;
  assign n1765 = ~n1760 & ~n1761 ;
  assign n1766 = \u3_u0_mast_dout_reg[0]/P0001  & ~n1004 ;
  assign n1767 = \u2_tsz_cnt_reg[0]/NET0131  & n1004 ;
  assign n1768 = ~n1766 & ~n1767 ;
  assign n1769 = ~n1757 & ~n1768 ;
  assign n1770 = ~n1765 & n1769 ;
  assign n1771 = ~n1764 & ~n1770 ;
  assign n1772 = \u3_u1_slv_dout_reg[0]/P0001  & n1756 ;
  assign n1773 = n1755 & n1772 ;
  assign n1774 = n1771 & ~n1773 ;
  assign n1775 = \u0_u0_ch_tot_sz_r_reg[1]/P0001  & ~n1761 ;
  assign n1776 = ~n1760 & n1775 ;
  assign n1777 = ~n1757 & n1776 ;
  assign n1778 = \u3_u0_mast_dout_reg[1]/P0001  & ~n1004 ;
  assign n1779 = \u2_tsz_cnt_reg[1]/NET0131  & n1004 ;
  assign n1780 = ~n1778 & ~n1779 ;
  assign n1781 = ~n1757 & ~n1780 ;
  assign n1782 = ~n1765 & n1781 ;
  assign n1783 = ~n1777 & ~n1782 ;
  assign n1784 = \u3_u1_slv_dout_reg[1]/P0001  & n1756 ;
  assign n1785 = n1755 & n1784 ;
  assign n1786 = n1783 & ~n1785 ;
  assign n1787 = \u2_tsz_cnt_reg[10]/NET0131  & n1004 ;
  assign n1788 = \u3_u0_mast_dout_reg[10]/P0001  & ~n1004 ;
  assign n1789 = ~n1787 & ~n1788 ;
  assign n1790 = ~n1757 & ~n1789 ;
  assign n1791 = ~n1765 & n1790 ;
  assign n1792 = \u3_u1_slv_dout_reg[10]/P0001  & n1756 ;
  assign n1793 = n1755 & n1792 ;
  assign n1794 = \u0_u0_ch_tot_sz_r_reg[10]/P0001  & ~n1757 ;
  assign n1795 = n1765 & n1794 ;
  assign n1796 = ~n1793 & ~n1795 ;
  assign n1797 = ~n1791 & n1796 ;
  assign n1798 = \u2_tsz_cnt_reg[11]/NET0131  & n1004 ;
  assign n1799 = \u3_u0_mast_dout_reg[11]/P0001  & ~n1004 ;
  assign n1800 = ~n1798 & ~n1799 ;
  assign n1801 = ~n1757 & ~n1800 ;
  assign n1802 = ~n1765 & n1801 ;
  assign n1803 = \u3_u1_slv_dout_reg[11]/P0001  & n1756 ;
  assign n1804 = n1755 & n1803 ;
  assign n1805 = \u0_u0_ch_tot_sz_r_reg[11]/P0001  & ~n1757 ;
  assign n1806 = n1765 & n1805 ;
  assign n1807 = ~n1804 & ~n1806 ;
  assign n1808 = ~n1802 & n1807 ;
  assign n1809 = \u2_tsz_cnt_reg[2]/NET0131  & n1004 ;
  assign n1810 = \u3_u0_mast_dout_reg[2]/P0001  & ~n1004 ;
  assign n1811 = ~n1809 & ~n1810 ;
  assign n1812 = ~n1757 & ~n1811 ;
  assign n1813 = ~n1765 & n1812 ;
  assign n1814 = \u3_u1_slv_dout_reg[2]/P0001  & n1756 ;
  assign n1815 = n1755 & n1814 ;
  assign n1816 = \u0_u0_ch_tot_sz_r_reg[2]/P0001  & ~n1757 ;
  assign n1817 = n1765 & n1816 ;
  assign n1818 = ~n1815 & ~n1817 ;
  assign n1819 = ~n1813 & n1818 ;
  assign n1820 = \u2_tsz_cnt_reg[3]/NET0131  & n1004 ;
  assign n1821 = \u3_u0_mast_dout_reg[3]/P0001  & ~n1004 ;
  assign n1822 = ~n1820 & ~n1821 ;
  assign n1823 = ~n1757 & ~n1822 ;
  assign n1824 = ~n1765 & n1823 ;
  assign n1825 = \u3_u1_slv_dout_reg[3]/P0001  & n1756 ;
  assign n1826 = n1755 & n1825 ;
  assign n1827 = \u0_u0_ch_tot_sz_r_reg[3]/P0001  & ~n1757 ;
  assign n1828 = n1765 & n1827 ;
  assign n1829 = ~n1826 & ~n1828 ;
  assign n1830 = ~n1824 & n1829 ;
  assign n1831 = \u2_tsz_cnt_reg[4]/NET0131  & n1004 ;
  assign n1832 = \u3_u0_mast_dout_reg[4]/P0001  & ~n1004 ;
  assign n1833 = ~n1831 & ~n1832 ;
  assign n1834 = ~n1757 & ~n1833 ;
  assign n1835 = ~n1765 & n1834 ;
  assign n1836 = \u3_u1_slv_dout_reg[4]/P0001  & n1756 ;
  assign n1837 = n1755 & n1836 ;
  assign n1838 = \u0_u0_ch_tot_sz_r_reg[4]/P0001  & ~n1757 ;
  assign n1839 = n1765 & n1838 ;
  assign n1840 = ~n1837 & ~n1839 ;
  assign n1841 = ~n1835 & n1840 ;
  assign n1842 = \u2_tsz_cnt_reg[5]/NET0131  & n1004 ;
  assign n1843 = \u3_u0_mast_dout_reg[5]/P0001  & ~n1004 ;
  assign n1844 = ~n1842 & ~n1843 ;
  assign n1845 = ~n1757 & ~n1844 ;
  assign n1846 = ~n1765 & n1845 ;
  assign n1847 = \u3_u1_slv_dout_reg[5]/P0001  & n1756 ;
  assign n1848 = n1755 & n1847 ;
  assign n1849 = \u0_u0_ch_tot_sz_r_reg[5]/P0001  & ~n1757 ;
  assign n1850 = n1765 & n1849 ;
  assign n1851 = ~n1848 & ~n1850 ;
  assign n1852 = ~n1846 & n1851 ;
  assign n1853 = \u2_tsz_cnt_reg[6]/NET0131  & n1004 ;
  assign n1854 = \u3_u0_mast_dout_reg[6]/P0001  & ~n1004 ;
  assign n1855 = ~n1853 & ~n1854 ;
  assign n1856 = ~n1757 & ~n1855 ;
  assign n1857 = ~n1765 & n1856 ;
  assign n1858 = \u3_u1_slv_dout_reg[6]/P0001  & n1756 ;
  assign n1859 = n1755 & n1858 ;
  assign n1860 = \u0_u0_ch_tot_sz_r_reg[6]/P0001  & ~n1757 ;
  assign n1861 = n1765 & n1860 ;
  assign n1862 = ~n1859 & ~n1861 ;
  assign n1863 = ~n1857 & n1862 ;
  assign n1864 = \u2_tsz_cnt_reg[7]/NET0131  & n1004 ;
  assign n1865 = \u3_u0_mast_dout_reg[7]/P0001  & ~n1004 ;
  assign n1866 = ~n1864 & ~n1865 ;
  assign n1867 = ~n1757 & ~n1866 ;
  assign n1868 = ~n1765 & n1867 ;
  assign n1869 = \u3_u1_slv_dout_reg[7]/P0001  & n1756 ;
  assign n1870 = n1755 & n1869 ;
  assign n1871 = \u0_u0_ch_tot_sz_r_reg[7]/P0001  & ~n1757 ;
  assign n1872 = n1765 & n1871 ;
  assign n1873 = ~n1870 & ~n1872 ;
  assign n1874 = ~n1868 & n1873 ;
  assign n1875 = \u2_tsz_cnt_reg[8]/NET0131  & n1004 ;
  assign n1876 = \u3_u0_mast_dout_reg[8]/P0001  & ~n1004 ;
  assign n1877 = ~n1875 & ~n1876 ;
  assign n1878 = ~n1757 & ~n1877 ;
  assign n1879 = ~n1765 & n1878 ;
  assign n1880 = \u3_u1_slv_dout_reg[8]/P0001  & n1756 ;
  assign n1881 = n1755 & n1880 ;
  assign n1882 = \u0_u0_ch_tot_sz_r_reg[8]/P0001  & ~n1757 ;
  assign n1883 = n1765 & n1882 ;
  assign n1884 = ~n1881 & ~n1883 ;
  assign n1885 = ~n1879 & n1884 ;
  assign n1886 = \u2_tsz_cnt_reg[9]/NET0131  & n1004 ;
  assign n1887 = \u3_u0_mast_dout_reg[9]/P0001  & ~n1004 ;
  assign n1888 = ~n1886 & ~n1887 ;
  assign n1889 = ~n1757 & ~n1888 ;
  assign n1890 = ~n1765 & n1889 ;
  assign n1891 = \u3_u1_slv_dout_reg[9]/P0001  & n1756 ;
  assign n1892 = n1755 & n1891 ;
  assign n1893 = \u0_u0_ch_tot_sz_r_reg[9]/P0001  & ~n1757 ;
  assign n1894 = n1765 & n1893 ;
  assign n1895 = ~n1892 & ~n1894 ;
  assign n1896 = ~n1890 & n1895 ;
  assign n1897 = \u0_u0_ch_chk_sz_r_reg[0]/P0001  & ~n1389 ;
  assign n1898 = ~\u2_chunk_cnt_reg[0]/NET0131  & n1738 ;
  assign n1899 = \u2_chunk_cnt_reg[0]/NET0131  & ~n1738 ;
  assign n1900 = ~n1898 & ~n1899 ;
  assign n1901 = n1389 & ~n1900 ;
  assign n1902 = ~n1897 & ~n1901 ;
  assign n1903 = \u0_u0_ch_chk_sz_r_reg[1]/P0001  & ~n1389 ;
  assign n1904 = \u2_chunk_cnt_reg[1]/NET0131  & ~n1898 ;
  assign n1905 = ~n1739 & ~n1904 ;
  assign n1906 = n1389 & ~n1905 ;
  assign n1907 = ~n1903 & ~n1906 ;
  assign n1908 = \u0_u0_ch_chk_sz_r_reg[2]/P0001  & ~n1389 ;
  assign n1909 = ~\u2_chunk_cnt_reg[2]/NET0131  & n1739 ;
  assign n1910 = \u2_chunk_cnt_reg[2]/NET0131  & ~n1739 ;
  assign n1911 = ~n1909 & ~n1910 ;
  assign n1912 = n1389 & ~n1911 ;
  assign n1913 = ~n1908 & ~n1912 ;
  assign n1914 = \u0_u0_ch_chk_sz_r_reg[3]/P0001  & ~n1389 ;
  assign n1915 = n915 & n1739 ;
  assign n1916 = \u2_chunk_cnt_reg[3]/NET0131  & ~n1909 ;
  assign n1917 = ~n1915 & ~n1916 ;
  assign n1918 = n1389 & ~n1917 ;
  assign n1919 = ~n1914 & ~n1918 ;
  assign n1920 = \u0_u0_ch_chk_sz_r_reg[4]/P0001  & ~n1389 ;
  assign n1921 = \u2_chunk_cnt_reg[4]/NET0131  & ~n1915 ;
  assign n1922 = ~n1742 & ~n1921 ;
  assign n1923 = n1389 & ~n1922 ;
  assign n1924 = ~n1920 & ~n1923 ;
  assign n1925 = \u0_u0_ch_chk_sz_r_reg[5]/P0001  & ~n1389 ;
  assign n1926 = ~\u2_chunk_cnt_reg[5]/NET0131  & n1742 ;
  assign n1927 = \u2_chunk_cnt_reg[5]/NET0131  & ~n1742 ;
  assign n1928 = ~n1926 & ~n1927 ;
  assign n1929 = n1389 & ~n1928 ;
  assign n1930 = ~n1925 & ~n1929 ;
  assign n1931 = \u0_u0_ch_chk_sz_r_reg[6]/P0001  & ~n1389 ;
  assign n1932 = ~\u1_next_start_reg/P0001  & \u2_chunk_cnt_reg[6]/NET0131  ;
  assign n1933 = ~n755 & n1932 ;
  assign n1934 = ~n1926 & n1933 ;
  assign n1935 = ~\u1_next_start_reg/P0001  & ~\u2_chunk_cnt_reg[6]/NET0131  ;
  assign n1936 = ~n755 & n1935 ;
  assign n1937 = n1926 & n1936 ;
  assign n1938 = ~n1934 & ~n1937 ;
  assign n1939 = ~n1931 & n1938 ;
  assign n1940 = ~\u0_u0_ch_chk_sz_r_reg[7]/P0001  & ~n1389 ;
  assign n1941 = ~\u2_chunk_cnt_reg[5]/NET0131  & ~\u2_chunk_cnt_reg[6]/NET0131  ;
  assign n1942 = n1742 & n1941 ;
  assign n1943 = \u2_chunk_cnt_reg[7]/NET0131  & ~n1942 ;
  assign n1944 = n1389 & ~n1744 ;
  assign n1945 = ~n1943 & n1944 ;
  assign n1946 = ~n1940 & ~n1945 ;
  assign n1947 = ~\u0_u0_ch_chk_sz_r_reg[6]/P0001  & ~\u0_u0_ch_chk_sz_r_reg[7]/P0001  ;
  assign n1948 = ~\u0_u0_ch_chk_sz_r_reg[8]/P0001  & n1947 ;
  assign n1949 = ~\u0_u0_ch_chk_sz_r_reg[0]/P0001  & ~\u0_u0_ch_chk_sz_r_reg[1]/P0001  ;
  assign n1950 = ~\u0_u0_ch_chk_sz_r_reg[2]/P0001  & ~\u0_u0_ch_chk_sz_r_reg[3]/P0001  ;
  assign n1951 = ~\u0_u0_ch_chk_sz_r_reg[4]/P0001  & ~\u0_u0_ch_chk_sz_r_reg[5]/P0001  ;
  assign n1952 = n1950 & n1951 ;
  assign n1953 = n1949 & n1952 ;
  assign n1954 = n1948 & n1953 ;
  assign n1955 = \u2_adr0_cnt_reg[0]/P0001  & \u2_adr0_cnt_reg[1]/P0001  ;
  assign n1956 = \u2_adr0_cnt_reg[2]/P0001  & \u2_adr0_cnt_reg[3]/P0001  ;
  assign n1957 = n1955 & n1956 ;
  assign n1958 = \u2_adr0_cnt_reg[4]/P0001  & \u2_adr0_cnt_reg[6]/P0001  ;
  assign n1959 = \u2_adr0_cnt_reg[5]/P0001  & n1958 ;
  assign n1960 = n1957 & n1959 ;
  assign n1961 = \u2_adr0_cnt_reg[7]/P0001  & \u2_adr0_cnt_reg[9]/P0001  ;
  assign n1962 = \u2_adr0_cnt_reg[8]/P0001  & n1961 ;
  assign n1963 = n1960 & n1962 ;
  assign n1964 = \u2_adr0_cnt_reg[10]/P0001  & \u2_adr0_cnt_reg[11]/P0001  ;
  assign n1965 = n1963 & n1964 ;
  assign n1966 = ~\u2_adr0_cnt_reg[12]/P0001  & ~n1965 ;
  assign n1967 = \u2_adr0_cnt_reg[11]/P0001  & \u2_adr0_cnt_reg[12]/P0001  ;
  assign n1968 = \u2_adr0_cnt_reg[10]/P0001  & n1967 ;
  assign n1969 = n1963 & n1968 ;
  assign n1970 = ~n1966 & ~n1969 ;
  assign n1971 = \u2_adr1_cnt_reg[0]/P0001  & \u2_adr1_cnt_reg[1]/P0001  ;
  assign n1972 = \u2_adr1_cnt_reg[2]/P0001  & \u2_adr1_cnt_reg[3]/P0001  ;
  assign n1973 = n1971 & n1972 ;
  assign n1974 = \u2_adr1_cnt_reg[4]/P0001  & \u2_adr1_cnt_reg[6]/P0001  ;
  assign n1975 = \u2_adr1_cnt_reg[5]/P0001  & n1974 ;
  assign n1976 = n1973 & n1975 ;
  assign n1977 = \u2_adr1_cnt_reg[7]/P0001  & \u2_adr1_cnt_reg[9]/P0001  ;
  assign n1978 = \u2_adr1_cnt_reg[8]/P0001  & n1977 ;
  assign n1979 = n1976 & n1978 ;
  assign n1980 = \u2_adr1_cnt_reg[10]/P0001  & \u2_adr1_cnt_reg[11]/P0001  ;
  assign n1981 = n1979 & n1980 ;
  assign n1982 = ~\u2_adr1_cnt_reg[12]/P0001  & ~n1981 ;
  assign n1983 = \u2_adr1_cnt_reg[11]/P0001  & \u2_adr1_cnt_reg[12]/P0001  ;
  assign n1984 = \u2_adr1_cnt_reg[10]/P0001  & n1983 ;
  assign n1985 = n1979 & n1984 ;
  assign n1986 = ~n1982 & ~n1985 ;
  assign n1987 = ~\u3_u1_slv_adr_reg[5]/P0001  & n1355 ;
  assign n1988 = \u3_u1_slv_adr_reg[2]/NET0131  & \u3_u1_slv_adr_reg[3]/P0001  ;
  assign n1989 = ~\u3_u1_slv_adr_reg[4]/NET0131  & ~n1988 ;
  assign n1990 = n1987 & ~n1989 ;
  assign n1991 = \u3_u1_slv_adr_reg[3]/P0001  & \u3_u1_slv_adr_reg[4]/NET0131  ;
  assign n1992 = n1355 & n1991 ;
  assign n1993 = ~n1424 & ~n1992 ;
  assign n1994 = ~n1990 & n1993 ;
  assign n1995 = ~\u3_u1_slv_adr_reg[2]/NET0131  & ~\u3_u1_slv_adr_reg[5]/P0001  ;
  assign n1996 = ~\u3_u1_slv_adr_reg[3]/P0001  & n1995 ;
  assign n1997 = \u3_u1_slv_adr_reg[3]/P0001  & ~n1995 ;
  assign n1998 = n1355 & ~n1997 ;
  assign n1999 = ~n1996 & n1998 ;
  assign n2000 = ~\u3_u1_slv_adr_reg[2]/NET0131  & \u3_u1_slv_adr_reg[5]/P0001  ;
  assign n2001 = ~n1422 & n2000 ;
  assign n2002 = n1355 & n2001 ;
  assign n2003 = \u0_u0_ch_adr1_r_reg[7]/P0001  & n2002 ;
  assign n2004 = n1999 & n2003 ;
  assign n2005 = n1994 & n2004 ;
  assign n2006 = \u3_u1_slv_adr_reg[2]/NET0131  & \u3_u1_slv_adr_reg[5]/P0001  ;
  assign n2007 = ~n1422 & n2006 ;
  assign n2008 = n1355 & n2007 ;
  assign n2009 = n1994 & n2008 ;
  assign n2010 = ~n2005 & ~n2009 ;
  assign n2011 = \u3_u1_slv_adr_reg[5]/P0001  & ~n1422 ;
  assign n2012 = n1355 & n2011 ;
  assign n2013 = ~n1995 & ~n2006 ;
  assign n2014 = n1355 & ~n2013 ;
  assign n2015 = ~n2012 & n2014 ;
  assign n2016 = n1999 & n2015 ;
  assign n2017 = ~n1994 & n2016 ;
  assign n2018 = \u0_u0_ch_tot_sz_r_reg[9]/P0001  & n2017 ;
  assign n2019 = ~n2012 & ~n2014 ;
  assign n2020 = n1999 & n2019 ;
  assign n2021 = n1994 & n2020 ;
  assign n2022 = \u0_int_maska_r_reg[9]/NET0131  & n2021 ;
  assign n2023 = ~n2018 & ~n2022 ;
  assign n2024 = n1994 & n2016 ;
  assign n2025 = \u0_int_maskb_r_reg[9]/NET0131  & n2024 ;
  assign n2026 = \u0_u0_ch_adr0_r_reg[7]/P0001  & n2002 ;
  assign n2027 = ~n1999 & n2026 ;
  assign n2028 = n1994 & n2027 ;
  assign n2029 = ~n2025 & ~n2028 ;
  assign n2030 = n2023 & n2029 ;
  assign n2031 = n2010 & n2030 ;
  assign n2032 = ~n1994 & n2020 ;
  assign n2033 = \u0_u0_ch_err_reg/NET0131  & n2032 ;
  assign n2034 = ~n2009 & ~n2033 ;
  assign n2035 = \u0_u0_ch_adr1_r_reg[10]/P0001  & n2002 ;
  assign n2036 = n1999 & n2035 ;
  assign n2037 = n1994 & n2036 ;
  assign n2038 = \u0_u0_ch_adr0_r_reg[10]/P0001  & n2002 ;
  assign n2039 = ~n1999 & n2038 ;
  assign n2040 = n1994 & n2039 ;
  assign n2041 = ~n2037 & ~n2040 ;
  assign n2042 = \u0_int_maska_r_reg[12]/NET0131  & n2021 ;
  assign n2043 = \u0_int_maskb_r_reg[12]/NET0131  & n2024 ;
  assign n2044 = ~n2042 & ~n2043 ;
  assign n2045 = n2041 & n2044 ;
  assign n2046 = n2034 & n2045 ;
  assign n2047 = \u0_u0_ch_adr0_r_reg[11]/P0001  & n2002 ;
  assign n2048 = ~n1999 & n2047 ;
  assign n2049 = n1994 & n2048 ;
  assign n2050 = ~n2009 & ~n2049 ;
  assign n2051 = \u0_u0_ch_csr_r2_reg[0]/NET0131  & n2032 ;
  assign n2052 = \u0_int_maska_r_reg[13]/NET0131  & n2021 ;
  assign n2053 = ~n2051 & ~n2052 ;
  assign n2054 = \u0_int_maskb_r_reg[13]/NET0131  & n2024 ;
  assign n2055 = \u0_u0_ch_adr1_r_reg[11]/P0001  & n2002 ;
  assign n2056 = n1999 & n2055 ;
  assign n2057 = n1994 & n2056 ;
  assign n2058 = ~n2054 & ~n2057 ;
  assign n2059 = n2053 & n2058 ;
  assign n2060 = n2050 & n2059 ;
  assign n2061 = \u0_u0_ch_adr0_r_reg[12]/P0001  & n2002 ;
  assign n2062 = ~n1999 & n2061 ;
  assign n2063 = n1994 & n2062 ;
  assign n2064 = ~n2009 & ~n2063 ;
  assign n2065 = \u0_u0_ch_csr_r2_reg[1]/NET0131  & n2032 ;
  assign n2066 = \u0_int_maska_r_reg[14]/NET0131  & n2021 ;
  assign n2067 = ~n2065 & ~n2066 ;
  assign n2068 = \u0_int_maskb_r_reg[14]/NET0131  & n2024 ;
  assign n2069 = \u0_u0_ch_adr1_r_reg[12]/P0001  & n2002 ;
  assign n2070 = n1999 & n2069 ;
  assign n2071 = n1994 & n2070 ;
  assign n2072 = ~n2068 & ~n2071 ;
  assign n2073 = n2067 & n2072 ;
  assign n2074 = n2064 & n2073 ;
  assign n2075 = \u0_u0_ch_adr0_r_reg[21]/P0001  & n2002 ;
  assign n2076 = ~n1999 & n2075 ;
  assign n2077 = n1994 & n2076 ;
  assign n2078 = ~n2009 & ~n2077 ;
  assign n2079 = \u0_int_maskb_r_reg[23]/NET0131  & n2024 ;
  assign n2080 = \u0_u0_ch_adr1_r_reg[21]/P0001  & n2002 ;
  assign n2081 = n1999 & n2080 ;
  assign n2082 = n1994 & n2081 ;
  assign n2083 = ~n2079 & ~n2082 ;
  assign n2084 = \u0_int_maska_r_reg[23]/NET0131  & n2021 ;
  assign n2085 = \u0_u0_ch_chk_sz_r_reg[7]/P0001  & n2017 ;
  assign n2086 = ~n2084 & ~n2085 ;
  assign n2087 = n2083 & n2086 ;
  assign n2088 = n2078 & n2087 ;
  assign n2089 = \u0_u0_ch_adr0_r_reg[22]/P0001  & n2002 ;
  assign n2090 = ~n1999 & n2089 ;
  assign n2091 = n1994 & n2090 ;
  assign n2092 = ~n2009 & ~n2091 ;
  assign n2093 = \u0_int_maskb_r_reg[24]/NET0131  & n2024 ;
  assign n2094 = \u0_u0_ch_adr1_r_reg[22]/P0001  & n2002 ;
  assign n2095 = n1999 & n2094 ;
  assign n2096 = n1994 & n2095 ;
  assign n2097 = ~n2093 & ~n2096 ;
  assign n2098 = \u0_int_maska_r_reg[24]/NET0131  & n2021 ;
  assign n2099 = \u0_u0_ch_chk_sz_r_reg[8]/P0001  & n2017 ;
  assign n2100 = ~n2098 & ~n2099 ;
  assign n2101 = n2097 & n2100 ;
  assign n2102 = n2092 & n2101 ;
  assign n2103 = \u0_u0_ch_adr0_r_reg[23]/P0001  & n2002 ;
  assign n2104 = ~n1999 & n2103 ;
  assign n2105 = n1994 & n2104 ;
  assign n2106 = ~n2009 & ~n2105 ;
  assign n2107 = \u0_u0_ch_chk_sz_r_reg[9]/P0001  & n2017 ;
  assign n2108 = \u0_int_maska_r_reg[25]/NET0131  & n2021 ;
  assign n2109 = ~n2107 & ~n2108 ;
  assign n2110 = \u0_int_maskb_r_reg[25]/NET0131  & n2024 ;
  assign n2111 = \u0_u0_ch_adr1_r_reg[23]/P0001  & n2002 ;
  assign n2112 = n1999 & n2111 ;
  assign n2113 = n1994 & n2112 ;
  assign n2114 = ~n2110 & ~n2113 ;
  assign n2115 = n2109 & n2114 ;
  assign n2116 = n2106 & n2115 ;
  assign n2117 = \u0_u0_ch_adr0_r_reg[24]/P0001  & n2002 ;
  assign n2118 = ~n1999 & n2117 ;
  assign n2119 = n1994 & n2118 ;
  assign n2120 = ~n2009 & ~n2119 ;
  assign n2121 = \u0_u0_ch_chk_sz_r_reg[10]/P0001  & n2017 ;
  assign n2122 = \u0_int_maska_r_reg[26]/NET0131  & n2021 ;
  assign n2123 = ~n2121 & ~n2122 ;
  assign n2124 = \u0_int_maskb_r_reg[26]/NET0131  & n2024 ;
  assign n2125 = \u0_u0_ch_adr1_r_reg[24]/P0001  & n2002 ;
  assign n2126 = n1999 & n2125 ;
  assign n2127 = n1994 & n2126 ;
  assign n2128 = ~n2124 & ~n2127 ;
  assign n2129 = n2123 & n2128 ;
  assign n2130 = n2120 & n2129 ;
  assign n2131 = \u0_u0_ch_adr0_r_reg[0]/P0001  & n2002 ;
  assign n2132 = ~n1999 & n2131 ;
  assign n2133 = n1994 & n2132 ;
  assign n2134 = \u0_u0_ch_adr1_r_reg[0]/P0001  & n2002 ;
  assign n2135 = n1999 & n2134 ;
  assign n2136 = n1994 & n2135 ;
  assign n2137 = ~n2133 & ~n2136 ;
  assign n2138 = \u0_u0_ch_csr_r_reg[2]/NET0131  & n2032 ;
  assign n2139 = \u0_int_maska_r_reg[2]/NET0131  & n2021 ;
  assign n2140 = ~n2138 & ~n2139 ;
  assign n2141 = \u0_u0_ch_tot_sz_r_reg[2]/P0001  & n2017 ;
  assign n2142 = \u0_int_maskb_r_reg[2]/NET0131  & n2024 ;
  assign n2143 = ~n2141 & ~n2142 ;
  assign n2144 = n2140 & n2143 ;
  assign n2145 = n2137 & n2144 ;
  assign n2146 = \u0_u0_ch_adr0_r_reg[1]/P0001  & n2002 ;
  assign n2147 = ~n1999 & n2146 ;
  assign n2148 = n1994 & n2147 ;
  assign n2149 = \u0_u0_ch_adr1_r_reg[1]/P0001  & n2002 ;
  assign n2150 = n1999 & n2149 ;
  assign n2151 = n1994 & n2150 ;
  assign n2152 = ~n2148 & ~n2151 ;
  assign n2153 = \u0_u0_ch_csr_r_reg[3]/NET0131  & n2032 ;
  assign n2154 = \u0_int_maska_r_reg[3]/NET0131  & n2021 ;
  assign n2155 = ~n2153 & ~n2154 ;
  assign n2156 = \u0_u0_ch_tot_sz_r_reg[3]/P0001  & n2017 ;
  assign n2157 = \u0_int_maskb_r_reg[3]/NET0131  & n2024 ;
  assign n2158 = ~n2156 & ~n2157 ;
  assign n2159 = n2155 & n2158 ;
  assign n2160 = n2152 & n2159 ;
  assign n2161 = \u2_adr0_cnt_reg[13]/P0001  & \u2_adr0_cnt_reg[14]/P0001  ;
  assign n2162 = n1968 & n2161 ;
  assign n2163 = n1963 & n2162 ;
  assign n2164 = \u2_adr0_cnt_reg[15]/P0001  & n2163 ;
  assign n2165 = \u2_adr1_cnt_reg[13]/P0001  & \u2_adr1_cnt_reg[14]/P0001  ;
  assign n2166 = n1984 & n2165 ;
  assign n2167 = n1979 & n2166 ;
  assign n2168 = \u2_adr1_cnt_reg[15]/P0001  & n2167 ;
  assign n2169 = \u0_int_maskb_r_reg[0]/NET0131  & n2024 ;
  assign n2170 = n1994 & ~n1999 ;
  assign n2171 = \u2_state_reg[10]/NET0131  & n2015 ;
  assign n2172 = n2170 & n2171 ;
  assign n2173 = \u0_u0_ch_csr_r3_reg[2]/NET0131  & \u0_u0_int_src_r_reg[2]/NET0131  ;
  assign n2174 = \u0_u0_ch_csr_r3_reg[1]/NET0131  & \u0_u0_int_src_r_reg[1]/NET0131  ;
  assign n2175 = \u0_u0_ch_csr_r3_reg[0]/NET0131  & \u0_u0_ch_err_reg/NET0131  ;
  assign n2176 = ~n2174 & ~n2175 ;
  assign n2177 = ~n2173 & n2176 ;
  assign n2178 = \u0_int_maska_r_reg[0]/NET0131  & ~n2177 ;
  assign n2179 = n2019 & n2178 ;
  assign n2180 = \u0_int_maskb_r_reg[0]/NET0131  & ~n2177 ;
  assign n2181 = n2015 & n2180 ;
  assign n2182 = ~n2179 & ~n2181 ;
  assign n2183 = ~n1994 & ~n1999 ;
  assign n2184 = ~n2182 & n2183 ;
  assign n2185 = ~n2172 & ~n2184 ;
  assign n2186 = ~n2169 & n2185 ;
  assign n2187 = \u0_int_maska_r_reg[0]/NET0131  & n2021 ;
  assign n2188 = \u0_u0_ch_tot_sz_r_reg[0]/P0001  & n2017 ;
  assign n2189 = \u0_u0_ch_csr_r_reg[0]/NET0131  & n2032 ;
  assign n2190 = ~n2188 & ~n2189 ;
  assign n2191 = ~n2187 & n2190 ;
  assign n2192 = n2186 & n2191 ;
  assign n2193 = \u2_adr0_cnt_reg[7]/P0001  & \u2_adr0_cnt_reg[8]/P0001  ;
  assign n2194 = n1960 & n2193 ;
  assign n2195 = \u2_adr0_cnt_reg[7]/P0001  & n1960 ;
  assign n2196 = ~\u2_adr0_cnt_reg[8]/P0001  & ~n2195 ;
  assign n2197 = ~n2194 & ~n2196 ;
  assign n2198 = \u2_adr1_cnt_reg[7]/P0001  & \u2_adr1_cnt_reg[8]/P0001  ;
  assign n2199 = n1976 & n2198 ;
  assign n2200 = \u2_adr1_cnt_reg[7]/P0001  & n1976 ;
  assign n2201 = ~\u2_adr1_cnt_reg[8]/P0001  & ~n2200 ;
  assign n2202 = ~n2199 & ~n2201 ;
  assign n2203 = ~\u3_u1_slv_adr_reg[2]/NET0131  & \u3_u1_slv_adr_reg[3]/P0001  ;
  assign n2204 = n1755 & n2203 ;
  assign n2205 = \u2_mast0_drdy_r_reg/P0001  & \u2_state_reg[6]/NET0131  ;
  assign n2206 = ~\u0_u0_ch_adr0_r_reg[10]/P0001  & ~n2205 ;
  assign n2207 = ~n1409 & n2206 ;
  assign n2208 = ~n2204 & n2207 ;
  assign n2209 = ~n1409 & ~n2205 ;
  assign n2210 = \u3_u0_mast_dout_reg[12]/P0001  & ~n1004 ;
  assign n2211 = \u2_adr0_cnt_reg[10]/P0001  & n1004 ;
  assign n2212 = ~n2210 & ~n2211 ;
  assign n2213 = ~n2204 & n2212 ;
  assign n2214 = ~n2209 & n2213 ;
  assign n2215 = ~n2208 & ~n2214 ;
  assign n2216 = ~\u3_u1_slv_dout_reg[12]/P0001  & n2203 ;
  assign n2217 = n1755 & n2216 ;
  assign n2218 = n2215 & ~n2217 ;
  assign n2219 = ~\u0_u0_ch_adr0_r_reg[11]/P0001  & ~n2205 ;
  assign n2220 = ~n1409 & n2219 ;
  assign n2221 = ~n2204 & n2220 ;
  assign n2222 = \u2_adr0_cnt_reg[11]/P0001  & n1004 ;
  assign n2223 = \u3_u0_mast_dout_reg[13]/P0001  & ~n1004 ;
  assign n2224 = ~n2222 & ~n2223 ;
  assign n2225 = ~n2204 & n2224 ;
  assign n2226 = ~n2209 & n2225 ;
  assign n2227 = ~n2221 & ~n2226 ;
  assign n2228 = ~\u3_u1_slv_dout_reg[13]/P0001  & n2203 ;
  assign n2229 = n1755 & n2228 ;
  assign n2230 = n2227 & ~n2229 ;
  assign n2231 = ~\u0_u0_ch_adr0_r_reg[12]/P0001  & ~n2205 ;
  assign n2232 = ~n1409 & n2231 ;
  assign n2233 = ~n2204 & n2232 ;
  assign n2234 = \u2_adr0_cnt_reg[12]/P0001  & n1004 ;
  assign n2235 = \u3_u0_mast_dout_reg[14]/P0001  & ~n1004 ;
  assign n2236 = ~n2234 & ~n2235 ;
  assign n2237 = ~n2204 & n2236 ;
  assign n2238 = ~n2209 & n2237 ;
  assign n2239 = ~n2233 & ~n2238 ;
  assign n2240 = ~\u3_u1_slv_dout_reg[14]/P0001  & n2203 ;
  assign n2241 = n1755 & n2240 ;
  assign n2242 = n2239 & ~n2241 ;
  assign n2243 = ~\u0_u0_ch_adr0_r_reg[13]/P0001  & ~n2205 ;
  assign n2244 = ~n1409 & n2243 ;
  assign n2245 = ~n2204 & n2244 ;
  assign n2246 = \u2_adr0_cnt_reg[13]/P0001  & n1004 ;
  assign n2247 = \u3_u0_mast_dout_reg[15]/P0001  & ~n1004 ;
  assign n2248 = ~n2246 & ~n2247 ;
  assign n2249 = ~n2204 & n2248 ;
  assign n2250 = ~n2209 & n2249 ;
  assign n2251 = ~n2245 & ~n2250 ;
  assign n2252 = ~\u3_u1_slv_dout_reg[15]/P0001  & n2203 ;
  assign n2253 = n1755 & n2252 ;
  assign n2254 = n2251 & ~n2253 ;
  assign n2255 = ~\u0_u0_ch_adr0_r_reg[14]/P0001  & ~n2205 ;
  assign n2256 = ~n1409 & n2255 ;
  assign n2257 = ~n2204 & n2256 ;
  assign n2258 = \u2_adr0_cnt_reg[14]/P0001  & n1004 ;
  assign n2259 = \u3_u0_mast_dout_reg[16]/P0001  & ~n1004 ;
  assign n2260 = ~n2258 & ~n2259 ;
  assign n2261 = ~n2204 & n2260 ;
  assign n2262 = ~n2209 & n2261 ;
  assign n2263 = ~n2257 & ~n2262 ;
  assign n2264 = ~\u3_u1_slv_dout_reg[16]/P0001  & n2203 ;
  assign n2265 = n1755 & n2264 ;
  assign n2266 = n2263 & ~n2265 ;
  assign n2267 = ~\u0_u0_ch_adr0_r_reg[15]/P0001  & ~n2205 ;
  assign n2268 = ~n1409 & n2267 ;
  assign n2269 = ~n2204 & n2268 ;
  assign n2270 = \u2_adr0_cnt_reg[15]/P0001  & n1004 ;
  assign n2271 = \u3_u0_mast_dout_reg[17]/P0001  & ~n1004 ;
  assign n2272 = ~n2270 & ~n2271 ;
  assign n2273 = ~n2204 & n2272 ;
  assign n2274 = ~n2209 & n2273 ;
  assign n2275 = ~n2269 & ~n2274 ;
  assign n2276 = ~\u3_u1_slv_dout_reg[17]/P0001  & n2203 ;
  assign n2277 = n1755 & n2276 ;
  assign n2278 = n2275 & ~n2277 ;
  assign n2279 = ~\u0_u0_ch_adr0_r_reg[16]/P0001  & ~n2205 ;
  assign n2280 = ~n1409 & n2279 ;
  assign n2281 = ~n2204 & n2280 ;
  assign n2282 = \u2_adr0_cnt_reg[16]/NET0131  & n1004 ;
  assign n2283 = \u3_u0_mast_dout_reg[18]/P0001  & ~n1004 ;
  assign n2284 = ~n2282 & ~n2283 ;
  assign n2285 = ~n2204 & n2284 ;
  assign n2286 = ~n2209 & n2285 ;
  assign n2287 = ~n2281 & ~n2286 ;
  assign n2288 = ~\u3_u1_slv_dout_reg[18]/P0001  & n2203 ;
  assign n2289 = n1755 & n2288 ;
  assign n2290 = n2287 & ~n2289 ;
  assign n2291 = ~\u0_u0_ch_adr0_r_reg[17]/P0001  & ~n2205 ;
  assign n2292 = ~n1409 & n2291 ;
  assign n2293 = ~n2204 & n2292 ;
  assign n2294 = \u2_adr0_cnt_reg[17]/P0001  & n1004 ;
  assign n2295 = \u3_u0_mast_dout_reg[19]/P0001  & ~n1004 ;
  assign n2296 = ~n2294 & ~n2295 ;
  assign n2297 = ~n2204 & n2296 ;
  assign n2298 = ~n2209 & n2297 ;
  assign n2299 = ~n2293 & ~n2298 ;
  assign n2300 = ~\u3_u1_slv_dout_reg[19]/P0001  & n2203 ;
  assign n2301 = n1755 & n2300 ;
  assign n2302 = n2299 & ~n2301 ;
  assign n2303 = ~\u0_u0_ch_adr0_r_reg[18]/P0001  & ~n2205 ;
  assign n2304 = ~n1409 & n2303 ;
  assign n2305 = ~n2204 & n2304 ;
  assign n2306 = \u2_adr0_cnt_reg[18]/P0001  & n1004 ;
  assign n2307 = \u3_u0_mast_dout_reg[20]/P0001  & ~n1004 ;
  assign n2308 = ~n2306 & ~n2307 ;
  assign n2309 = ~n2204 & n2308 ;
  assign n2310 = ~n2209 & n2309 ;
  assign n2311 = ~n2305 & ~n2310 ;
  assign n2312 = ~\u3_u1_slv_dout_reg[20]/P0001  & n2203 ;
  assign n2313 = n1755 & n2312 ;
  assign n2314 = n2311 & ~n2313 ;
  assign n2315 = ~\u0_u0_ch_adr0_r_reg[19]/P0001  & ~n2205 ;
  assign n2316 = ~n1409 & n2315 ;
  assign n2317 = ~n2204 & n2316 ;
  assign n2318 = \u2_adr0_cnt_reg[19]/P0001  & n1004 ;
  assign n2319 = \u3_u0_mast_dout_reg[21]/P0001  & ~n1004 ;
  assign n2320 = ~n2318 & ~n2319 ;
  assign n2321 = ~n2204 & n2320 ;
  assign n2322 = ~n2209 & n2321 ;
  assign n2323 = ~n2317 & ~n2322 ;
  assign n2324 = ~\u3_u1_slv_dout_reg[21]/P0001  & n2203 ;
  assign n2325 = n1755 & n2324 ;
  assign n2326 = n2323 & ~n2325 ;
  assign n2327 = ~\u0_u0_ch_adr0_r_reg[20]/P0001  & ~n2205 ;
  assign n2328 = ~n1409 & n2327 ;
  assign n2329 = ~n2204 & n2328 ;
  assign n2330 = \u2_adr0_cnt_reg[20]/P0001  & n1004 ;
  assign n2331 = \u3_u0_mast_dout_reg[22]/P0001  & ~n1004 ;
  assign n2332 = ~n2330 & ~n2331 ;
  assign n2333 = ~n2204 & n2332 ;
  assign n2334 = ~n2209 & n2333 ;
  assign n2335 = ~n2329 & ~n2334 ;
  assign n2336 = ~\u3_u1_slv_dout_reg[22]/P0001  & n2203 ;
  assign n2337 = n1755 & n2336 ;
  assign n2338 = n2335 & ~n2337 ;
  assign n2339 = ~\u0_u0_ch_adr0_r_reg[21]/P0001  & ~n2205 ;
  assign n2340 = ~n1409 & n2339 ;
  assign n2341 = ~n2204 & n2340 ;
  assign n2342 = \u2_adr0_cnt_reg[21]/P0001  & n1004 ;
  assign n2343 = \u3_u0_mast_dout_reg[23]/P0001  & ~n1004 ;
  assign n2344 = ~n2342 & ~n2343 ;
  assign n2345 = ~n2204 & n2344 ;
  assign n2346 = ~n2209 & n2345 ;
  assign n2347 = ~n2341 & ~n2346 ;
  assign n2348 = ~\u3_u1_slv_dout_reg[23]/P0001  & n2203 ;
  assign n2349 = n1755 & n2348 ;
  assign n2350 = n2347 & ~n2349 ;
  assign n2351 = ~\u0_u0_ch_adr0_r_reg[22]/P0001  & ~n2205 ;
  assign n2352 = ~n1409 & n2351 ;
  assign n2353 = ~n2204 & n2352 ;
  assign n2354 = \u2_adr0_cnt_reg[22]/P0001  & n1004 ;
  assign n2355 = \u3_u0_mast_dout_reg[24]/P0001  & ~n1004 ;
  assign n2356 = ~n2354 & ~n2355 ;
  assign n2357 = ~n2204 & n2356 ;
  assign n2358 = ~n2209 & n2357 ;
  assign n2359 = ~n2353 & ~n2358 ;
  assign n2360 = ~\u3_u1_slv_dout_reg[24]/P0001  & n2203 ;
  assign n2361 = n1755 & n2360 ;
  assign n2362 = n2359 & ~n2361 ;
  assign n2363 = ~\u0_u0_ch_adr0_r_reg[23]/P0001  & ~n2205 ;
  assign n2364 = ~n1409 & n2363 ;
  assign n2365 = ~n2204 & n2364 ;
  assign n2366 = \u2_adr0_cnt_reg[23]/P0001  & n1004 ;
  assign n2367 = \u3_u0_mast_dout_reg[25]/P0001  & ~n1004 ;
  assign n2368 = ~n2366 & ~n2367 ;
  assign n2369 = ~n2204 & n2368 ;
  assign n2370 = ~n2209 & n2369 ;
  assign n2371 = ~n2365 & ~n2370 ;
  assign n2372 = ~\u3_u1_slv_dout_reg[25]/P0001  & n2203 ;
  assign n2373 = n1755 & n2372 ;
  assign n2374 = n2371 & ~n2373 ;
  assign n2375 = ~\u0_u0_ch_adr0_r_reg[24]/P0001  & ~n2205 ;
  assign n2376 = ~n1409 & n2375 ;
  assign n2377 = ~n2204 & n2376 ;
  assign n2378 = \u2_adr0_cnt_reg[24]/P0001  & n1004 ;
  assign n2379 = \u3_u0_mast_dout_reg[26]/P0001  & ~n1004 ;
  assign n2380 = ~n2378 & ~n2379 ;
  assign n2381 = ~n2204 & n2380 ;
  assign n2382 = ~n2209 & n2381 ;
  assign n2383 = ~n2377 & ~n2382 ;
  assign n2384 = ~\u3_u1_slv_dout_reg[26]/P0001  & n2203 ;
  assign n2385 = n1755 & n2384 ;
  assign n2386 = n2383 & ~n2385 ;
  assign n2387 = ~\u0_u0_ch_adr0_r_reg[25]/P0001  & ~n2205 ;
  assign n2388 = ~n1409 & n2387 ;
  assign n2389 = ~n2204 & n2388 ;
  assign n2390 = \u2_adr0_cnt_reg[25]/P0001  & n1004 ;
  assign n2391 = \u3_u0_mast_dout_reg[27]/P0001  & ~n1004 ;
  assign n2392 = ~n2390 & ~n2391 ;
  assign n2393 = ~n2204 & n2392 ;
  assign n2394 = ~n2209 & n2393 ;
  assign n2395 = ~n2389 & ~n2394 ;
  assign n2396 = ~\u3_u1_slv_dout_reg[27]/P0001  & n2203 ;
  assign n2397 = n1755 & n2396 ;
  assign n2398 = n2395 & ~n2397 ;
  assign n2399 = ~\u0_u0_ch_adr0_r_reg[26]/P0001  & ~n2205 ;
  assign n2400 = ~n1409 & n2399 ;
  assign n2401 = ~n2204 & n2400 ;
  assign n2402 = \u2_adr0_cnt_reg[26]/P0001  & n1004 ;
  assign n2403 = \u3_u0_mast_dout_reg[28]/P0001  & ~n1004 ;
  assign n2404 = ~n2402 & ~n2403 ;
  assign n2405 = ~n2204 & n2404 ;
  assign n2406 = ~n2209 & n2405 ;
  assign n2407 = ~n2401 & ~n2406 ;
  assign n2408 = ~\u3_u1_slv_dout_reg[28]/P0001  & n2203 ;
  assign n2409 = n1755 & n2408 ;
  assign n2410 = n2407 & ~n2409 ;
  assign n2411 = ~\u0_u0_ch_adr0_r_reg[27]/P0001  & ~n2205 ;
  assign n2412 = ~n1409 & n2411 ;
  assign n2413 = ~n2204 & n2412 ;
  assign n2414 = \u2_adr0_cnt_reg[27]/P0001  & n1004 ;
  assign n2415 = \u3_u0_mast_dout_reg[29]/P0001  & ~n1004 ;
  assign n2416 = ~n2414 & ~n2415 ;
  assign n2417 = ~n2204 & n2416 ;
  assign n2418 = ~n2209 & n2417 ;
  assign n2419 = ~n2413 & ~n2418 ;
  assign n2420 = ~\u3_u1_slv_dout_reg[29]/P0001  & n2203 ;
  assign n2421 = n1755 & n2420 ;
  assign n2422 = n2419 & ~n2421 ;
  assign n2423 = ~\u0_u0_ch_adr0_r_reg[28]/P0001  & ~n2205 ;
  assign n2424 = ~n1409 & n2423 ;
  assign n2425 = ~n2204 & n2424 ;
  assign n2426 = \u2_adr0_cnt_reg[28]/P0001  & n1004 ;
  assign n2427 = \u3_u0_mast_dout_reg[30]/P0001  & ~n1004 ;
  assign n2428 = ~n2426 & ~n2427 ;
  assign n2429 = ~n2204 & n2428 ;
  assign n2430 = ~n2209 & n2429 ;
  assign n2431 = ~n2425 & ~n2430 ;
  assign n2432 = ~\u3_u1_slv_dout_reg[30]/P0001  & n2203 ;
  assign n2433 = n1755 & n2432 ;
  assign n2434 = n2431 & ~n2433 ;
  assign n2435 = ~\u0_u0_ch_adr0_r_reg[29]/P0001  & ~n2205 ;
  assign n2436 = ~n1409 & n2435 ;
  assign n2437 = ~n2204 & n2436 ;
  assign n2438 = \u2_adr0_cnt_reg[29]/P0001  & n1004 ;
  assign n2439 = \u3_u0_mast_dout_reg[31]/P0001  & ~n1004 ;
  assign n2440 = ~n2438 & ~n2439 ;
  assign n2441 = ~n2204 & n2440 ;
  assign n2442 = ~n2209 & n2441 ;
  assign n2443 = ~n2437 & ~n2442 ;
  assign n2444 = ~\u3_u1_slv_dout_reg[31]/P0001  & n2203 ;
  assign n2445 = n1755 & n2444 ;
  assign n2446 = n2443 & ~n2445 ;
  assign n2447 = \u3_u1_slv_adr_reg[4]/NET0131  & \u3_u1_slv_we_reg/P0001  ;
  assign n2448 = n1358 & n2447 ;
  assign n2449 = ~\u2_mast0_drdy_r_reg/P0001  & \u2_state_reg[7]/NET0131  ;
  assign n2450 = ~\u0_u0_ch_adr1_r_reg[10]/P0001  & n2449 ;
  assign n2451 = ~\u0_u0_ch_adr1_r_reg[10]/P0001  & ~\u2_state_reg[7]/NET0131  ;
  assign n2452 = ~n1409 & n2451 ;
  assign n2453 = ~n2450 & ~n2452 ;
  assign n2454 = ~\u2_state_reg[7]/NET0131  & ~n1409 ;
  assign n2455 = \u2_adr1_cnt_reg[10]/P0001  & n1004 ;
  assign n2456 = ~n2210 & ~n2455 ;
  assign n2457 = ~n2449 & n2456 ;
  assign n2458 = ~n2454 & n2457 ;
  assign n2459 = n2453 & ~n2458 ;
  assign n2460 = ~n2448 & ~n2459 ;
  assign n2461 = ~\u3_u1_slv_dout_reg[12]/P0001  & n2447 ;
  assign n2462 = n1358 & n2461 ;
  assign n2463 = ~n2460 & ~n2462 ;
  assign n2464 = ~\u0_u0_ch_adr1_r_reg[11]/P0001  & n2449 ;
  assign n2465 = ~\u0_u0_ch_adr1_r_reg[11]/P0001  & ~\u2_state_reg[7]/NET0131  ;
  assign n2466 = ~n1409 & n2465 ;
  assign n2467 = ~n2464 & ~n2466 ;
  assign n2468 = \u2_adr1_cnt_reg[11]/P0001  & n1004 ;
  assign n2469 = ~n2223 & ~n2468 ;
  assign n2470 = ~n2449 & n2469 ;
  assign n2471 = ~n2454 & n2470 ;
  assign n2472 = n2467 & ~n2471 ;
  assign n2473 = ~n2448 & ~n2472 ;
  assign n2474 = ~\u3_u1_slv_dout_reg[13]/P0001  & n2447 ;
  assign n2475 = n1358 & n2474 ;
  assign n2476 = ~n2473 & ~n2475 ;
  assign n2477 = ~\u0_u0_ch_adr1_r_reg[12]/P0001  & n2449 ;
  assign n2478 = ~\u0_u0_ch_adr1_r_reg[12]/P0001  & ~\u2_state_reg[7]/NET0131  ;
  assign n2479 = ~n1409 & n2478 ;
  assign n2480 = ~n2477 & ~n2479 ;
  assign n2481 = \u2_adr1_cnt_reg[12]/P0001  & n1004 ;
  assign n2482 = ~n2235 & ~n2481 ;
  assign n2483 = ~n2449 & n2482 ;
  assign n2484 = ~n2454 & n2483 ;
  assign n2485 = n2480 & ~n2484 ;
  assign n2486 = ~n2448 & ~n2485 ;
  assign n2487 = ~\u3_u1_slv_dout_reg[14]/P0001  & n2447 ;
  assign n2488 = n1358 & n2487 ;
  assign n2489 = ~n2486 & ~n2488 ;
  assign n2490 = ~\u0_u0_ch_adr1_r_reg[13]/P0001  & n2449 ;
  assign n2491 = ~\u0_u0_ch_adr1_r_reg[13]/P0001  & ~\u2_state_reg[7]/NET0131  ;
  assign n2492 = ~n1409 & n2491 ;
  assign n2493 = ~n2490 & ~n2492 ;
  assign n2494 = \u2_adr1_cnt_reg[13]/P0001  & n1004 ;
  assign n2495 = ~n2247 & ~n2494 ;
  assign n2496 = ~n2449 & n2495 ;
  assign n2497 = ~n2454 & n2496 ;
  assign n2498 = n2493 & ~n2497 ;
  assign n2499 = ~n2448 & ~n2498 ;
  assign n2500 = ~\u3_u1_slv_dout_reg[15]/P0001  & n2447 ;
  assign n2501 = n1358 & n2500 ;
  assign n2502 = ~n2499 & ~n2501 ;
  assign n2503 = ~\u0_u0_ch_adr1_r_reg[14]/P0001  & n2449 ;
  assign n2504 = ~\u0_u0_ch_adr1_r_reg[14]/P0001  & ~\u2_state_reg[7]/NET0131  ;
  assign n2505 = ~n1409 & n2504 ;
  assign n2506 = ~n2503 & ~n2505 ;
  assign n2507 = \u2_adr1_cnt_reg[14]/P0001  & n1004 ;
  assign n2508 = ~n2259 & ~n2507 ;
  assign n2509 = ~n2449 & n2508 ;
  assign n2510 = ~n2454 & n2509 ;
  assign n2511 = n2506 & ~n2510 ;
  assign n2512 = ~n2448 & ~n2511 ;
  assign n2513 = ~\u3_u1_slv_dout_reg[16]/P0001  & n2447 ;
  assign n2514 = n1358 & n2513 ;
  assign n2515 = ~n2512 & ~n2514 ;
  assign n2516 = ~\u0_u0_ch_adr1_r_reg[15]/P0001  & n2449 ;
  assign n2517 = ~\u0_u0_ch_adr1_r_reg[15]/P0001  & ~\u2_state_reg[7]/NET0131  ;
  assign n2518 = ~n1409 & n2517 ;
  assign n2519 = ~n2516 & ~n2518 ;
  assign n2520 = \u2_adr1_cnt_reg[15]/P0001  & n1004 ;
  assign n2521 = ~n2271 & ~n2520 ;
  assign n2522 = ~n2449 & n2521 ;
  assign n2523 = ~n2454 & n2522 ;
  assign n2524 = n2519 & ~n2523 ;
  assign n2525 = ~n2448 & ~n2524 ;
  assign n2526 = ~\u3_u1_slv_dout_reg[17]/P0001  & n2447 ;
  assign n2527 = n1358 & n2526 ;
  assign n2528 = ~n2525 & ~n2527 ;
  assign n2529 = ~\u0_u0_ch_adr1_r_reg[16]/P0001  & n2449 ;
  assign n2530 = ~\u0_u0_ch_adr1_r_reg[16]/P0001  & ~\u2_state_reg[7]/NET0131  ;
  assign n2531 = ~n1409 & n2530 ;
  assign n2532 = ~n2529 & ~n2531 ;
  assign n2533 = \u2_adr1_cnt_reg[16]/NET0131  & n1004 ;
  assign n2534 = ~n2283 & ~n2533 ;
  assign n2535 = ~n2449 & n2534 ;
  assign n2536 = ~n2454 & n2535 ;
  assign n2537 = n2532 & ~n2536 ;
  assign n2538 = ~n2448 & ~n2537 ;
  assign n2539 = ~\u3_u1_slv_dout_reg[18]/P0001  & n2447 ;
  assign n2540 = n1358 & n2539 ;
  assign n2541 = ~n2538 & ~n2540 ;
  assign n2542 = ~\u0_u0_ch_adr1_r_reg[17]/P0001  & n2449 ;
  assign n2543 = ~\u0_u0_ch_adr1_r_reg[17]/P0001  & ~\u2_state_reg[7]/NET0131  ;
  assign n2544 = ~n1409 & n2543 ;
  assign n2545 = ~n2542 & ~n2544 ;
  assign n2546 = \u2_adr1_cnt_reg[17]/P0001  & n1004 ;
  assign n2547 = ~n2295 & ~n2546 ;
  assign n2548 = ~n2449 & n2547 ;
  assign n2549 = ~n2454 & n2548 ;
  assign n2550 = n2545 & ~n2549 ;
  assign n2551 = ~n2448 & ~n2550 ;
  assign n2552 = ~\u3_u1_slv_dout_reg[19]/P0001  & n2447 ;
  assign n2553 = n1358 & n2552 ;
  assign n2554 = ~n2551 & ~n2553 ;
  assign n2555 = ~\u0_u0_ch_adr1_r_reg[18]/P0001  & n2449 ;
  assign n2556 = ~\u0_u0_ch_adr1_r_reg[18]/P0001  & ~\u2_state_reg[7]/NET0131  ;
  assign n2557 = ~n1409 & n2556 ;
  assign n2558 = ~n2555 & ~n2557 ;
  assign n2559 = \u2_adr1_cnt_reg[18]/P0001  & n1004 ;
  assign n2560 = ~n2307 & ~n2559 ;
  assign n2561 = ~n2449 & n2560 ;
  assign n2562 = ~n2454 & n2561 ;
  assign n2563 = n2558 & ~n2562 ;
  assign n2564 = ~n2448 & ~n2563 ;
  assign n2565 = ~\u3_u1_slv_dout_reg[20]/P0001  & n2447 ;
  assign n2566 = n1358 & n2565 ;
  assign n2567 = ~n2564 & ~n2566 ;
  assign n2568 = ~\u0_u0_ch_adr1_r_reg[19]/P0001  & n2449 ;
  assign n2569 = ~\u0_u0_ch_adr1_r_reg[19]/P0001  & ~\u2_state_reg[7]/NET0131  ;
  assign n2570 = ~n1409 & n2569 ;
  assign n2571 = ~n2568 & ~n2570 ;
  assign n2572 = \u2_adr1_cnt_reg[19]/P0001  & n1004 ;
  assign n2573 = ~n2319 & ~n2572 ;
  assign n2574 = ~n2449 & n2573 ;
  assign n2575 = ~n2454 & n2574 ;
  assign n2576 = n2571 & ~n2575 ;
  assign n2577 = ~n2448 & ~n2576 ;
  assign n2578 = ~\u3_u1_slv_dout_reg[21]/P0001  & n2447 ;
  assign n2579 = n1358 & n2578 ;
  assign n2580 = ~n2577 & ~n2579 ;
  assign n2581 = ~\u0_u0_ch_adr1_r_reg[20]/P0001  & n2449 ;
  assign n2582 = ~\u0_u0_ch_adr1_r_reg[20]/P0001  & ~\u2_state_reg[7]/NET0131  ;
  assign n2583 = ~n1409 & n2582 ;
  assign n2584 = ~n2581 & ~n2583 ;
  assign n2585 = \u2_adr1_cnt_reg[20]/P0001  & n1004 ;
  assign n2586 = ~n2331 & ~n2585 ;
  assign n2587 = ~n2449 & n2586 ;
  assign n2588 = ~n2454 & n2587 ;
  assign n2589 = n2584 & ~n2588 ;
  assign n2590 = ~n2448 & ~n2589 ;
  assign n2591 = ~\u3_u1_slv_dout_reg[22]/P0001  & n2447 ;
  assign n2592 = n1358 & n2591 ;
  assign n2593 = ~n2590 & ~n2592 ;
  assign n2594 = ~\u0_u0_ch_adr1_r_reg[21]/P0001  & n2449 ;
  assign n2595 = ~\u0_u0_ch_adr1_r_reg[21]/P0001  & ~\u2_state_reg[7]/NET0131  ;
  assign n2596 = ~n1409 & n2595 ;
  assign n2597 = ~n2594 & ~n2596 ;
  assign n2598 = \u2_adr1_cnt_reg[21]/P0001  & n1004 ;
  assign n2599 = ~n2343 & ~n2598 ;
  assign n2600 = ~n2449 & n2599 ;
  assign n2601 = ~n2454 & n2600 ;
  assign n2602 = n2597 & ~n2601 ;
  assign n2603 = ~n2448 & ~n2602 ;
  assign n2604 = ~\u3_u1_slv_dout_reg[23]/P0001  & n2447 ;
  assign n2605 = n1358 & n2604 ;
  assign n2606 = ~n2603 & ~n2605 ;
  assign n2607 = ~\u0_u0_ch_adr1_r_reg[22]/P0001  & n2449 ;
  assign n2608 = ~\u0_u0_ch_adr1_r_reg[22]/P0001  & ~\u2_state_reg[7]/NET0131  ;
  assign n2609 = ~n1409 & n2608 ;
  assign n2610 = ~n2607 & ~n2609 ;
  assign n2611 = \u2_adr1_cnt_reg[22]/P0001  & n1004 ;
  assign n2612 = ~n2355 & ~n2611 ;
  assign n2613 = ~n2449 & n2612 ;
  assign n2614 = ~n2454 & n2613 ;
  assign n2615 = n2610 & ~n2614 ;
  assign n2616 = ~n2448 & ~n2615 ;
  assign n2617 = ~\u3_u1_slv_dout_reg[24]/P0001  & n2447 ;
  assign n2618 = n1358 & n2617 ;
  assign n2619 = ~n2616 & ~n2618 ;
  assign n2620 = ~\u0_u0_ch_adr1_r_reg[23]/P0001  & n2449 ;
  assign n2621 = ~\u0_u0_ch_adr1_r_reg[23]/P0001  & ~\u2_state_reg[7]/NET0131  ;
  assign n2622 = ~n1409 & n2621 ;
  assign n2623 = ~n2620 & ~n2622 ;
  assign n2624 = \u2_adr1_cnt_reg[23]/P0001  & n1004 ;
  assign n2625 = ~n2367 & ~n2624 ;
  assign n2626 = ~n2449 & n2625 ;
  assign n2627 = ~n2454 & n2626 ;
  assign n2628 = n2623 & ~n2627 ;
  assign n2629 = ~n2448 & ~n2628 ;
  assign n2630 = ~\u3_u1_slv_dout_reg[25]/P0001  & n2447 ;
  assign n2631 = n1358 & n2630 ;
  assign n2632 = ~n2629 & ~n2631 ;
  assign n2633 = ~\u0_u0_ch_adr1_r_reg[24]/P0001  & n2449 ;
  assign n2634 = ~\u0_u0_ch_adr1_r_reg[24]/P0001  & ~\u2_state_reg[7]/NET0131  ;
  assign n2635 = ~n1409 & n2634 ;
  assign n2636 = ~n2633 & ~n2635 ;
  assign n2637 = \u2_adr1_cnt_reg[24]/P0001  & n1004 ;
  assign n2638 = ~n2379 & ~n2637 ;
  assign n2639 = ~n2449 & n2638 ;
  assign n2640 = ~n2454 & n2639 ;
  assign n2641 = n2636 & ~n2640 ;
  assign n2642 = ~n2448 & ~n2641 ;
  assign n2643 = ~\u3_u1_slv_dout_reg[26]/P0001  & n2447 ;
  assign n2644 = n1358 & n2643 ;
  assign n2645 = ~n2642 & ~n2644 ;
  assign n2646 = ~\u0_u0_ch_adr1_r_reg[25]/P0001  & n2449 ;
  assign n2647 = ~\u0_u0_ch_adr1_r_reg[25]/P0001  & ~\u2_state_reg[7]/NET0131  ;
  assign n2648 = ~n1409 & n2647 ;
  assign n2649 = ~n2646 & ~n2648 ;
  assign n2650 = \u2_adr1_cnt_reg[25]/P0001  & n1004 ;
  assign n2651 = ~n2391 & ~n2650 ;
  assign n2652 = ~n2449 & n2651 ;
  assign n2653 = ~n2454 & n2652 ;
  assign n2654 = n2649 & ~n2653 ;
  assign n2655 = ~n2448 & ~n2654 ;
  assign n2656 = ~\u3_u1_slv_dout_reg[27]/P0001  & n2447 ;
  assign n2657 = n1358 & n2656 ;
  assign n2658 = ~n2655 & ~n2657 ;
  assign n2659 = ~\u0_u0_ch_adr1_r_reg[26]/P0001  & n2449 ;
  assign n2660 = ~\u0_u0_ch_adr1_r_reg[26]/P0001  & ~\u2_state_reg[7]/NET0131  ;
  assign n2661 = ~n1409 & n2660 ;
  assign n2662 = ~n2659 & ~n2661 ;
  assign n2663 = \u2_adr1_cnt_reg[26]/P0001  & n1004 ;
  assign n2664 = ~n2403 & ~n2663 ;
  assign n2665 = ~n2449 & n2664 ;
  assign n2666 = ~n2454 & n2665 ;
  assign n2667 = n2662 & ~n2666 ;
  assign n2668 = ~n2448 & ~n2667 ;
  assign n2669 = ~\u3_u1_slv_dout_reg[28]/P0001  & n2447 ;
  assign n2670 = n1358 & n2669 ;
  assign n2671 = ~n2668 & ~n2670 ;
  assign n2672 = ~\u0_u0_ch_adr1_r_reg[27]/P0001  & n2449 ;
  assign n2673 = ~\u0_u0_ch_adr1_r_reg[27]/P0001  & ~\u2_state_reg[7]/NET0131  ;
  assign n2674 = ~n1409 & n2673 ;
  assign n2675 = ~n2672 & ~n2674 ;
  assign n2676 = \u2_adr1_cnt_reg[27]/P0001  & n1004 ;
  assign n2677 = ~n2415 & ~n2676 ;
  assign n2678 = ~n2449 & n2677 ;
  assign n2679 = ~n2454 & n2678 ;
  assign n2680 = n2675 & ~n2679 ;
  assign n2681 = ~n2448 & ~n2680 ;
  assign n2682 = ~\u3_u1_slv_dout_reg[29]/P0001  & n2447 ;
  assign n2683 = n1358 & n2682 ;
  assign n2684 = ~n2681 & ~n2683 ;
  assign n2685 = ~\u0_u0_ch_adr1_r_reg[28]/P0001  & n2449 ;
  assign n2686 = ~\u0_u0_ch_adr1_r_reg[28]/P0001  & ~\u2_state_reg[7]/NET0131  ;
  assign n2687 = ~n1409 & n2686 ;
  assign n2688 = ~n2685 & ~n2687 ;
  assign n2689 = \u2_adr1_cnt_reg[28]/P0001  & n1004 ;
  assign n2690 = ~n2427 & ~n2689 ;
  assign n2691 = ~n2449 & n2690 ;
  assign n2692 = ~n2454 & n2691 ;
  assign n2693 = n2688 & ~n2692 ;
  assign n2694 = ~n2448 & ~n2693 ;
  assign n2695 = ~\u3_u1_slv_dout_reg[30]/P0001  & n2447 ;
  assign n2696 = n1358 & n2695 ;
  assign n2697 = ~n2694 & ~n2696 ;
  assign n2698 = ~\u0_u0_ch_adr1_r_reg[29]/P0001  & n2449 ;
  assign n2699 = ~\u0_u0_ch_adr1_r_reg[29]/P0001  & ~\u2_state_reg[7]/NET0131  ;
  assign n2700 = ~n1409 & n2699 ;
  assign n2701 = ~n2698 & ~n2700 ;
  assign n2702 = \u2_adr1_cnt_reg[29]/P0001  & n1004 ;
  assign n2703 = ~n2439 & ~n2702 ;
  assign n2704 = ~n2449 & n2703 ;
  assign n2705 = ~n2454 & n2704 ;
  assign n2706 = n2701 & ~n2705 ;
  assign n2707 = ~n2448 & ~n2706 ;
  assign n2708 = ~\u3_u1_slv_dout_reg[31]/P0001  & n2447 ;
  assign n2709 = n1358 & n2708 ;
  assign n2710 = ~n2707 & ~n2709 ;
  assign n2711 = \u2_state_reg[4]/NET0131  & ~\u2_state_reg[6]/NET0131  ;
  assign n2712 = ~\u2_state_reg[7]/NET0131  & n2711 ;
  assign n2713 = n1011 & n2712 ;
  assign n2714 = n1010 & n2713 ;
  assign n2715 = \u0_u0_ch_csr_r_reg[1]/NET0131  & ~n1761 ;
  assign n2716 = ~n2714 & n2715 ;
  assign n2717 = ~n1362 & n2716 ;
  assign n2718 = ~n1761 & ~n2714 ;
  assign n2719 = \u3_u0_mast_dout_reg[16]/P0001  & ~n1362 ;
  assign n2720 = ~n2718 & n2719 ;
  assign n2721 = ~n2717 & ~n2720 ;
  assign n2722 = \u3_u1_slv_dout_reg[1]/P0001  & n1359 ;
  assign n2723 = n1358 & n2722 ;
  assign n2724 = n2721 & ~n2723 ;
  assign n2725 = \u0_u0_ch_csr_r_reg[2]/NET0131  & ~n1761 ;
  assign n2726 = ~n2714 & n2725 ;
  assign n2727 = ~n1362 & n2726 ;
  assign n2728 = \u3_u0_mast_dout_reg[17]/P0001  & ~n1362 ;
  assign n2729 = ~n2718 & n2728 ;
  assign n2730 = ~n2727 & ~n2729 ;
  assign n2731 = \u3_u1_slv_dout_reg[2]/P0001  & n1359 ;
  assign n2732 = n1358 & n2731 ;
  assign n2733 = n2730 & ~n2732 ;
  assign n2734 = \u0_u0_ch_csr_r_reg[3]/NET0131  & ~n1761 ;
  assign n2735 = ~n2714 & n2734 ;
  assign n2736 = ~n1362 & n2735 ;
  assign n2737 = \u3_u0_mast_dout_reg[18]/P0001  & ~n1362 ;
  assign n2738 = ~n2718 & n2737 ;
  assign n2739 = ~n2736 & ~n2738 ;
  assign n2740 = \u3_u1_slv_dout_reg[3]/P0001  & n1359 ;
  assign n2741 = n1358 & n2740 ;
  assign n2742 = n2739 & ~n2741 ;
  assign n2743 = \u0_u0_ch_csr_r_reg[4]/NET0131  & ~n1761 ;
  assign n2744 = ~n2714 & n2743 ;
  assign n2745 = ~n1362 & n2744 ;
  assign n2746 = \u3_u0_mast_dout_reg[19]/P0001  & ~n1362 ;
  assign n2747 = ~n2718 & n2746 ;
  assign n2748 = ~n2745 & ~n2747 ;
  assign n2749 = \u3_u1_slv_dout_reg[4]/P0001  & n1359 ;
  assign n2750 = n1358 & n2749 ;
  assign n2751 = n2748 & ~n2750 ;
  assign n2752 = \u2_adr1_cnt_reg[0]/P0001  & n1004 ;
  assign n2753 = ~n1810 & ~n2752 ;
  assign n2754 = ~n2448 & ~n2449 ;
  assign n2755 = ~n2454 & n2754 ;
  assign n2756 = ~n2753 & n2755 ;
  assign n2757 = \u3_u1_slv_dout_reg[2]/P0001  & n2447 ;
  assign n2758 = n1358 & n2757 ;
  assign n2759 = ~n2449 & ~n2454 ;
  assign n2760 = \u0_u0_ch_adr1_r_reg[0]/P0001  & ~n2448 ;
  assign n2761 = ~n2759 & n2760 ;
  assign n2762 = ~n2758 & ~n2761 ;
  assign n2763 = ~n2756 & n2762 ;
  assign n2764 = \u2_adr1_cnt_reg[2]/P0001  & n1004 ;
  assign n2765 = ~n1832 & ~n2764 ;
  assign n2766 = n2755 & ~n2765 ;
  assign n2767 = \u3_u1_slv_dout_reg[4]/P0001  & n2447 ;
  assign n2768 = n1358 & n2767 ;
  assign n2769 = \u0_u0_ch_adr1_r_reg[2]/P0001  & ~n2448 ;
  assign n2770 = ~n2759 & n2769 ;
  assign n2771 = ~n2768 & ~n2770 ;
  assign n2772 = ~n2766 & n2771 ;
  assign n2773 = \u2_adr1_cnt_reg[1]/P0001  & n1004 ;
  assign n2774 = ~n1821 & ~n2773 ;
  assign n2775 = n2755 & ~n2774 ;
  assign n2776 = \u3_u1_slv_dout_reg[3]/P0001  & n2447 ;
  assign n2777 = n1358 & n2776 ;
  assign n2778 = \u0_u0_ch_adr1_r_reg[1]/P0001  & ~n2448 ;
  assign n2779 = ~n2759 & n2778 ;
  assign n2780 = ~n2777 & ~n2779 ;
  assign n2781 = ~n2775 & n2780 ;
  assign n2782 = \u2_adr1_cnt_reg[3]/P0001  & n1004 ;
  assign n2783 = ~n1843 & ~n2782 ;
  assign n2784 = n2755 & ~n2783 ;
  assign n2785 = \u3_u1_slv_dout_reg[5]/P0001  & n2447 ;
  assign n2786 = n1358 & n2785 ;
  assign n2787 = \u0_u0_ch_adr1_r_reg[3]/P0001  & ~n2448 ;
  assign n2788 = ~n2759 & n2787 ;
  assign n2789 = ~n2786 & ~n2788 ;
  assign n2790 = ~n2784 & n2789 ;
  assign n2791 = \u2_adr1_cnt_reg[4]/P0001  & n1004 ;
  assign n2792 = ~n1854 & ~n2791 ;
  assign n2793 = n2755 & ~n2792 ;
  assign n2794 = \u3_u1_slv_dout_reg[6]/P0001  & n2447 ;
  assign n2795 = n1358 & n2794 ;
  assign n2796 = \u0_u0_ch_adr1_r_reg[4]/P0001  & ~n2448 ;
  assign n2797 = ~n2759 & n2796 ;
  assign n2798 = ~n2795 & ~n2797 ;
  assign n2799 = ~n2793 & n2798 ;
  assign n2800 = \u2_adr1_cnt_reg[5]/P0001  & n1004 ;
  assign n2801 = ~n1865 & ~n2800 ;
  assign n2802 = n2755 & ~n2801 ;
  assign n2803 = \u3_u1_slv_dout_reg[7]/P0001  & n2447 ;
  assign n2804 = n1358 & n2803 ;
  assign n2805 = \u0_u0_ch_adr1_r_reg[5]/P0001  & ~n2448 ;
  assign n2806 = ~n2759 & n2805 ;
  assign n2807 = ~n2804 & ~n2806 ;
  assign n2808 = ~n2802 & n2807 ;
  assign n2809 = \u2_adr1_cnt_reg[6]/P0001  & n1004 ;
  assign n2810 = ~n1876 & ~n2809 ;
  assign n2811 = n2755 & ~n2810 ;
  assign n2812 = \u3_u1_slv_dout_reg[8]/P0001  & n2447 ;
  assign n2813 = n1358 & n2812 ;
  assign n2814 = \u0_u0_ch_adr1_r_reg[6]/P0001  & ~n2448 ;
  assign n2815 = ~n2759 & n2814 ;
  assign n2816 = ~n2813 & ~n2815 ;
  assign n2817 = ~n2811 & n2816 ;
  assign n2818 = \u2_adr1_cnt_reg[7]/P0001  & n1004 ;
  assign n2819 = ~n1887 & ~n2818 ;
  assign n2820 = n2755 & ~n2819 ;
  assign n2821 = \u3_u1_slv_dout_reg[9]/P0001  & n2447 ;
  assign n2822 = n1358 & n2821 ;
  assign n2823 = \u0_u0_ch_adr1_r_reg[7]/P0001  & ~n2448 ;
  assign n2824 = ~n2759 & n2823 ;
  assign n2825 = ~n2822 & ~n2824 ;
  assign n2826 = ~n2820 & n2825 ;
  assign n2827 = \u2_adr1_cnt_reg[8]/P0001  & n1004 ;
  assign n2828 = ~n1788 & ~n2827 ;
  assign n2829 = n2755 & ~n2828 ;
  assign n2830 = \u3_u1_slv_dout_reg[10]/P0001  & n2447 ;
  assign n2831 = n1358 & n2830 ;
  assign n2832 = \u0_u0_ch_adr1_r_reg[8]/P0001  & ~n2448 ;
  assign n2833 = ~n2759 & n2832 ;
  assign n2834 = ~n2831 & ~n2833 ;
  assign n2835 = ~n2829 & n2834 ;
  assign n2836 = \u2_adr1_cnt_reg[9]/P0001  & n1004 ;
  assign n2837 = ~n1799 & ~n2836 ;
  assign n2838 = n2755 & ~n2837 ;
  assign n2839 = \u3_u1_slv_dout_reg[11]/P0001  & n2447 ;
  assign n2840 = n1358 & n2839 ;
  assign n2841 = \u0_u0_ch_adr1_r_reg[9]/P0001  & ~n2448 ;
  assign n2842 = ~n2759 & n2841 ;
  assign n2843 = ~n2840 & ~n2842 ;
  assign n2844 = ~n2838 & n2843 ;
  assign n2845 = \u0_int_maska_r_reg[27]/NET0131  & n2021 ;
  assign n2846 = \u0_int_maskb_r_reg[27]/NET0131  & n2024 ;
  assign n2847 = ~n2845 & ~n2846 ;
  assign n2848 = \u0_u0_ch_adr1_r_reg[25]/P0001  & n2002 ;
  assign n2849 = n1999 & n2848 ;
  assign n2850 = n1994 & n2849 ;
  assign n2851 = \u0_u0_ch_adr0_r_reg[25]/P0001  & n2002 ;
  assign n2852 = ~n1999 & n2851 ;
  assign n2853 = n1994 & n2852 ;
  assign n2854 = ~n2009 & ~n2853 ;
  assign n2855 = ~n2850 & n2854 ;
  assign n2856 = n2847 & n2855 ;
  assign n2857 = \u0_int_maska_r_reg[28]/NET0131  & n2021 ;
  assign n2858 = \u0_int_maskb_r_reg[28]/NET0131  & n2024 ;
  assign n2859 = ~n2857 & ~n2858 ;
  assign n2860 = \u0_u0_ch_adr1_r_reg[26]/P0001  & n2002 ;
  assign n2861 = n1999 & n2860 ;
  assign n2862 = n1994 & n2861 ;
  assign n2863 = \u0_u0_ch_adr0_r_reg[26]/P0001  & n2002 ;
  assign n2864 = ~n1999 & n2863 ;
  assign n2865 = n1994 & n2864 ;
  assign n2866 = ~n2009 & ~n2865 ;
  assign n2867 = ~n2862 & n2866 ;
  assign n2868 = n2859 & n2867 ;
  assign n2869 = \u0_int_maska_r_reg[29]/NET0131  & n2021 ;
  assign n2870 = \u0_int_maskb_r_reg[29]/NET0131  & n2024 ;
  assign n2871 = ~n2869 & ~n2870 ;
  assign n2872 = \u0_u0_ch_adr1_r_reg[27]/P0001  & n2002 ;
  assign n2873 = n1999 & n2872 ;
  assign n2874 = n1994 & n2873 ;
  assign n2875 = \u0_u0_ch_adr0_r_reg[27]/P0001  & n2002 ;
  assign n2876 = ~n1999 & n2875 ;
  assign n2877 = n1994 & n2876 ;
  assign n2878 = ~n2009 & ~n2877 ;
  assign n2879 = ~n2874 & n2878 ;
  assign n2880 = n2871 & n2879 ;
  assign n2881 = \u0_int_maska_r_reg[30]/NET0131  & n2021 ;
  assign n2882 = \u0_int_maskb_r_reg[30]/NET0131  & n2024 ;
  assign n2883 = ~n2881 & ~n2882 ;
  assign n2884 = \u0_u0_ch_adr1_r_reg[28]/P0001  & n2002 ;
  assign n2885 = n1999 & n2884 ;
  assign n2886 = n1994 & n2885 ;
  assign n2887 = \u0_u0_ch_adr0_r_reg[28]/P0001  & n2002 ;
  assign n2888 = ~n1999 & n2887 ;
  assign n2889 = n1994 & n2888 ;
  assign n2890 = ~n2009 & ~n2889 ;
  assign n2891 = ~n2886 & n2890 ;
  assign n2892 = n2883 & n2891 ;
  assign n2893 = \u2_adr0_cnt_reg[9]/P0001  & n1004 ;
  assign n2894 = ~n1799 & ~n2893 ;
  assign n2895 = ~n2204 & ~n2894 ;
  assign n2896 = ~n2209 & n2895 ;
  assign n2897 = \u3_u1_slv_dout_reg[11]/P0001  & n2203 ;
  assign n2898 = n1755 & n2897 ;
  assign n2899 = \u0_u0_ch_adr0_r_reg[9]/P0001  & ~n2204 ;
  assign n2900 = n2209 & n2899 ;
  assign n2901 = ~n2898 & ~n2900 ;
  assign n2902 = ~n2896 & n2901 ;
  assign n2903 = \u2_adr0_cnt_reg[0]/P0001  & n1004 ;
  assign n2904 = ~n1810 & ~n2903 ;
  assign n2905 = ~n2204 & ~n2904 ;
  assign n2906 = ~n2209 & n2905 ;
  assign n2907 = \u3_u1_slv_dout_reg[2]/P0001  & n2203 ;
  assign n2908 = n1755 & n2907 ;
  assign n2909 = \u0_u0_ch_adr0_r_reg[0]/P0001  & ~n2204 ;
  assign n2910 = n2209 & n2909 ;
  assign n2911 = ~n2908 & ~n2910 ;
  assign n2912 = ~n2906 & n2911 ;
  assign n2913 = \u2_adr0_cnt_reg[1]/P0001  & n1004 ;
  assign n2914 = ~n1821 & ~n2913 ;
  assign n2915 = ~n2204 & ~n2914 ;
  assign n2916 = ~n2209 & n2915 ;
  assign n2917 = \u3_u1_slv_dout_reg[3]/P0001  & n2203 ;
  assign n2918 = n1755 & n2917 ;
  assign n2919 = \u0_u0_ch_adr0_r_reg[1]/P0001  & ~n2204 ;
  assign n2920 = n2209 & n2919 ;
  assign n2921 = ~n2918 & ~n2920 ;
  assign n2922 = ~n2916 & n2921 ;
  assign n2923 = \u2_adr0_cnt_reg[2]/P0001  & n1004 ;
  assign n2924 = ~n1832 & ~n2923 ;
  assign n2925 = ~n2204 & ~n2924 ;
  assign n2926 = ~n2209 & n2925 ;
  assign n2927 = \u3_u1_slv_dout_reg[4]/P0001  & n2203 ;
  assign n2928 = n1755 & n2927 ;
  assign n2929 = \u0_u0_ch_adr0_r_reg[2]/P0001  & ~n2204 ;
  assign n2930 = n2209 & n2929 ;
  assign n2931 = ~n2928 & ~n2930 ;
  assign n2932 = ~n2926 & n2931 ;
  assign n2933 = \u2_adr0_cnt_reg[3]/P0001  & n1004 ;
  assign n2934 = ~n1843 & ~n2933 ;
  assign n2935 = ~n2204 & ~n2934 ;
  assign n2936 = ~n2209 & n2935 ;
  assign n2937 = \u3_u1_slv_dout_reg[5]/P0001  & n2203 ;
  assign n2938 = n1755 & n2937 ;
  assign n2939 = \u0_u0_ch_adr0_r_reg[3]/P0001  & ~n2204 ;
  assign n2940 = n2209 & n2939 ;
  assign n2941 = ~n2938 & ~n2940 ;
  assign n2942 = ~n2936 & n2941 ;
  assign n2943 = \u2_adr0_cnt_reg[4]/P0001  & n1004 ;
  assign n2944 = ~n1854 & ~n2943 ;
  assign n2945 = ~n2204 & ~n2944 ;
  assign n2946 = ~n2209 & n2945 ;
  assign n2947 = \u3_u1_slv_dout_reg[6]/P0001  & n2203 ;
  assign n2948 = n1755 & n2947 ;
  assign n2949 = \u0_u0_ch_adr0_r_reg[4]/P0001  & ~n2204 ;
  assign n2950 = n2209 & n2949 ;
  assign n2951 = ~n2948 & ~n2950 ;
  assign n2952 = ~n2946 & n2951 ;
  assign n2953 = \u2_adr0_cnt_reg[5]/P0001  & n1004 ;
  assign n2954 = ~n1865 & ~n2953 ;
  assign n2955 = ~n2204 & ~n2954 ;
  assign n2956 = ~n2209 & n2955 ;
  assign n2957 = \u3_u1_slv_dout_reg[7]/P0001  & n2203 ;
  assign n2958 = n1755 & n2957 ;
  assign n2959 = \u0_u0_ch_adr0_r_reg[5]/P0001  & ~n2204 ;
  assign n2960 = n2209 & n2959 ;
  assign n2961 = ~n2958 & ~n2960 ;
  assign n2962 = ~n2956 & n2961 ;
  assign n2963 = \u2_adr0_cnt_reg[6]/P0001  & n1004 ;
  assign n2964 = ~n1876 & ~n2963 ;
  assign n2965 = ~n2204 & ~n2964 ;
  assign n2966 = ~n2209 & n2965 ;
  assign n2967 = \u3_u1_slv_dout_reg[8]/P0001  & n2203 ;
  assign n2968 = n1755 & n2967 ;
  assign n2969 = \u0_u0_ch_adr0_r_reg[6]/P0001  & ~n2204 ;
  assign n2970 = n2209 & n2969 ;
  assign n2971 = ~n2968 & ~n2970 ;
  assign n2972 = ~n2966 & n2971 ;
  assign n2973 = \u2_adr0_cnt_reg[7]/P0001  & n1004 ;
  assign n2974 = ~n1887 & ~n2973 ;
  assign n2975 = ~n2204 & ~n2974 ;
  assign n2976 = ~n2209 & n2975 ;
  assign n2977 = \u3_u1_slv_dout_reg[9]/P0001  & n2203 ;
  assign n2978 = n1755 & n2977 ;
  assign n2979 = \u0_u0_ch_adr0_r_reg[7]/P0001  & ~n2204 ;
  assign n2980 = n2209 & n2979 ;
  assign n2981 = ~n2978 & ~n2980 ;
  assign n2982 = ~n2976 & n2981 ;
  assign n2983 = \u2_adr0_cnt_reg[8]/P0001  & n1004 ;
  assign n2984 = ~n1788 & ~n2983 ;
  assign n2985 = ~n2204 & ~n2984 ;
  assign n2986 = ~n2209 & n2985 ;
  assign n2987 = \u3_u1_slv_dout_reg[10]/P0001  & n2203 ;
  assign n2988 = n1755 & n2987 ;
  assign n2989 = \u0_u0_ch_adr0_r_reg[8]/P0001  & ~n2204 ;
  assign n2990 = n2209 & n2989 ;
  assign n2991 = ~n2988 & ~n2990 ;
  assign n2992 = ~n2986 & n2991 ;
  assign n2993 = \u0_u0_ch_tot_sz_r_reg[11]/P0001  & n2017 ;
  assign n2994 = \u0_int_maskb_r_reg[11]/NET0131  & n2024 ;
  assign n2995 = \u0_u0_ch_adr0_r_reg[9]/P0001  & n2002 ;
  assign n2996 = ~n1999 & n2995 ;
  assign n2997 = n1994 & n2996 ;
  assign n2998 = ~n2994 & ~n2997 ;
  assign n2999 = ~n2993 & n2998 ;
  assign n3000 = \u0_int_maska_r_reg[11]/NET0131  & n2021 ;
  assign n3001 = ~n2009 & ~n3000 ;
  assign n3002 = \u0_u0_ch_adr1_r_reg[9]/P0001  & n2002 ;
  assign n3003 = n1999 & n3002 ;
  assign n3004 = n1994 & n3003 ;
  assign n3005 = \u0_u0_ch_done_reg/P0002  & n2032 ;
  assign n3006 = ~n3004 & ~n3005 ;
  assign n3007 = n3001 & n3006 ;
  assign n3008 = n2999 & n3007 ;
  assign n3009 = \u0_u0_ch_csr_r2_reg[2]/NET0131  & n2032 ;
  assign n3010 = \u0_int_maska_r_reg[15]/NET0131  & n2021 ;
  assign n3011 = \u0_int_maskb_r_reg[15]/NET0131  & n2024 ;
  assign n3012 = ~n3010 & ~n3011 ;
  assign n3013 = ~n3009 & n3012 ;
  assign n3014 = \u0_u0_ch_adr1_r_reg[13]/P0001  & n2002 ;
  assign n3015 = n1999 & n3014 ;
  assign n3016 = n1994 & n3015 ;
  assign n3017 = ~n2009 & ~n3016 ;
  assign n3018 = \u0_u0_ch_sz_inf_reg/NET0131  & n2017 ;
  assign n3019 = \u0_u0_ch_adr0_r_reg[13]/P0001  & n2002 ;
  assign n3020 = ~n1999 & n3019 ;
  assign n3021 = n1994 & n3020 ;
  assign n3022 = ~n3018 & ~n3021 ;
  assign n3023 = n3017 & n3022 ;
  assign n3024 = n3013 & n3023 ;
  assign n3025 = \u0_int_maskb_r_reg[16]/NET0131  & n2024 ;
  assign n3026 = \u0_u0_rest_en_reg/NET0131  & n2032 ;
  assign n3027 = \u0_int_maska_r_reg[16]/NET0131  & n2021 ;
  assign n3028 = ~n3026 & ~n3027 ;
  assign n3029 = ~n3025 & n3028 ;
  assign n3030 = \u0_u0_ch_adr1_r_reg[14]/P0001  & n2002 ;
  assign n3031 = n1999 & n3030 ;
  assign n3032 = n1994 & n3031 ;
  assign n3033 = ~n2009 & ~n3032 ;
  assign n3034 = \u0_u0_ch_chk_sz_r_reg[0]/P0001  & n2017 ;
  assign n3035 = \u0_u0_ch_adr0_r_reg[14]/P0001  & n2002 ;
  assign n3036 = ~n1999 & n3035 ;
  assign n3037 = n1994 & n3036 ;
  assign n3038 = ~n3034 & ~n3037 ;
  assign n3039 = n3033 & n3038 ;
  assign n3040 = n3029 & n3039 ;
  assign n3041 = \u0_u0_ch_adr1_r_reg[15]/P0001  & n2002 ;
  assign n3042 = n1999 & n3041 ;
  assign n3043 = n1994 & n3042 ;
  assign n3044 = \u0_int_maska_r_reg[17]/NET0131  & n2021 ;
  assign n3045 = \u0_int_maskb_r_reg[17]/NET0131  & n2024 ;
  assign n3046 = ~n3044 & ~n3045 ;
  assign n3047 = ~n3043 & n3046 ;
  assign n3048 = \u0_u0_ch_chk_sz_r_reg[1]/P0001  & n2017 ;
  assign n3049 = ~n2009 & ~n3048 ;
  assign n3050 = \u0_u0_ch_adr0_r_reg[15]/P0001  & n2002 ;
  assign n3051 = ~n1999 & n3050 ;
  assign n3052 = n1994 & n3051 ;
  assign n3053 = \u0_u0_ch_csr_r3_reg[0]/NET0131  & n2032 ;
  assign n3054 = ~n3052 & ~n3053 ;
  assign n3055 = n3049 & n3054 ;
  assign n3056 = n3047 & n3055 ;
  assign n3057 = \u0_u0_ch_adr1_r_reg[16]/P0001  & n2002 ;
  assign n3058 = n1999 & n3057 ;
  assign n3059 = n1994 & n3058 ;
  assign n3060 = \u0_int_maska_r_reg[18]/NET0131  & n2021 ;
  assign n3061 = \u0_int_maskb_r_reg[18]/NET0131  & n2024 ;
  assign n3062 = ~n3060 & ~n3061 ;
  assign n3063 = ~n3059 & n3062 ;
  assign n3064 = \u0_u0_ch_chk_sz_r_reg[2]/P0001  & n2017 ;
  assign n3065 = ~n2009 & ~n3064 ;
  assign n3066 = \u0_u0_ch_adr0_r_reg[16]/P0001  & n2002 ;
  assign n3067 = ~n1999 & n3066 ;
  assign n3068 = n1994 & n3067 ;
  assign n3069 = \u0_u0_ch_csr_r3_reg[1]/NET0131  & n2032 ;
  assign n3070 = ~n3068 & ~n3069 ;
  assign n3071 = n3065 & n3070 ;
  assign n3072 = n3063 & n3071 ;
  assign n3073 = \u0_u0_ch_adr1_r_reg[17]/P0001  & n2002 ;
  assign n3074 = n1999 & n3073 ;
  assign n3075 = n1994 & n3074 ;
  assign n3076 = \u0_int_maska_r_reg[19]/NET0131  & n2021 ;
  assign n3077 = \u0_int_maskb_r_reg[19]/NET0131  & n2024 ;
  assign n3078 = ~n3076 & ~n3077 ;
  assign n3079 = ~n3075 & n3078 ;
  assign n3080 = \u0_u0_ch_chk_sz_r_reg[3]/P0001  & n2017 ;
  assign n3081 = ~n2009 & ~n3080 ;
  assign n3082 = \u0_u0_ch_adr0_r_reg[17]/P0001  & n2002 ;
  assign n3083 = ~n1999 & n3082 ;
  assign n3084 = n1994 & n3083 ;
  assign n3085 = \u0_u0_ch_csr_r3_reg[2]/NET0131  & n2032 ;
  assign n3086 = ~n3084 & ~n3085 ;
  assign n3087 = n3081 & n3086 ;
  assign n3088 = n3079 & n3087 ;
  assign n3089 = \u0_int_maskb_r_reg[20]/NET0131  & n2024 ;
  assign n3090 = \u0_int_maska_r_reg[20]/NET0131  & n2021 ;
  assign n3091 = \u0_u0_ch_adr1_r_reg[18]/P0001  & n2002 ;
  assign n3092 = n1999 & n3091 ;
  assign n3093 = n1994 & n3092 ;
  assign n3094 = ~n3090 & ~n3093 ;
  assign n3095 = ~n3089 & n3094 ;
  assign n3096 = \u0_u0_ch_chk_sz_r_reg[4]/P0001  & n2017 ;
  assign n3097 = \u0_u0_ch_adr0_r_reg[18]/P0001  & n2002 ;
  assign n3098 = ~n1999 & n3097 ;
  assign n3099 = n1994 & n3098 ;
  assign n3100 = ~n3096 & ~n3099 ;
  assign n3101 = n2034 & n3100 ;
  assign n3102 = n3095 & n3101 ;
  assign n3103 = \u0_u0_ch_adr1_r_reg[19]/P0001  & n2002 ;
  assign n3104 = n1999 & n3103 ;
  assign n3105 = n1994 & n3104 ;
  assign n3106 = \u0_int_maska_r_reg[21]/NET0131  & n2021 ;
  assign n3107 = \u0_int_maskb_r_reg[21]/NET0131  & n2024 ;
  assign n3108 = ~n3106 & ~n3107 ;
  assign n3109 = ~n3105 & n3108 ;
  assign n3110 = \u0_u0_ch_chk_sz_r_reg[5]/P0001  & n2017 ;
  assign n3111 = ~n2009 & ~n3110 ;
  assign n3112 = \u0_u0_ch_adr0_r_reg[19]/P0001  & n2002 ;
  assign n3113 = ~n1999 & n3112 ;
  assign n3114 = n1994 & n3113 ;
  assign n3115 = \u0_u0_int_src_r_reg[1]/NET0131  & n2032 ;
  assign n3116 = ~n3114 & ~n3115 ;
  assign n3117 = n3111 & n3116 ;
  assign n3118 = n3109 & n3117 ;
  assign n3119 = \u0_u0_ch_adr1_r_reg[20]/P0001  & n2002 ;
  assign n3120 = n1999 & n3119 ;
  assign n3121 = n1994 & n3120 ;
  assign n3122 = \u0_int_maska_r_reg[22]/NET0131  & n2021 ;
  assign n3123 = \u0_int_maskb_r_reg[22]/NET0131  & n2024 ;
  assign n3124 = ~n3122 & ~n3123 ;
  assign n3125 = ~n3121 & n3124 ;
  assign n3126 = \u0_u0_ch_chk_sz_r_reg[6]/P0001  & n2017 ;
  assign n3127 = ~n2009 & ~n3126 ;
  assign n3128 = \u0_u0_ch_adr0_r_reg[20]/P0001  & n2002 ;
  assign n3129 = ~n1999 & n3128 ;
  assign n3130 = n1994 & n3129 ;
  assign n3131 = \u0_u0_int_src_r_reg[2]/NET0131  & n2032 ;
  assign n3132 = ~n3130 & ~n3131 ;
  assign n3133 = n3127 & n3132 ;
  assign n3134 = n3125 & n3133 ;
  assign n3135 = \u0_u0_ch_adr0_r_reg[2]/P0001  & n2002 ;
  assign n3136 = ~n1999 & n3135 ;
  assign n3137 = n1994 & n3136 ;
  assign n3138 = \u0_int_maska_r_reg[4]/NET0131  & n2021 ;
  assign n3139 = \u0_int_maskb_r_reg[4]/NET0131  & n2024 ;
  assign n3140 = ~n3138 & ~n3139 ;
  assign n3141 = ~n3137 & n3140 ;
  assign n3142 = \u0_u0_ch_csr_r_reg[4]/NET0131  & n2032 ;
  assign n3143 = ~n2009 & ~n3142 ;
  assign n3144 = \u0_u0_ch_adr1_r_reg[2]/P0001  & n2002 ;
  assign n3145 = n1999 & n3144 ;
  assign n3146 = n1994 & n3145 ;
  assign n3147 = \u0_u0_ch_tot_sz_r_reg[4]/P0001  & n2017 ;
  assign n3148 = ~n3146 & ~n3147 ;
  assign n3149 = n3143 & n3148 ;
  assign n3150 = n3141 & n3149 ;
  assign n3151 = \u0_u0_ch_tot_sz_r_reg[5]/P0001  & n2017 ;
  assign n3152 = \u0_u0_ch_adr0_r_reg[3]/P0001  & n2002 ;
  assign n3153 = ~n1999 & n3152 ;
  assign n3154 = n1994 & n3153 ;
  assign n3155 = \u0_int_maskb_r_reg[5]/NET0131  & n2024 ;
  assign n3156 = ~n3154 & ~n3155 ;
  assign n3157 = ~n3151 & n3156 ;
  assign n3158 = \u0_u0_ch_csr_r_reg[5]/NET0131  & n2032 ;
  assign n3159 = ~n2009 & ~n3158 ;
  assign n3160 = \u0_u0_ch_adr1_r_reg[3]/P0001  & n2002 ;
  assign n3161 = n1999 & n3160 ;
  assign n3162 = n1994 & n3161 ;
  assign n3163 = \u0_int_maska_r_reg[5]/NET0131  & n2021 ;
  assign n3164 = ~n3162 & ~n3163 ;
  assign n3165 = n3159 & n3164 ;
  assign n3166 = n3157 & n3165 ;
  assign n3167 = \u0_u0_ch_tot_sz_r_reg[6]/P0001  & n2017 ;
  assign n3168 = \u0_u0_ch_adr0_r_reg[4]/P0001  & n2002 ;
  assign n3169 = ~n1999 & n3168 ;
  assign n3170 = n1994 & n3169 ;
  assign n3171 = \u0_int_maskb_r_reg[6]/NET0131  & n2024 ;
  assign n3172 = ~n3170 & ~n3171 ;
  assign n3173 = ~n3167 & n3172 ;
  assign n3174 = \u0_u0_ch_csr_r_reg[6]/NET0131  & n2032 ;
  assign n3175 = ~n2009 & ~n3174 ;
  assign n3176 = \u0_u0_ch_adr1_r_reg[4]/P0001  & n2002 ;
  assign n3177 = n1999 & n3176 ;
  assign n3178 = n1994 & n3177 ;
  assign n3179 = \u0_int_maska_r_reg[6]/NET0131  & n2021 ;
  assign n3180 = ~n3178 & ~n3179 ;
  assign n3181 = n3175 & n3180 ;
  assign n3182 = n3173 & n3181 ;
  assign n3183 = \u0_u0_ch_tot_sz_r_reg[7]/P0001  & n2017 ;
  assign n3184 = \u0_u0_ch_adr0_r_reg[5]/P0001  & n2002 ;
  assign n3185 = ~n1999 & n3184 ;
  assign n3186 = n1994 & n3185 ;
  assign n3187 = \u0_int_maskb_r_reg[7]/NET0131  & n2024 ;
  assign n3188 = ~n3186 & ~n3187 ;
  assign n3189 = ~n3183 & n3188 ;
  assign n3190 = \u0_u0_ch_csr_r_reg[7]/NET0131  & n2032 ;
  assign n3191 = ~n2009 & ~n3190 ;
  assign n3192 = \u0_u0_ch_adr1_r_reg[5]/P0001  & n2002 ;
  assign n3193 = n1999 & n3192 ;
  assign n3194 = n1994 & n3193 ;
  assign n3195 = \u0_int_maska_r_reg[7]/NET0131  & n2021 ;
  assign n3196 = ~n3194 & ~n3195 ;
  assign n3197 = n3191 & n3196 ;
  assign n3198 = n3189 & n3197 ;
  assign n3199 = \u0_u0_ch_tot_sz_r_reg[8]/P0001  & n2017 ;
  assign n3200 = \u0_int_maskb_r_reg[8]/NET0131  & n2024 ;
  assign n3201 = \u0_u0_ch_adr0_r_reg[6]/P0001  & n2002 ;
  assign n3202 = ~n1999 & n3201 ;
  assign n3203 = n1994 & n3202 ;
  assign n3204 = ~n3200 & ~n3203 ;
  assign n3205 = ~n3199 & n3204 ;
  assign n3206 = \u0_int_maska_r_reg[8]/NET0131  & n2021 ;
  assign n3207 = ~n2009 & ~n3206 ;
  assign n3208 = \u0_u0_ch_adr1_r_reg[6]/P0001  & n2002 ;
  assign n3209 = n1999 & n3208 ;
  assign n3210 = n1994 & n3209 ;
  assign n3211 = \u0_u0_ch_csr_r_reg[8]/NET0131  & n2032 ;
  assign n3212 = ~n3210 & ~n3211 ;
  assign n3213 = n3207 & n3212 ;
  assign n3214 = n3205 & n3213 ;
  assign n3215 = \u0_u0_ch_adr0_r_reg[29]/P0001  & n2002 ;
  assign n3216 = ~n1999 & n3215 ;
  assign n3217 = n1994 & n3216 ;
  assign n3218 = \u0_u0_ch_adr1_r_reg[29]/P0001  & n2002 ;
  assign n3219 = n1999 & n3218 ;
  assign n3220 = n1994 & n3219 ;
  assign n3221 = ~n2009 & ~n3220 ;
  assign n3222 = ~n3217 & n3221 ;
  assign n3223 = \u0_u0_ch_csr_r_reg[1]/NET0131  & n2032 ;
  assign n3224 = \u0_u0_ch_tot_sz_r_reg[1]/P0001  & n2017 ;
  assign n3225 = ~n3223 & ~n3224 ;
  assign n3226 = \u0_int_maska_r_reg[1]/NET0131  & n2021 ;
  assign n3227 = \u0_int_maskb_r_reg[1]/NET0131  & n2024 ;
  assign n3228 = ~n3226 & ~n3227 ;
  assign n3229 = n3225 & n3228 ;
  assign n3230 = ~\u0_u0_ch_err_reg/NET0131  & ~\u2_dma_abort_r_reg/NET0131  ;
  assign n3231 = ~\u2_dma_abort_r_reg/NET0131  & n1425 ;
  assign n3232 = n1424 & n3231 ;
  assign n3233 = ~n3230 & ~n3232 ;
  assign n3234 = ~\u2_adr0_cnt_reg[15]/P0001  & ~n2163 ;
  assign n3235 = ~n2164 & ~n3234 ;
  assign n3236 = ~\u2_adr1_cnt_reg[15]/P0001  & ~n2167 ;
  assign n3237 = ~n2168 & ~n3236 ;
  assign n3238 = \u2_adr0_cnt_reg[10]/P0001  & n1963 ;
  assign n3239 = ~\u2_adr0_cnt_reg[11]/P0001  & ~n3238 ;
  assign n3240 = ~n1965 & ~n3239 ;
  assign n3241 = \u2_adr1_cnt_reg[10]/P0001  & n1979 ;
  assign n3242 = ~\u2_adr1_cnt_reg[11]/P0001  & ~n3241 ;
  assign n3243 = ~n1981 & ~n3242 ;
  assign n3244 = \u2_adr0_cnt_reg[4]/P0001  & n1957 ;
  assign n3245 = ~\u2_adr0_cnt_reg[4]/P0001  & ~n1957 ;
  assign n3246 = ~n3244 & ~n3245 ;
  assign n3247 = \u2_adr1_cnt_reg[4]/P0001  & n1973 ;
  assign n3248 = ~\u2_adr1_cnt_reg[4]/P0001  & ~n1973 ;
  assign n3249 = ~n3247 & ~n3248 ;
  assign n3250 = ~\u0_u0_ch_stop_reg/P0001  & ~\wb0_err_i_pad  ;
  assign n3251 = ~\wb1_err_i_pad  & n3250 ;
  assign n3252 = ~\u2_state_reg[7]/NET0131  & ~\wb0_ack_i_pad  ;
  assign n3253 = n1511 & ~n3252 ;
  assign n3254 = n1513 & n3253 ;
  assign n3255 = \u2_state_reg[7]/NET0131  & ~\u2_state_reg[9]/NET0131  ;
  assign n3256 = n948 & n3255 ;
  assign n3257 = ~\wb0_ack_i_pad  & n3256 ;
  assign n3258 = n1385 & n3257 ;
  assign n3259 = ~n3254 & ~n3258 ;
  assign n3260 = ~\u2_state_reg[5]/NET0131  & ~\wb0_ack_i_pad  ;
  assign n3261 = \u2_state_reg[5]/NET0131  & n956 ;
  assign n3262 = n953 & n3261 ;
  assign n3263 = n950 & n3252 ;
  assign n3264 = n3262 & n3263 ;
  assign n3265 = ~n1655 & ~n3264 ;
  assign n3266 = ~n3260 & ~n3265 ;
  assign n3267 = \wb0_ack_i_pad  & n3256 ;
  assign n3268 = n1385 & n3267 ;
  assign n3269 = ~\u2_state_reg[6]/NET0131  & ~\wb0_ack_i_pad  ;
  assign n3270 = ~\u2_state_reg[7]/NET0131  & ~n3269 ;
  assign n3271 = n950 & n3270 ;
  assign n3272 = n3262 & n3271 ;
  assign n3273 = ~\wb0_ack_i_pad  & n1511 ;
  assign n3274 = n1513 & n3273 ;
  assign n3275 = ~n3272 & ~n3274 ;
  assign n3276 = \u2_adr0_cnt_reg[10]/P0001  & \u2_adr0_cnt_reg[13]/P0001  ;
  assign n3277 = n1967 & n3276 ;
  assign n3278 = n1963 & n3277 ;
  assign n3279 = ~\u2_adr0_cnt_reg[14]/P0001  & ~n3278 ;
  assign n3280 = ~n2163 & ~n3279 ;
  assign n3281 = \u2_adr1_cnt_reg[10]/P0001  & \u2_adr1_cnt_reg[13]/P0001  ;
  assign n3282 = n1983 & n3281 ;
  assign n3283 = n1979 & n3282 ;
  assign n3284 = ~\u2_adr1_cnt_reg[14]/P0001  & ~n3283 ;
  assign n3285 = ~n2167 & ~n3284 ;
  assign n3286 = ~\u2_adr0_cnt_reg[7]/P0001  & ~n1960 ;
  assign n3287 = ~n2195 & ~n3286 ;
  assign n3288 = ~\u2_adr1_cnt_reg[7]/P0001  & ~n1976 ;
  assign n3289 = ~n2200 & ~n3288 ;
  assign n3290 = ~\u4_u1_rf_ack_reg/P0001  & \wb1_stb_i_pad  ;
  assign n3291 = ~\u4_u1_slv_re_reg/P0001  & ~\u4_u1_slv_we_reg/P0001  ;
  assign n3292 = \wb1_cyc_i_pad  & ~n3291 ;
  assign n3293 = n3290 & n3292 ;
  assign n3294 = n917 & n919 ;
  assign n3295 = \u0_u0_ch_csr_r_reg[5]/NET0131  & ~n1362 ;
  assign n3296 = \u3_u1_slv_dout_reg[5]/P0001  & n1359 ;
  assign n3297 = n1358 & n3296 ;
  assign n3298 = ~n3295 & ~n3297 ;
  assign n3299 = \u0_u0_ch_csr_r_reg[6]/NET0131  & ~n1362 ;
  assign n3300 = \u3_u1_slv_dout_reg[6]/P0001  & n1359 ;
  assign n3301 = n1358 & n3300 ;
  assign n3302 = ~n3299 & ~n3301 ;
  assign n3303 = \u0_u0_ch_csr_r_reg[7]/NET0131  & ~n1362 ;
  assign n3304 = \u3_u1_slv_dout_reg[7]/P0001  & n1359 ;
  assign n3305 = n1358 & n3304 ;
  assign n3306 = ~n3303 & ~n3305 ;
  assign n3307 = \u0_u0_ch_csr_r_reg[8]/NET0131  & ~n1362 ;
  assign n3308 = \u3_u1_slv_dout_reg[8]/P0001  & n1359 ;
  assign n3309 = n1358 & n3308 ;
  assign n3310 = ~n3307 & ~n3309 ;
  assign n3311 = \u3_u1_slv_dout_reg[9]/P0001  & n1359 ;
  assign n3312 = n1358 & n3311 ;
  assign n3313 = \u2_adr1_cnt_reg[2]/P0001  & n1971 ;
  assign n3314 = ~\u2_adr1_cnt_reg[3]/P0001  & ~n3313 ;
  assign n3315 = ~n1973 & ~n3314 ;
  assign n3316 = ~\u3_u1_slv_adr_reg[5]/P0001  & n1359 ;
  assign n3317 = n1355 & n3316 ;
  assign n3318 = n1756 & n3317 ;
  assign n3319 = \u0_int_maska_r_reg[0]/NET0131  & ~n3318 ;
  assign n3320 = n1772 & n3317 ;
  assign n3321 = ~n3319 & ~n3320 ;
  assign n3322 = \u0_int_maska_r_reg[10]/NET0131  & ~n3318 ;
  assign n3323 = n1792 & n3317 ;
  assign n3324 = ~n3322 & ~n3323 ;
  assign n3325 = \u0_int_maska_r_reg[11]/NET0131  & ~n3318 ;
  assign n3326 = n1803 & n3317 ;
  assign n3327 = ~n3325 & ~n3326 ;
  assign n3328 = \u0_int_maska_r_reg[8]/NET0131  & ~n3318 ;
  assign n3329 = n1880 & n3317 ;
  assign n3330 = ~n3328 & ~n3329 ;
  assign n3331 = \u0_int_maska_r_reg[5]/NET0131  & ~n3318 ;
  assign n3332 = n1847 & n3317 ;
  assign n3333 = ~n3331 & ~n3332 ;
  assign n3334 = \u0_int_maska_r_reg[6]/NET0131  & ~n3318 ;
  assign n3335 = n1858 & n3317 ;
  assign n3336 = ~n3334 & ~n3335 ;
  assign n3337 = \u0_int_maska_r_reg[7]/NET0131  & ~n3318 ;
  assign n3338 = n1869 & n3317 ;
  assign n3339 = ~n3337 & ~n3338 ;
  assign n3340 = \u0_int_maska_r_reg[9]/NET0131  & ~n3318 ;
  assign n3341 = n1891 & n3317 ;
  assign n3342 = ~n3340 & ~n3341 ;
  assign n3343 = \u3_u1_slv_dout_reg[0]/P0001  & n1356 ;
  assign n3344 = n3317 & n3343 ;
  assign n3345 = n1356 & n3317 ;
  assign n3346 = \u0_csr_r_reg[0]/NET0131  & ~n3345 ;
  assign n3347 = ~n3344 & ~n3346 ;
  assign n3348 = \u2_adr0_cnt_reg[2]/P0001  & n1955 ;
  assign n3349 = ~\u2_adr0_cnt_reg[3]/P0001  & ~n3348 ;
  assign n3350 = ~n1957 & ~n3349 ;
  assign n3351 = ~\u2_adr1_cnt_reg[10]/P0001  & ~n1979 ;
  assign n3352 = ~n3241 & ~n3351 ;
  assign n3353 = ~\u2_adr0_cnt_reg[10]/P0001  & ~n1963 ;
  assign n3354 = ~n3238 & ~n3353 ;
  assign n3355 = \u2_adr0_cnt_reg[4]/P0001  & \u2_adr0_cnt_reg[5]/P0001  ;
  assign n3356 = n1957 & n3355 ;
  assign n3357 = ~\u2_adr0_cnt_reg[6]/P0001  & ~n3356 ;
  assign n3358 = ~n1960 & ~n3357 ;
  assign n3359 = ~\u2_adr0_cnt_reg[13]/P0001  & ~n1969 ;
  assign n3360 = ~n3278 & ~n3359 ;
  assign n3361 = ~\u2_adr1_cnt_reg[13]/P0001  & ~n1985 ;
  assign n3362 = ~n3283 & ~n3361 ;
  assign n3363 = \u2_adr1_cnt_reg[4]/P0001  & \u2_adr1_cnt_reg[5]/P0001  ;
  assign n3364 = n1973 & n3363 ;
  assign n3365 = ~\u2_adr1_cnt_reg[6]/P0001  & ~n3364 ;
  assign n3366 = ~n1976 & ~n3365 ;
  assign n3367 = n2203 & n3317 ;
  assign n3368 = \u0_int_maskb_r_reg[11]/NET0131  & ~n3367 ;
  assign n3369 = n2897 & n3317 ;
  assign n3370 = ~n3368 & ~n3369 ;
  assign n3371 = \u0_int_maskb_r_reg[10]/NET0131  & ~n3367 ;
  assign n3372 = n2987 & n3317 ;
  assign n3373 = ~n3371 & ~n3372 ;
  assign n3374 = \u0_int_maskb_r_reg[0]/NET0131  & ~n3367 ;
  assign n3375 = \u3_u1_slv_dout_reg[0]/P0001  & n2203 ;
  assign n3376 = n3317 & n3375 ;
  assign n3377 = ~n3374 & ~n3376 ;
  assign n3378 = \u0_int_maskb_r_reg[5]/NET0131  & ~n3367 ;
  assign n3379 = n2937 & n3317 ;
  assign n3380 = ~n3378 & ~n3379 ;
  assign n3381 = \u0_int_maskb_r_reg[6]/NET0131  & ~n3367 ;
  assign n3382 = n2947 & n3317 ;
  assign n3383 = ~n3381 & ~n3382 ;
  assign n3384 = \u0_int_maskb_r_reg[7]/NET0131  & ~n3367 ;
  assign n3385 = n2957 & n3317 ;
  assign n3386 = ~n3384 & ~n3385 ;
  assign n3387 = \u0_int_maskb_r_reg[8]/NET0131  & ~n3367 ;
  assign n3388 = n2967 & n3317 ;
  assign n3389 = ~n3387 & ~n3388 ;
  assign n3390 = \u0_int_maskb_r_reg[9]/NET0131  & ~n3367 ;
  assign n3391 = n2977 & n3317 ;
  assign n3392 = ~n3390 & ~n3391 ;
  assign n3393 = ~\u2_adr0_cnt_reg[9]/P0001  & ~n2194 ;
  assign n3394 = ~n1963 & ~n3393 ;
  assign n3395 = ~\u2_adr1_cnt_reg[9]/P0001  & ~n2199 ;
  assign n3396 = ~n1979 & ~n3395 ;
  assign n3397 = ~\wb1_addr_i[28]_pad  & ~\wb1_addr_i[29]_pad  ;
  assign n3398 = ~\wb1_addr_i[30]_pad  & ~\wb1_addr_i[31]_pad  ;
  assign n3399 = n3397 & n3398 ;
  assign n3400 = \wb1_cyc_i_pad  & n3399 ;
  assign n3401 = ~\u4_u1_slv_re_reg/P0001  & ~\wb1_we_i_pad  ;
  assign n3402 = n3290 & n3401 ;
  assign n3403 = n3400 & n3402 ;
  assign n3404 = ~\wb0_addr_i[28]_pad  & ~\wb0_addr_i[29]_pad  ;
  assign n3405 = ~\wb0_addr_i[30]_pad  & ~\wb0_addr_i[31]_pad  ;
  assign n3406 = n3404 & n3405 ;
  assign n3407 = ~\u3_u1_rf_ack_reg/P0001  & \wb0_cyc_i_pad  ;
  assign n3408 = \wb0_stb_i_pad  & n3407 ;
  assign n3409 = ~\u3_u1_slv_re_reg/P0001  & ~\wb0_we_i_pad  ;
  assign n3410 = n3408 & n3409 ;
  assign n3411 = n3406 & n3410 ;
  assign n3412 = \wb1_cyc_i_pad  & \wb1_we_i_pad  ;
  assign n3413 = n3290 & n3412 ;
  assign n3414 = n3399 & n3413 ;
  assign n3415 = ~\u2_adr0_cnt_reg[5]/P0001  & ~n3244 ;
  assign n3416 = ~n3356 & ~n3415 ;
  assign n3417 = ~\u2_adr1_cnt_reg[5]/P0001  & ~n3247 ;
  assign n3418 = ~n3364 & ~n3417 ;
  assign n3419 = \wb0_stb_i_pad  & \wb0_we_i_pad  ;
  assign n3420 = n3407 & n3419 ;
  assign n3421 = n3406 & n3420 ;
  assign n3422 = ~\u2_adr0_cnt_reg[2]/P0001  & ~n1955 ;
  assign n3423 = ~n3348 & ~n3422 ;
  assign n3424 = ~\u2_adr1_cnt_reg[2]/P0001  & ~n1971 ;
  assign n3425 = ~n3313 & ~n3424 ;
  assign n3426 = \u0_u0_ch_csr_r_reg[0]/NET0131  & ~n753 ;
  assign n3427 = ~\u3_u1_slv_re_reg/P0001  & ~\u3_u1_slv_we_reg/P0001  ;
  assign n3428 = n3408 & ~n3427 ;
  assign n3429 = ~\u2_adr0_cnt_reg[0]/P0001  & ~\u2_adr0_cnt_reg[1]/P0001  ;
  assign n3430 = ~n1955 & ~n3429 ;
  assign n3431 = ~\u2_adr1_cnt_reg[0]/P0001  & ~\u2_adr1_cnt_reg[1]/P0001  ;
  assign n3432 = ~n1971 & ~n3431 ;
  assign n3433 = dma_nd_i_pad & ~dma_req_i_pad ;
  assign n3434 = ~dma_ack_o_pad & dma_req_i_pad ;
  assign n3435 = dma_nd_i_pad & dma_req_i_pad ;
  assign n3436 = \u2_tsz_cnt_reg[2]/NET0131  & ~n1664 ;
  assign n3437 = ~n1691 & ~n3436 ;
  assign n3438 = n757 & ~n3437 ;
  assign n3439 = \u0_u0_ch_tot_sz_r_reg[2]/P0001  & ~n757 ;
  assign n3440 = ~n3438 & ~n3439 ;
  assign n3441 = \u0_u0_ch_adr1_r_reg[25]/P0001  & ~n757 ;
  assign n3442 = ~\u2_adr1_cnt_reg[25]/P0001  & ~n831 ;
  assign n3443 = n757 & ~n806 ;
  assign n3444 = ~n3442 & n3443 ;
  assign n3445 = ~n3441 & ~n3444 ;
  assign n3446 = \u2_adr0_cnt_reg[13]/P0001  & ~n1036 ;
  assign n3447 = \u2_u0_out_r_reg[13]/P0001  & n768 ;
  assign n3448 = ~n767 & n3447 ;
  assign n3449 = ~n3446 & ~n3448 ;
  assign n3450 = n757 & ~n3449 ;
  assign n3451 = \u0_u0_ch_adr0_r_reg[13]/P0001  & ~n757 ;
  assign n3452 = ~n3450 & ~n3451 ;
  assign n3453 = \u0_u0_ch_tot_sz_r_reg[10]/P0001  & n2017 ;
  assign n3454 = \u0_int_maskb_r_reg[10]/NET0131  & n2024 ;
  assign n3455 = \u0_u0_ch_busy_reg/P0001  & n2032 ;
  assign n3456 = ~n3454 & ~n3455 ;
  assign n3457 = ~n3453 & n3456 ;
  assign n3458 = \u0_int_maska_r_reg[10]/NET0131  & n2021 ;
  assign n3459 = ~n2009 & ~n3458 ;
  assign n3460 = \u0_u0_ch_adr0_r_reg[8]/P0001  & n2002 ;
  assign n3461 = ~n1999 & n3460 ;
  assign n3462 = n1994 & n3461 ;
  assign n3463 = \u0_u0_ch_adr1_r_reg[8]/P0001  & n2002 ;
  assign n3464 = n1999 & n3463 ;
  assign n3465 = n1994 & n3464 ;
  assign n3466 = ~n3462 & ~n3465 ;
  assign n3467 = n3459 & n3466 ;
  assign n3468 = n3457 & n3467 ;
  assign n3469 = \u0_u0_ch_done_reg/P0002  & ~n1362 ;
  assign n3470 = ~n1372 & ~n3469 ;
  assign n3471 = ~n1361 & n3470 ;
  assign n3472 = ~n1000 & n1008 ;
  assign n3473 = ~n970 & ~n3472 ;
  assign n3474 = \wb0_cyc_i_pad  & ~n3406 ;
  assign n3475 = \u3_u1_rf_ack_reg/P0001  & ~n3474 ;
  assign n3476 = \wb0_cyc_i_pad  & \wb1_ack_i_pad  ;
  assign n3477 = ~n3406 & n3476 ;
  assign n3478 = ~n3475 & ~n3477 ;
  assign n3479 = \wb1_addr_i[0]_pad  & \wb1_cyc_i_pad  ;
  assign n3480 = ~n3399 & n3479 ;
  assign n3481 = \wb1_cyc_i_pad  & ~n3399 ;
  assign n3482 = \u2_mast0_adr_reg[10]/P0001  & ~n3481 ;
  assign n3483 = \wb1_addr_i[10]_pad  & \wb1_cyc_i_pad  ;
  assign n3484 = ~n3399 & n3483 ;
  assign n3485 = ~n3482 & ~n3484 ;
  assign n3486 = \u2_mast0_adr_reg[11]/P0001  & ~n3481 ;
  assign n3487 = \wb1_addr_i[11]_pad  & \wb1_cyc_i_pad  ;
  assign n3488 = ~n3399 & n3487 ;
  assign n3489 = ~n3486 & ~n3488 ;
  assign n3490 = \u2_mast0_adr_reg[12]/P0001  & ~n3481 ;
  assign n3491 = \wb1_addr_i[12]_pad  & \wb1_cyc_i_pad  ;
  assign n3492 = ~n3399 & n3491 ;
  assign n3493 = ~n3490 & ~n3492 ;
  assign n3494 = \u2_mast0_adr_reg[13]/P0001  & ~n3481 ;
  assign n3495 = \wb1_addr_i[13]_pad  & \wb1_cyc_i_pad  ;
  assign n3496 = ~n3399 & n3495 ;
  assign n3497 = ~n3494 & ~n3496 ;
  assign n3498 = \u2_mast0_adr_reg[14]/P0001  & ~n3481 ;
  assign n3499 = \wb1_addr_i[14]_pad  & \wb1_cyc_i_pad  ;
  assign n3500 = ~n3399 & n3499 ;
  assign n3501 = ~n3498 & ~n3500 ;
  assign n3502 = \u2_mast0_adr_reg[15]/P0001  & ~n3481 ;
  assign n3503 = \wb1_addr_i[15]_pad  & \wb1_cyc_i_pad  ;
  assign n3504 = ~n3399 & n3503 ;
  assign n3505 = ~n3502 & ~n3504 ;
  assign n3506 = \u2_mast0_adr_reg[16]/P0001  & ~n3481 ;
  assign n3507 = \wb1_addr_i[16]_pad  & \wb1_cyc_i_pad  ;
  assign n3508 = ~n3399 & n3507 ;
  assign n3509 = ~n3506 & ~n3508 ;
  assign n3510 = \u2_mast0_adr_reg[17]/P0001  & ~n3481 ;
  assign n3511 = \wb1_addr_i[17]_pad  & \wb1_cyc_i_pad  ;
  assign n3512 = ~n3399 & n3511 ;
  assign n3513 = ~n3510 & ~n3512 ;
  assign n3514 = \u2_mast0_adr_reg[18]/P0001  & ~n3481 ;
  assign n3515 = \wb1_addr_i[18]_pad  & \wb1_cyc_i_pad  ;
  assign n3516 = ~n3399 & n3515 ;
  assign n3517 = ~n3514 & ~n3516 ;
  assign n3518 = \u2_mast0_adr_reg[19]/P0001  & ~n3481 ;
  assign n3519 = \wb1_addr_i[19]_pad  & \wb1_cyc_i_pad  ;
  assign n3520 = ~n3399 & n3519 ;
  assign n3521 = ~n3518 & ~n3520 ;
  assign n3522 = \wb1_addr_i[1]_pad  & \wb1_cyc_i_pad  ;
  assign n3523 = ~n3399 & n3522 ;
  assign n3524 = \u2_mast0_adr_reg[20]/P0001  & ~n3481 ;
  assign n3525 = \wb1_addr_i[20]_pad  & \wb1_cyc_i_pad  ;
  assign n3526 = ~n3399 & n3525 ;
  assign n3527 = ~n3524 & ~n3526 ;
  assign n3528 = \u2_mast0_adr_reg[21]/P0001  & ~n3481 ;
  assign n3529 = \wb1_addr_i[21]_pad  & \wb1_cyc_i_pad  ;
  assign n3530 = ~n3399 & n3529 ;
  assign n3531 = ~n3528 & ~n3530 ;
  assign n3532 = \u2_mast0_adr_reg[22]/P0001  & ~n3481 ;
  assign n3533 = \wb1_addr_i[22]_pad  & \wb1_cyc_i_pad  ;
  assign n3534 = ~n3399 & n3533 ;
  assign n3535 = ~n3532 & ~n3534 ;
  assign n3536 = \u2_mast0_adr_reg[23]/P0001  & ~n3481 ;
  assign n3537 = \wb1_addr_i[23]_pad  & \wb1_cyc_i_pad  ;
  assign n3538 = ~n3399 & n3537 ;
  assign n3539 = ~n3536 & ~n3538 ;
  assign n3540 = \u2_mast0_adr_reg[24]/P0001  & ~n3481 ;
  assign n3541 = \wb1_addr_i[24]_pad  & \wb1_cyc_i_pad  ;
  assign n3542 = ~n3399 & n3541 ;
  assign n3543 = ~n3540 & ~n3542 ;
  assign n3544 = \u2_mast0_adr_reg[25]/P0001  & ~n3481 ;
  assign n3545 = \wb1_addr_i[25]_pad  & \wb1_cyc_i_pad  ;
  assign n3546 = ~n3399 & n3545 ;
  assign n3547 = ~n3544 & ~n3546 ;
  assign n3548 = \u2_mast0_adr_reg[26]/P0001  & ~n3481 ;
  assign n3549 = \wb1_addr_i[26]_pad  & \wb1_cyc_i_pad  ;
  assign n3550 = ~n3399 & n3549 ;
  assign n3551 = ~n3548 & ~n3550 ;
  assign n3552 = \u2_mast0_adr_reg[27]/P0001  & ~n3481 ;
  assign n3553 = \wb1_addr_i[27]_pad  & \wb1_cyc_i_pad  ;
  assign n3554 = ~n3399 & n3553 ;
  assign n3555 = ~n3552 & ~n3554 ;
  assign n3556 = \wb1_addr_i[28]_pad  & \wb1_cyc_i_pad  ;
  assign n3557 = ~\u2_mast0_adr_reg[28]/P0001  & ~n3556 ;
  assign n3558 = \wb1_cyc_i_pad  & ~n3556 ;
  assign n3559 = ~n3399 & n3558 ;
  assign n3560 = ~n3557 & ~n3559 ;
  assign n3561 = \wb1_addr_i[29]_pad  & \wb1_cyc_i_pad  ;
  assign n3562 = ~\u2_mast0_adr_reg[29]/P0001  & ~n3561 ;
  assign n3563 = \wb1_cyc_i_pad  & ~n3561 ;
  assign n3564 = ~n3399 & n3563 ;
  assign n3565 = ~n3562 & ~n3564 ;
  assign n3566 = \u2_mast0_adr_reg[2]/P0001  & ~n3481 ;
  assign n3567 = \wb1_addr_i[2]_pad  & \wb1_cyc_i_pad  ;
  assign n3568 = ~n3399 & n3567 ;
  assign n3569 = ~n3566 & ~n3568 ;
  assign n3570 = \wb1_addr_i[30]_pad  & \wb1_cyc_i_pad  ;
  assign n3571 = ~\u2_mast0_adr_reg[30]/P0001  & ~n3570 ;
  assign n3572 = \wb1_cyc_i_pad  & ~n3570 ;
  assign n3573 = ~n3399 & n3572 ;
  assign n3574 = ~n3571 & ~n3573 ;
  assign n3575 = \wb1_addr_i[31]_pad  & \wb1_cyc_i_pad  ;
  assign n3576 = ~\u2_mast0_adr_reg[31]/P0001  & ~n3575 ;
  assign n3577 = \wb1_cyc_i_pad  & ~n3575 ;
  assign n3578 = ~n3399 & n3577 ;
  assign n3579 = ~n3576 & ~n3578 ;
  assign n3580 = \u2_mast0_adr_reg[3]/NET0131  & ~n3481 ;
  assign n3581 = \wb1_addr_i[3]_pad  & \wb1_cyc_i_pad  ;
  assign n3582 = ~n3399 & n3581 ;
  assign n3583 = ~n3580 & ~n3582 ;
  assign n3584 = \u2_mast0_adr_reg[4]/P0001  & ~n3481 ;
  assign n3585 = \wb1_addr_i[4]_pad  & \wb1_cyc_i_pad  ;
  assign n3586 = ~n3399 & n3585 ;
  assign n3587 = ~n3584 & ~n3586 ;
  assign n3588 = \u2_mast0_adr_reg[5]/P0001  & ~n3481 ;
  assign n3589 = \wb1_addr_i[5]_pad  & \wb1_cyc_i_pad  ;
  assign n3590 = ~n3399 & n3589 ;
  assign n3591 = ~n3588 & ~n3590 ;
  assign n3592 = \u2_mast0_adr_reg[6]/P0001  & ~n3481 ;
  assign n3593 = \wb1_addr_i[6]_pad  & \wb1_cyc_i_pad  ;
  assign n3594 = ~n3399 & n3593 ;
  assign n3595 = ~n3592 & ~n3594 ;
  assign n3596 = \u2_mast0_adr_reg[7]/P0001  & ~n3481 ;
  assign n3597 = \wb1_addr_i[7]_pad  & \wb1_cyc_i_pad  ;
  assign n3598 = ~n3399 & n3597 ;
  assign n3599 = ~n3596 & ~n3598 ;
  assign n3600 = \u2_mast0_adr_reg[8]/P0001  & ~n3481 ;
  assign n3601 = \wb1_addr_i[8]_pad  & \wb1_cyc_i_pad  ;
  assign n3602 = ~n3399 & n3601 ;
  assign n3603 = ~n3600 & ~n3602 ;
  assign n3604 = \u2_mast0_adr_reg[9]/P0001  & ~n3481 ;
  assign n3605 = \wb1_addr_i[9]_pad  & \wb1_cyc_i_pad  ;
  assign n3606 = ~n3399 & n3605 ;
  assign n3607 = ~n3604 & ~n3606 ;
  assign n3608 = ~\u3_u0_mast_cyc_reg/P0001  & ~n3481 ;
  assign n3609 = \wb0_cyc_i_pad  & \wb1_err_i_pad  ;
  assign n3610 = ~n3406 & n3609 ;
  assign n3611 = \wb0_cyc_i_pad  & \wb1_rty_i_pad  ;
  assign n3612 = ~n3406 & n3611 ;
  assign n3613 = \wb1_cyc_i_pad  & ~\wb1_sel_i[0]_pad  ;
  assign n3614 = ~n3399 & n3613 ;
  assign n3615 = \wb1_cyc_i_pad  & ~\wb1_sel_i[1]_pad  ;
  assign n3616 = ~n3399 & n3615 ;
  assign n3617 = \wb1_cyc_i_pad  & ~\wb1_sel_i[2]_pad  ;
  assign n3618 = ~n3399 & n3617 ;
  assign n3619 = \wb1_cyc_i_pad  & ~\wb1_sel_i[3]_pad  ;
  assign n3620 = ~n3399 & n3619 ;
  assign n3621 = \u3_u0_mast_stb_reg/P0001  & ~n3481 ;
  assign n3622 = \wb1_cyc_i_pad  & \wb1_stb_i_pad  ;
  assign n3623 = ~n3399 & n3622 ;
  assign n3624 = ~n3621 & ~n3623 ;
  assign n3625 = \u3_u0_mast_we_r_reg/P0002  & ~n3481 ;
  assign n3626 = ~n3399 & n3412 ;
  assign n3627 = ~n3625 & ~n3626 ;
  assign n3628 = \u0_wb_rf_dout_reg[0]/P0001  & ~n3474 ;
  assign n3629 = \wb0_cyc_i_pad  & \wb1s_data_i[0]_pad  ;
  assign n3630 = ~n3406 & n3629 ;
  assign n3631 = ~n3628 & ~n3630 ;
  assign n3632 = \u0_wb_rf_dout_reg[10]/P0001  & ~n3474 ;
  assign n3633 = \wb0_cyc_i_pad  & \wb1s_data_i[10]_pad  ;
  assign n3634 = ~n3406 & n3633 ;
  assign n3635 = ~n3632 & ~n3634 ;
  assign n3636 = \u0_wb_rf_dout_reg[11]/P0001  & ~n3474 ;
  assign n3637 = \wb0_cyc_i_pad  & \wb1s_data_i[11]_pad  ;
  assign n3638 = ~n3406 & n3637 ;
  assign n3639 = ~n3636 & ~n3638 ;
  assign n3640 = \u0_wb_rf_dout_reg[12]/P0001  & ~n3474 ;
  assign n3641 = \wb0_cyc_i_pad  & \wb1s_data_i[12]_pad  ;
  assign n3642 = ~n3406 & n3641 ;
  assign n3643 = ~n3640 & ~n3642 ;
  assign n3644 = \u0_wb_rf_dout_reg[13]/P0001  & ~n3474 ;
  assign n3645 = \wb0_cyc_i_pad  & \wb1s_data_i[13]_pad  ;
  assign n3646 = ~n3406 & n3645 ;
  assign n3647 = ~n3644 & ~n3646 ;
  assign n3648 = \u0_wb_rf_dout_reg[14]/P0001  & ~n3474 ;
  assign n3649 = \wb0_cyc_i_pad  & \wb1s_data_i[14]_pad  ;
  assign n3650 = ~n3406 & n3649 ;
  assign n3651 = ~n3648 & ~n3650 ;
  assign n3652 = \u0_wb_rf_dout_reg[15]/P0001  & ~n3474 ;
  assign n3653 = \wb0_cyc_i_pad  & \wb1s_data_i[15]_pad  ;
  assign n3654 = ~n3406 & n3653 ;
  assign n3655 = ~n3652 & ~n3654 ;
  assign n3656 = \u0_wb_rf_dout_reg[16]/P0001  & ~n3474 ;
  assign n3657 = \wb0_cyc_i_pad  & \wb1s_data_i[16]_pad  ;
  assign n3658 = ~n3406 & n3657 ;
  assign n3659 = ~n3656 & ~n3658 ;
  assign n3660 = \u0_wb_rf_dout_reg[17]/P0001  & ~n3474 ;
  assign n3661 = \wb0_cyc_i_pad  & \wb1s_data_i[17]_pad  ;
  assign n3662 = ~n3406 & n3661 ;
  assign n3663 = ~n3660 & ~n3662 ;
  assign n3664 = \u0_wb_rf_dout_reg[18]/P0001  & ~n3474 ;
  assign n3665 = \wb0_cyc_i_pad  & \wb1s_data_i[18]_pad  ;
  assign n3666 = ~n3406 & n3665 ;
  assign n3667 = ~n3664 & ~n3666 ;
  assign n3668 = \u0_wb_rf_dout_reg[19]/P0001  & ~n3474 ;
  assign n3669 = \wb0_cyc_i_pad  & \wb1s_data_i[19]_pad  ;
  assign n3670 = ~n3406 & n3669 ;
  assign n3671 = ~n3668 & ~n3670 ;
  assign n3672 = \u0_wb_rf_dout_reg[1]/P0001  & ~n3474 ;
  assign n3673 = \wb0_cyc_i_pad  & \wb1s_data_i[1]_pad  ;
  assign n3674 = ~n3406 & n3673 ;
  assign n3675 = ~n3672 & ~n3674 ;
  assign n3676 = \u0_wb_rf_dout_reg[20]/P0001  & ~n3474 ;
  assign n3677 = \wb0_cyc_i_pad  & \wb1s_data_i[20]_pad  ;
  assign n3678 = ~n3406 & n3677 ;
  assign n3679 = ~n3676 & ~n3678 ;
  assign n3680 = \u0_wb_rf_dout_reg[21]/P0001  & ~n3474 ;
  assign n3681 = \wb0_cyc_i_pad  & \wb1s_data_i[21]_pad  ;
  assign n3682 = ~n3406 & n3681 ;
  assign n3683 = ~n3680 & ~n3682 ;
  assign n3684 = \u0_wb_rf_dout_reg[22]/P0001  & ~n3474 ;
  assign n3685 = \wb0_cyc_i_pad  & \wb1s_data_i[22]_pad  ;
  assign n3686 = ~n3406 & n3685 ;
  assign n3687 = ~n3684 & ~n3686 ;
  assign n3688 = \u0_wb_rf_dout_reg[23]/P0001  & ~n3474 ;
  assign n3689 = \wb0_cyc_i_pad  & \wb1s_data_i[23]_pad  ;
  assign n3690 = ~n3406 & n3689 ;
  assign n3691 = ~n3688 & ~n3690 ;
  assign n3692 = \u0_wb_rf_dout_reg[24]/P0001  & ~n3474 ;
  assign n3693 = \wb0_cyc_i_pad  & \wb1s_data_i[24]_pad  ;
  assign n3694 = ~n3406 & n3693 ;
  assign n3695 = ~n3692 & ~n3694 ;
  assign n3696 = \u0_wb_rf_dout_reg[25]/P0001  & ~n3474 ;
  assign n3697 = \wb0_cyc_i_pad  & \wb1s_data_i[25]_pad  ;
  assign n3698 = ~n3406 & n3697 ;
  assign n3699 = ~n3696 & ~n3698 ;
  assign n3700 = \u0_wb_rf_dout_reg[26]/P0001  & ~n3474 ;
  assign n3701 = \wb0_cyc_i_pad  & \wb1s_data_i[26]_pad  ;
  assign n3702 = ~n3406 & n3701 ;
  assign n3703 = ~n3700 & ~n3702 ;
  assign n3704 = \u0_wb_rf_dout_reg[27]/P0001  & ~n3474 ;
  assign n3705 = \wb0_cyc_i_pad  & \wb1s_data_i[27]_pad  ;
  assign n3706 = ~n3406 & n3705 ;
  assign n3707 = ~n3704 & ~n3706 ;
  assign n3708 = \u0_wb_rf_dout_reg[28]/P0001  & ~n3474 ;
  assign n3709 = \wb0_cyc_i_pad  & \wb1s_data_i[28]_pad  ;
  assign n3710 = ~n3406 & n3709 ;
  assign n3711 = ~n3708 & ~n3710 ;
  assign n3712 = \u0_wb_rf_dout_reg[29]/P0001  & ~n3474 ;
  assign n3713 = \wb0_cyc_i_pad  & \wb1s_data_i[29]_pad  ;
  assign n3714 = ~n3406 & n3713 ;
  assign n3715 = ~n3712 & ~n3714 ;
  assign n3716 = \u0_wb_rf_dout_reg[2]/P0001  & ~n3474 ;
  assign n3717 = \wb0_cyc_i_pad  & \wb1s_data_i[2]_pad  ;
  assign n3718 = ~n3406 & n3717 ;
  assign n3719 = ~n3716 & ~n3718 ;
  assign n3720 = \u0_wb_rf_dout_reg[30]/P0001  & ~n3474 ;
  assign n3721 = \wb0_cyc_i_pad  & \wb1s_data_i[30]_pad  ;
  assign n3722 = ~n3406 & n3721 ;
  assign n3723 = ~n3720 & ~n3722 ;
  assign n3724 = \u0_wb_rf_dout_reg[31]/P0001  & ~n3474 ;
  assign n3725 = \wb0_cyc_i_pad  & \wb1s_data_i[31]_pad  ;
  assign n3726 = ~n3406 & n3725 ;
  assign n3727 = ~n3724 & ~n3726 ;
  assign n3728 = \u0_wb_rf_dout_reg[3]/P0001  & ~n3474 ;
  assign n3729 = \wb0_cyc_i_pad  & \wb1s_data_i[3]_pad  ;
  assign n3730 = ~n3406 & n3729 ;
  assign n3731 = ~n3728 & ~n3730 ;
  assign n3732 = \u0_wb_rf_dout_reg[4]/P0001  & ~n3474 ;
  assign n3733 = \wb0_cyc_i_pad  & \wb1s_data_i[4]_pad  ;
  assign n3734 = ~n3406 & n3733 ;
  assign n3735 = ~n3732 & ~n3734 ;
  assign n3736 = \u0_wb_rf_dout_reg[5]/P0001  & ~n3474 ;
  assign n3737 = \wb0_cyc_i_pad  & \wb1s_data_i[5]_pad  ;
  assign n3738 = ~n3406 & n3737 ;
  assign n3739 = ~n3736 & ~n3738 ;
  assign n3740 = \u0_wb_rf_dout_reg[6]/P0001  & ~n3474 ;
  assign n3741 = \wb0_cyc_i_pad  & \wb1s_data_i[6]_pad  ;
  assign n3742 = ~n3406 & n3741 ;
  assign n3743 = ~n3740 & ~n3742 ;
  assign n3744 = \u0_wb_rf_dout_reg[7]/P0001  & ~n3474 ;
  assign n3745 = \wb0_cyc_i_pad  & \wb1s_data_i[7]_pad  ;
  assign n3746 = ~n3406 & n3745 ;
  assign n3747 = ~n3744 & ~n3746 ;
  assign n3748 = \u0_wb_rf_dout_reg[8]/P0001  & ~n3474 ;
  assign n3749 = \wb0_cyc_i_pad  & \wb1s_data_i[8]_pad  ;
  assign n3750 = ~n3406 & n3749 ;
  assign n3751 = ~n3748 & ~n3750 ;
  assign n3752 = \u0_wb_rf_dout_reg[9]/P0001  & ~n3474 ;
  assign n3753 = \wb0_cyc_i_pad  & \wb1s_data_i[9]_pad  ;
  assign n3754 = ~n3406 & n3753 ;
  assign n3755 = ~n3752 & ~n3754 ;
  assign n3756 = \wb1_cyc_i_pad  & \wb1m_data_i[0]_pad  ;
  assign n3757 = ~n3399 & n3756 ;
  assign n3758 = \u0_u0_ch_csr_r_reg[2]/NET0131  & \u4_u0_mast_dout_reg[0]/P0001  ;
  assign n3759 = ~\u0_u0_ch_csr_r_reg[2]/NET0131  & \u3_u0_mast_dout_reg[0]/P0001  ;
  assign n3760 = ~n3758 & ~n3759 ;
  assign n3761 = ~n965 & n3760 ;
  assign n3762 = ~n1007 & n3761 ;
  assign n3763 = ~\u2_tsz_cnt_reg[0]/NET0131  & n965 ;
  assign n3764 = ~\u2_tsz_cnt_reg[0]/NET0131  & n1002 ;
  assign n3765 = n1006 & n3764 ;
  assign n3766 = ~n3763 & ~n3765 ;
  assign n3767 = ~n3481 & n3766 ;
  assign n3768 = ~n3762 & n3767 ;
  assign n3769 = ~n3757 & ~n3768 ;
  assign n3770 = \wb1_cyc_i_pad  & \wb1m_data_i[10]_pad  ;
  assign n3771 = ~n3399 & n3770 ;
  assign n3772 = \u0_u0_ch_csr_r_reg[2]/NET0131  & \u4_u0_mast_dout_reg[10]/P0001  ;
  assign n3773 = ~\u0_u0_ch_csr_r_reg[2]/NET0131  & \u3_u0_mast_dout_reg[10]/P0001  ;
  assign n3774 = ~n3772 & ~n3773 ;
  assign n3775 = ~n965 & n3774 ;
  assign n3776 = ~n1007 & n3775 ;
  assign n3777 = ~\u2_tsz_cnt_reg[10]/NET0131  & n965 ;
  assign n3778 = ~\u2_tsz_cnt_reg[10]/NET0131  & n1002 ;
  assign n3779 = n1006 & n3778 ;
  assign n3780 = ~n3777 & ~n3779 ;
  assign n3781 = ~n3481 & n3780 ;
  assign n3782 = ~n3776 & n3781 ;
  assign n3783 = ~n3771 & ~n3782 ;
  assign n3784 = \wb1_cyc_i_pad  & \wb1m_data_i[11]_pad  ;
  assign n3785 = ~n3399 & n3784 ;
  assign n3786 = \u0_u0_ch_csr_r_reg[2]/NET0131  & \u4_u0_mast_dout_reg[11]/P0001  ;
  assign n3787 = ~\u0_u0_ch_csr_r_reg[2]/NET0131  & \u3_u0_mast_dout_reg[11]/P0001  ;
  assign n3788 = ~n3786 & ~n3787 ;
  assign n3789 = ~n965 & n3788 ;
  assign n3790 = ~n1007 & n3789 ;
  assign n3791 = ~\u2_tsz_cnt_reg[11]/NET0131  & n965 ;
  assign n3792 = ~\u2_tsz_cnt_reg[11]/NET0131  & n1002 ;
  assign n3793 = n1006 & n3792 ;
  assign n3794 = ~n3791 & ~n3793 ;
  assign n3795 = ~n3481 & n3794 ;
  assign n3796 = ~n3790 & n3795 ;
  assign n3797 = ~n3785 & ~n3796 ;
  assign n3798 = \wb1_cyc_i_pad  & \wb1m_data_i[12]_pad  ;
  assign n3799 = ~n3399 & n3798 ;
  assign n3800 = \u0_u0_ch_csr_r_reg[2]/NET0131  & \u4_u0_mast_dout_reg[12]/P0001  ;
  assign n3801 = ~\u0_u0_ch_csr_r_reg[2]/NET0131  & \u3_u0_mast_dout_reg[12]/P0001  ;
  assign n3802 = ~n3800 & ~n3801 ;
  assign n3803 = ~n965 & ~n3802 ;
  assign n3804 = ~n3481 & n3803 ;
  assign n3805 = ~n1007 & n3804 ;
  assign n3806 = ~n3799 & ~n3805 ;
  assign n3807 = \wb1_cyc_i_pad  & \wb1m_data_i[13]_pad  ;
  assign n3808 = ~n3399 & n3807 ;
  assign n3809 = \u0_u0_ch_csr_r_reg[2]/NET0131  & \u4_u0_mast_dout_reg[13]/P0001  ;
  assign n3810 = ~\u0_u0_ch_csr_r_reg[2]/NET0131  & \u3_u0_mast_dout_reg[13]/P0001  ;
  assign n3811 = ~n3809 & ~n3810 ;
  assign n3812 = ~n965 & ~n3811 ;
  assign n3813 = ~n3481 & n3812 ;
  assign n3814 = ~n1007 & n3813 ;
  assign n3815 = ~n3808 & ~n3814 ;
  assign n3816 = \wb1_cyc_i_pad  & \wb1m_data_i[14]_pad  ;
  assign n3817 = ~n3399 & n3816 ;
  assign n3818 = \u0_u0_ch_csr_r_reg[2]/NET0131  & \u4_u0_mast_dout_reg[14]/P0001  ;
  assign n3819 = ~\u0_u0_ch_csr_r_reg[2]/NET0131  & \u3_u0_mast_dout_reg[14]/P0001  ;
  assign n3820 = ~n3818 & ~n3819 ;
  assign n3821 = ~n965 & ~n3820 ;
  assign n3822 = ~n3481 & n3821 ;
  assign n3823 = ~n1007 & n3822 ;
  assign n3824 = ~n3817 & ~n3823 ;
  assign n3825 = \wb1_cyc_i_pad  & \wb1m_data_i[15]_pad  ;
  assign n3826 = ~n3399 & n3825 ;
  assign n3827 = \u0_u0_ch_csr_r_reg[2]/NET0131  & \u4_u0_mast_dout_reg[15]/P0001  ;
  assign n3828 = ~\u0_u0_ch_csr_r_reg[2]/NET0131  & \u3_u0_mast_dout_reg[15]/P0001  ;
  assign n3829 = ~n3827 & ~n3828 ;
  assign n3830 = ~n965 & ~n3829 ;
  assign n3831 = ~n3481 & n3830 ;
  assign n3832 = ~n1007 & n3831 ;
  assign n3833 = ~n3826 & ~n3832 ;
  assign n3834 = \wb1_cyc_i_pad  & \wb1m_data_i[16]_pad  ;
  assign n3835 = ~n3399 & n3834 ;
  assign n3836 = \u0_u0_ch_csr_r_reg[2]/NET0131  & \u4_u0_mast_dout_reg[16]/P0001  ;
  assign n3837 = ~\u0_u0_ch_csr_r_reg[2]/NET0131  & \u3_u0_mast_dout_reg[16]/P0001  ;
  assign n3838 = ~n3836 & ~n3837 ;
  assign n3839 = ~n965 & ~n3838 ;
  assign n3840 = ~n3481 & n3839 ;
  assign n3841 = ~n1007 & n3840 ;
  assign n3842 = ~n3835 & ~n3841 ;
  assign n3843 = \wb1_cyc_i_pad  & \wb1m_data_i[17]_pad  ;
  assign n3844 = ~n3399 & n3843 ;
  assign n3845 = \u0_u0_ch_csr_r_reg[2]/NET0131  & \u4_u0_mast_dout_reg[17]/P0001  ;
  assign n3846 = ~\u0_u0_ch_csr_r_reg[2]/NET0131  & \u3_u0_mast_dout_reg[17]/P0001  ;
  assign n3847 = ~n3845 & ~n3846 ;
  assign n3848 = ~n965 & ~n3847 ;
  assign n3849 = ~n3481 & n3848 ;
  assign n3850 = ~n1007 & n3849 ;
  assign n3851 = ~n3844 & ~n3850 ;
  assign n3852 = \wb1_cyc_i_pad  & \wb1m_data_i[18]_pad  ;
  assign n3853 = ~n3399 & n3852 ;
  assign n3854 = \u0_u0_ch_csr_r_reg[2]/NET0131  & \u4_u0_mast_dout_reg[18]/P0001  ;
  assign n3855 = ~\u0_u0_ch_csr_r_reg[2]/NET0131  & \u3_u0_mast_dout_reg[18]/P0001  ;
  assign n3856 = ~n3854 & ~n3855 ;
  assign n3857 = ~n965 & ~n3856 ;
  assign n3858 = ~n3481 & n3857 ;
  assign n3859 = ~n1007 & n3858 ;
  assign n3860 = ~n3853 & ~n3859 ;
  assign n3861 = \wb1_cyc_i_pad  & \wb1m_data_i[19]_pad  ;
  assign n3862 = ~n3399 & n3861 ;
  assign n3863 = \u0_u0_ch_csr_r_reg[2]/NET0131  & \u4_u0_mast_dout_reg[19]/P0001  ;
  assign n3864 = ~\u0_u0_ch_csr_r_reg[2]/NET0131  & \u3_u0_mast_dout_reg[19]/P0001  ;
  assign n3865 = ~n3863 & ~n3864 ;
  assign n3866 = ~n965 & ~n3865 ;
  assign n3867 = ~n3481 & n3866 ;
  assign n3868 = ~n1007 & n3867 ;
  assign n3869 = ~n3862 & ~n3868 ;
  assign n3870 = \wb1_cyc_i_pad  & \wb1m_data_i[1]_pad  ;
  assign n3871 = ~n3399 & n3870 ;
  assign n3872 = \u0_u0_ch_csr_r_reg[2]/NET0131  & \u4_u0_mast_dout_reg[1]/P0001  ;
  assign n3873 = ~\u0_u0_ch_csr_r_reg[2]/NET0131  & \u3_u0_mast_dout_reg[1]/P0001  ;
  assign n3874 = ~n3872 & ~n3873 ;
  assign n3875 = ~n965 & n3874 ;
  assign n3876 = ~n1007 & n3875 ;
  assign n3877 = ~\u2_tsz_cnt_reg[1]/NET0131  & n965 ;
  assign n3878 = ~\u2_tsz_cnt_reg[1]/NET0131  & n1002 ;
  assign n3879 = n1006 & n3878 ;
  assign n3880 = ~n3877 & ~n3879 ;
  assign n3881 = ~n3481 & n3880 ;
  assign n3882 = ~n3876 & n3881 ;
  assign n3883 = ~n3871 & ~n3882 ;
  assign n3884 = \wb1_cyc_i_pad  & \wb1m_data_i[20]_pad  ;
  assign n3885 = ~n3399 & n3884 ;
  assign n3886 = \u0_u0_ch_csr_r_reg[2]/NET0131  & \u4_u0_mast_dout_reg[20]/P0001  ;
  assign n3887 = ~\u0_u0_ch_csr_r_reg[2]/NET0131  & \u3_u0_mast_dout_reg[20]/P0001  ;
  assign n3888 = ~n3886 & ~n3887 ;
  assign n3889 = ~n965 & ~n3888 ;
  assign n3890 = ~n3481 & n3889 ;
  assign n3891 = ~n1007 & n3890 ;
  assign n3892 = ~n3885 & ~n3891 ;
  assign n3893 = \wb1_cyc_i_pad  & \wb1m_data_i[21]_pad  ;
  assign n3894 = ~n3399 & n3893 ;
  assign n3895 = \u0_u0_ch_csr_r_reg[2]/NET0131  & \u4_u0_mast_dout_reg[21]/P0001  ;
  assign n3896 = ~\u0_u0_ch_csr_r_reg[2]/NET0131  & \u3_u0_mast_dout_reg[21]/P0001  ;
  assign n3897 = ~n3895 & ~n3896 ;
  assign n3898 = ~n965 & ~n3897 ;
  assign n3899 = ~n3481 & n3898 ;
  assign n3900 = ~n1007 & n3899 ;
  assign n3901 = ~n3894 & ~n3900 ;
  assign n3902 = \wb1_cyc_i_pad  & \wb1m_data_i[22]_pad  ;
  assign n3903 = ~n3399 & n3902 ;
  assign n3904 = \u0_u0_ch_csr_r_reg[2]/NET0131  & \u4_u0_mast_dout_reg[22]/P0001  ;
  assign n3905 = ~\u0_u0_ch_csr_r_reg[2]/NET0131  & \u3_u0_mast_dout_reg[22]/P0001  ;
  assign n3906 = ~n3904 & ~n3905 ;
  assign n3907 = ~n965 & ~n3906 ;
  assign n3908 = ~n3481 & n3907 ;
  assign n3909 = ~n1007 & n3908 ;
  assign n3910 = ~n3903 & ~n3909 ;
  assign n3911 = \wb1_cyc_i_pad  & \wb1m_data_i[23]_pad  ;
  assign n3912 = ~n3399 & n3911 ;
  assign n3913 = \u0_u0_ch_csr_r_reg[2]/NET0131  & \u4_u0_mast_dout_reg[23]/P0001  ;
  assign n3914 = ~\u0_u0_ch_csr_r_reg[2]/NET0131  & \u3_u0_mast_dout_reg[23]/P0001  ;
  assign n3915 = ~n3913 & ~n3914 ;
  assign n3916 = ~n965 & ~n3915 ;
  assign n3917 = ~n3481 & n3916 ;
  assign n3918 = ~n1007 & n3917 ;
  assign n3919 = ~n3912 & ~n3918 ;
  assign n3920 = \wb1_cyc_i_pad  & \wb1m_data_i[24]_pad  ;
  assign n3921 = ~n3399 & n3920 ;
  assign n3922 = \u0_u0_ch_csr_r_reg[2]/NET0131  & \u4_u0_mast_dout_reg[24]/P0001  ;
  assign n3923 = ~\u0_u0_ch_csr_r_reg[2]/NET0131  & \u3_u0_mast_dout_reg[24]/P0001  ;
  assign n3924 = ~n3922 & ~n3923 ;
  assign n3925 = ~n965 & ~n3924 ;
  assign n3926 = ~n3481 & n3925 ;
  assign n3927 = ~n1007 & n3926 ;
  assign n3928 = ~n3921 & ~n3927 ;
  assign n3929 = \wb1_cyc_i_pad  & \wb1m_data_i[25]_pad  ;
  assign n3930 = ~n3399 & n3929 ;
  assign n3931 = \u0_u0_ch_csr_r_reg[2]/NET0131  & \u4_u0_mast_dout_reg[25]/P0001  ;
  assign n3932 = ~\u0_u0_ch_csr_r_reg[2]/NET0131  & \u3_u0_mast_dout_reg[25]/P0001  ;
  assign n3933 = ~n3931 & ~n3932 ;
  assign n3934 = ~n965 & ~n3933 ;
  assign n3935 = ~n3481 & n3934 ;
  assign n3936 = ~n1007 & n3935 ;
  assign n3937 = ~n3930 & ~n3936 ;
  assign n3938 = \wb1_cyc_i_pad  & \wb1m_data_i[26]_pad  ;
  assign n3939 = ~n3399 & n3938 ;
  assign n3940 = \u0_u0_ch_csr_r_reg[2]/NET0131  & \u4_u0_mast_dout_reg[26]/P0001  ;
  assign n3941 = ~\u0_u0_ch_csr_r_reg[2]/NET0131  & \u3_u0_mast_dout_reg[26]/P0001  ;
  assign n3942 = ~n3940 & ~n3941 ;
  assign n3943 = ~n965 & ~n3942 ;
  assign n3944 = ~n3481 & n3943 ;
  assign n3945 = ~n1007 & n3944 ;
  assign n3946 = ~n3939 & ~n3945 ;
  assign n3947 = \wb1_cyc_i_pad  & \wb1m_data_i[27]_pad  ;
  assign n3948 = ~n3399 & n3947 ;
  assign n3949 = \u0_u0_ch_csr_r_reg[2]/NET0131  & \u4_u0_mast_dout_reg[27]/P0001  ;
  assign n3950 = ~\u0_u0_ch_csr_r_reg[2]/NET0131  & \u3_u0_mast_dout_reg[27]/P0001  ;
  assign n3951 = ~n3949 & ~n3950 ;
  assign n3952 = ~n965 & ~n3951 ;
  assign n3953 = ~n3481 & n3952 ;
  assign n3954 = ~n1007 & n3953 ;
  assign n3955 = ~n3948 & ~n3954 ;
  assign n3956 = \wb1_cyc_i_pad  & \wb1m_data_i[28]_pad  ;
  assign n3957 = ~n3399 & n3956 ;
  assign n3958 = \u0_u0_ch_csr_r_reg[2]/NET0131  & \u4_u0_mast_dout_reg[28]/P0001  ;
  assign n3959 = ~\u0_u0_ch_csr_r_reg[2]/NET0131  & \u3_u0_mast_dout_reg[28]/P0001  ;
  assign n3960 = ~n3958 & ~n3959 ;
  assign n3961 = ~n965 & ~n3960 ;
  assign n3962 = ~n3481 & n3961 ;
  assign n3963 = ~n1007 & n3962 ;
  assign n3964 = ~n3957 & ~n3963 ;
  assign n3965 = \wb1_cyc_i_pad  & \wb1m_data_i[29]_pad  ;
  assign n3966 = ~n3399 & n3965 ;
  assign n3967 = \u0_u0_ch_csr_r_reg[2]/NET0131  & \u4_u0_mast_dout_reg[29]/P0001  ;
  assign n3968 = ~\u0_u0_ch_csr_r_reg[2]/NET0131  & \u3_u0_mast_dout_reg[29]/P0001  ;
  assign n3969 = ~n3967 & ~n3968 ;
  assign n3970 = ~n965 & ~n3969 ;
  assign n3971 = ~n3481 & n3970 ;
  assign n3972 = ~n1007 & n3971 ;
  assign n3973 = ~n3966 & ~n3972 ;
  assign n3974 = \wb1_cyc_i_pad  & \wb1m_data_i[2]_pad  ;
  assign n3975 = ~n3399 & n3974 ;
  assign n3976 = \u0_u0_ch_csr_r_reg[2]/NET0131  & \u4_u0_mast_dout_reg[2]/P0001  ;
  assign n3977 = ~\u0_u0_ch_csr_r_reg[2]/NET0131  & \u3_u0_mast_dout_reg[2]/P0001  ;
  assign n3978 = ~n3976 & ~n3977 ;
  assign n3979 = ~n965 & n3978 ;
  assign n3980 = ~n1007 & n3979 ;
  assign n3981 = ~\u2_tsz_cnt_reg[2]/NET0131  & n965 ;
  assign n3982 = ~\u2_tsz_cnt_reg[2]/NET0131  & n1002 ;
  assign n3983 = n1006 & n3982 ;
  assign n3984 = ~n3981 & ~n3983 ;
  assign n3985 = ~n3481 & n3984 ;
  assign n3986 = ~n3980 & n3985 ;
  assign n3987 = ~n3975 & ~n3986 ;
  assign n3988 = \wb1_cyc_i_pad  & \wb1m_data_i[30]_pad  ;
  assign n3989 = ~n3399 & n3988 ;
  assign n3990 = \u0_u0_ch_csr_r_reg[2]/NET0131  & \u4_u0_mast_dout_reg[30]/P0001  ;
  assign n3991 = ~\u0_u0_ch_csr_r_reg[2]/NET0131  & \u3_u0_mast_dout_reg[30]/P0001  ;
  assign n3992 = ~n3990 & ~n3991 ;
  assign n3993 = ~n965 & ~n3992 ;
  assign n3994 = ~n3481 & n3993 ;
  assign n3995 = ~n1007 & n3994 ;
  assign n3996 = ~n3989 & ~n3995 ;
  assign n3997 = \wb1_cyc_i_pad  & \wb1m_data_i[31]_pad  ;
  assign n3998 = ~n3399 & n3997 ;
  assign n3999 = \u0_u0_ch_csr_r_reg[2]/NET0131  & \u4_u0_mast_dout_reg[31]/P0001  ;
  assign n4000 = ~\u0_u0_ch_csr_r_reg[2]/NET0131  & \u3_u0_mast_dout_reg[31]/P0001  ;
  assign n4001 = ~n3999 & ~n4000 ;
  assign n4002 = ~n965 & ~n4001 ;
  assign n4003 = ~n3481 & n4002 ;
  assign n4004 = ~n1007 & n4003 ;
  assign n4005 = ~n3998 & ~n4004 ;
  assign n4006 = \wb1_cyc_i_pad  & \wb1m_data_i[3]_pad  ;
  assign n4007 = ~n3399 & n4006 ;
  assign n4008 = \u0_u0_ch_csr_r_reg[2]/NET0131  & \u4_u0_mast_dout_reg[3]/P0001  ;
  assign n4009 = ~\u0_u0_ch_csr_r_reg[2]/NET0131  & \u3_u0_mast_dout_reg[3]/P0001  ;
  assign n4010 = ~n4008 & ~n4009 ;
  assign n4011 = ~n965 & n4010 ;
  assign n4012 = ~n1007 & n4011 ;
  assign n4013 = ~\u2_tsz_cnt_reg[3]/NET0131  & n965 ;
  assign n4014 = ~\u2_tsz_cnt_reg[3]/NET0131  & n1002 ;
  assign n4015 = n1006 & n4014 ;
  assign n4016 = ~n4013 & ~n4015 ;
  assign n4017 = ~n3481 & n4016 ;
  assign n4018 = ~n4012 & n4017 ;
  assign n4019 = ~n4007 & ~n4018 ;
  assign n4020 = \wb1_cyc_i_pad  & \wb1m_data_i[4]_pad  ;
  assign n4021 = ~n3399 & n4020 ;
  assign n4022 = \u0_u0_ch_csr_r_reg[2]/NET0131  & \u4_u0_mast_dout_reg[4]/P0001  ;
  assign n4023 = ~\u0_u0_ch_csr_r_reg[2]/NET0131  & \u3_u0_mast_dout_reg[4]/P0001  ;
  assign n4024 = ~n4022 & ~n4023 ;
  assign n4025 = ~n965 & n4024 ;
  assign n4026 = ~n1007 & n4025 ;
  assign n4027 = ~\u2_tsz_cnt_reg[4]/NET0131  & n965 ;
  assign n4028 = ~\u2_tsz_cnt_reg[4]/NET0131  & n1002 ;
  assign n4029 = n1006 & n4028 ;
  assign n4030 = ~n4027 & ~n4029 ;
  assign n4031 = ~n3481 & n4030 ;
  assign n4032 = ~n4026 & n4031 ;
  assign n4033 = ~n4021 & ~n4032 ;
  assign n4034 = \wb1_cyc_i_pad  & \wb1m_data_i[5]_pad  ;
  assign n4035 = ~n3399 & n4034 ;
  assign n4036 = \u0_u0_ch_csr_r_reg[2]/NET0131  & \u4_u0_mast_dout_reg[5]/P0001  ;
  assign n4037 = ~\u0_u0_ch_csr_r_reg[2]/NET0131  & \u3_u0_mast_dout_reg[5]/P0001  ;
  assign n4038 = ~n4036 & ~n4037 ;
  assign n4039 = ~n965 & n4038 ;
  assign n4040 = ~n1007 & n4039 ;
  assign n4041 = ~\u2_tsz_cnt_reg[5]/NET0131  & n965 ;
  assign n4042 = ~\u2_tsz_cnt_reg[5]/NET0131  & n1002 ;
  assign n4043 = n1006 & n4042 ;
  assign n4044 = ~n4041 & ~n4043 ;
  assign n4045 = ~n3481 & n4044 ;
  assign n4046 = ~n4040 & n4045 ;
  assign n4047 = ~n4035 & ~n4046 ;
  assign n4048 = \wb1_cyc_i_pad  & \wb1m_data_i[6]_pad  ;
  assign n4049 = ~n3399 & n4048 ;
  assign n4050 = \u0_u0_ch_csr_r_reg[2]/NET0131  & \u4_u0_mast_dout_reg[6]/P0001  ;
  assign n4051 = ~\u0_u0_ch_csr_r_reg[2]/NET0131  & \u3_u0_mast_dout_reg[6]/P0001  ;
  assign n4052 = ~n4050 & ~n4051 ;
  assign n4053 = ~n965 & n4052 ;
  assign n4054 = ~n1007 & n4053 ;
  assign n4055 = ~\u2_tsz_cnt_reg[6]/NET0131  & n965 ;
  assign n4056 = ~\u2_tsz_cnt_reg[6]/NET0131  & n1002 ;
  assign n4057 = n1006 & n4056 ;
  assign n4058 = ~n4055 & ~n4057 ;
  assign n4059 = ~n3481 & n4058 ;
  assign n4060 = ~n4054 & n4059 ;
  assign n4061 = ~n4049 & ~n4060 ;
  assign n4062 = \wb1_cyc_i_pad  & \wb1m_data_i[7]_pad  ;
  assign n4063 = ~n3399 & n4062 ;
  assign n4064 = \u0_u0_ch_csr_r_reg[2]/NET0131  & \u4_u0_mast_dout_reg[7]/P0001  ;
  assign n4065 = ~\u0_u0_ch_csr_r_reg[2]/NET0131  & \u3_u0_mast_dout_reg[7]/P0001  ;
  assign n4066 = ~n4064 & ~n4065 ;
  assign n4067 = ~n965 & n4066 ;
  assign n4068 = ~n1007 & n4067 ;
  assign n4069 = ~\u2_tsz_cnt_reg[7]/NET0131  & n965 ;
  assign n4070 = ~\u2_tsz_cnt_reg[7]/NET0131  & n1002 ;
  assign n4071 = n1006 & n4070 ;
  assign n4072 = ~n4069 & ~n4071 ;
  assign n4073 = ~n3481 & n4072 ;
  assign n4074 = ~n4068 & n4073 ;
  assign n4075 = ~n4063 & ~n4074 ;
  assign n4076 = \wb1_cyc_i_pad  & \wb1m_data_i[8]_pad  ;
  assign n4077 = ~n3399 & n4076 ;
  assign n4078 = \u0_u0_ch_csr_r_reg[2]/NET0131  & \u4_u0_mast_dout_reg[8]/P0001  ;
  assign n4079 = ~\u0_u0_ch_csr_r_reg[2]/NET0131  & \u3_u0_mast_dout_reg[8]/P0001  ;
  assign n4080 = ~n4078 & ~n4079 ;
  assign n4081 = ~n965 & n4080 ;
  assign n4082 = ~n1007 & n4081 ;
  assign n4083 = ~\u2_tsz_cnt_reg[8]/NET0131  & n965 ;
  assign n4084 = ~\u2_tsz_cnt_reg[8]/NET0131  & n1002 ;
  assign n4085 = n1006 & n4084 ;
  assign n4086 = ~n4083 & ~n4085 ;
  assign n4087 = ~n3481 & n4086 ;
  assign n4088 = ~n4082 & n4087 ;
  assign n4089 = ~n4077 & ~n4088 ;
  assign n4090 = \wb1_cyc_i_pad  & \wb1m_data_i[9]_pad  ;
  assign n4091 = ~n3399 & n4090 ;
  assign n4092 = \u0_u0_ch_csr_r_reg[2]/NET0131  & \u4_u0_mast_dout_reg[9]/P0001  ;
  assign n4093 = ~\u0_u0_ch_csr_r_reg[2]/NET0131  & \u3_u0_mast_dout_reg[9]/P0001  ;
  assign n4094 = ~n4092 & ~n4093 ;
  assign n4095 = ~n965 & n4094 ;
  assign n4096 = ~n1007 & n4095 ;
  assign n4097 = ~\u2_tsz_cnt_reg[9]/NET0131  & n965 ;
  assign n4098 = ~\u2_tsz_cnt_reg[9]/NET0131  & n1002 ;
  assign n4099 = n1006 & n4098 ;
  assign n4100 = ~n4097 & ~n4099 ;
  assign n4101 = ~n3481 & n4100 ;
  assign n4102 = ~n4096 & n4101 ;
  assign n4103 = ~n4091 & ~n4102 ;
  assign n4104 = \u4_u1_rf_ack_reg/P0001  & ~n3481 ;
  assign n4105 = \wb0_ack_i_pad  & \wb1_cyc_i_pad  ;
  assign n4106 = ~n3399 & n4105 ;
  assign n4107 = ~n4104 & ~n4106 ;
  assign n4108 = \wb0_addr_i[0]_pad  & \wb0_cyc_i_pad  ;
  assign n4109 = ~n3406 & n4108 ;
  assign n4110 = \u2_mast1_adr_reg[10]/P0001  & ~n3474 ;
  assign n4111 = \wb0_addr_i[10]_pad  & \wb0_cyc_i_pad  ;
  assign n4112 = ~n3406 & n4111 ;
  assign n4113 = ~n4110 & ~n4112 ;
  assign n4114 = \u2_mast1_adr_reg[11]/P0001  & ~n3474 ;
  assign n4115 = \wb0_addr_i[11]_pad  & \wb0_cyc_i_pad  ;
  assign n4116 = ~n3406 & n4115 ;
  assign n4117 = ~n4114 & ~n4116 ;
  assign n4118 = \u2_mast1_adr_reg[12]/P0001  & ~n3474 ;
  assign n4119 = \wb0_addr_i[12]_pad  & \wb0_cyc_i_pad  ;
  assign n4120 = ~n3406 & n4119 ;
  assign n4121 = ~n4118 & ~n4120 ;
  assign n4122 = \u2_mast1_adr_reg[13]/P0001  & ~n3474 ;
  assign n4123 = \wb0_addr_i[13]_pad  & \wb0_cyc_i_pad  ;
  assign n4124 = ~n3406 & n4123 ;
  assign n4125 = ~n4122 & ~n4124 ;
  assign n4126 = \u2_mast1_adr_reg[14]/P0001  & ~n3474 ;
  assign n4127 = \wb0_addr_i[14]_pad  & \wb0_cyc_i_pad  ;
  assign n4128 = ~n3406 & n4127 ;
  assign n4129 = ~n4126 & ~n4128 ;
  assign n4130 = \u2_mast1_adr_reg[15]/P0001  & ~n3474 ;
  assign n4131 = \wb0_addr_i[15]_pad  & \wb0_cyc_i_pad  ;
  assign n4132 = ~n3406 & n4131 ;
  assign n4133 = ~n4130 & ~n4132 ;
  assign n4134 = \u2_mast1_adr_reg[16]/P0001  & ~n3474 ;
  assign n4135 = \wb0_addr_i[16]_pad  & \wb0_cyc_i_pad  ;
  assign n4136 = ~n3406 & n4135 ;
  assign n4137 = ~n4134 & ~n4136 ;
  assign n4138 = \u2_mast1_adr_reg[17]/P0001  & ~n3474 ;
  assign n4139 = \wb0_addr_i[17]_pad  & \wb0_cyc_i_pad  ;
  assign n4140 = ~n3406 & n4139 ;
  assign n4141 = ~n4138 & ~n4140 ;
  assign n4142 = \u2_mast1_adr_reg[18]/P0001  & ~n3474 ;
  assign n4143 = \wb0_addr_i[18]_pad  & \wb0_cyc_i_pad  ;
  assign n4144 = ~n3406 & n4143 ;
  assign n4145 = ~n4142 & ~n4144 ;
  assign n4146 = \u2_mast1_adr_reg[19]/P0001  & ~n3474 ;
  assign n4147 = \wb0_addr_i[19]_pad  & \wb0_cyc_i_pad  ;
  assign n4148 = ~n3406 & n4147 ;
  assign n4149 = ~n4146 & ~n4148 ;
  assign n4150 = \wb0_addr_i[1]_pad  & \wb0_cyc_i_pad  ;
  assign n4151 = ~n3406 & n4150 ;
  assign n4152 = \u2_mast1_adr_reg[20]/P0001  & ~n3474 ;
  assign n4153 = \wb0_addr_i[20]_pad  & \wb0_cyc_i_pad  ;
  assign n4154 = ~n3406 & n4153 ;
  assign n4155 = ~n4152 & ~n4154 ;
  assign n4156 = \u2_mast1_adr_reg[21]/P0001  & ~n3474 ;
  assign n4157 = \wb0_addr_i[21]_pad  & \wb0_cyc_i_pad  ;
  assign n4158 = ~n3406 & n4157 ;
  assign n4159 = ~n4156 & ~n4158 ;
  assign n4160 = \u2_mast1_adr_reg[22]/P0001  & ~n3474 ;
  assign n4161 = \wb0_addr_i[22]_pad  & \wb0_cyc_i_pad  ;
  assign n4162 = ~n3406 & n4161 ;
  assign n4163 = ~n4160 & ~n4162 ;
  assign n4164 = \u2_mast1_adr_reg[23]/P0001  & ~n3474 ;
  assign n4165 = \wb0_addr_i[23]_pad  & \wb0_cyc_i_pad  ;
  assign n4166 = ~n3406 & n4165 ;
  assign n4167 = ~n4164 & ~n4166 ;
  assign n4168 = \u2_mast1_adr_reg[24]/P0001  & ~n3474 ;
  assign n4169 = \wb0_addr_i[24]_pad  & \wb0_cyc_i_pad  ;
  assign n4170 = ~n3406 & n4169 ;
  assign n4171 = ~n4168 & ~n4170 ;
  assign n4172 = \u2_mast1_adr_reg[25]/P0001  & ~n3474 ;
  assign n4173 = \wb0_addr_i[25]_pad  & \wb0_cyc_i_pad  ;
  assign n4174 = ~n3406 & n4173 ;
  assign n4175 = ~n4172 & ~n4174 ;
  assign n4176 = \u2_mast1_adr_reg[26]/P0001  & ~n3474 ;
  assign n4177 = \wb0_addr_i[26]_pad  & \wb0_cyc_i_pad  ;
  assign n4178 = ~n3406 & n4177 ;
  assign n4179 = ~n4176 & ~n4178 ;
  assign n4180 = \u2_mast1_adr_reg[27]/P0001  & ~n3474 ;
  assign n4181 = \wb0_addr_i[27]_pad  & \wb0_cyc_i_pad  ;
  assign n4182 = ~n3406 & n4181 ;
  assign n4183 = ~n4180 & ~n4182 ;
  assign n4184 = \wb0_addr_i[28]_pad  & \wb0_cyc_i_pad  ;
  assign n4185 = ~\u2_mast1_adr_reg[28]/P0001  & ~n4184 ;
  assign n4186 = \wb0_cyc_i_pad  & ~n4184 ;
  assign n4187 = ~n3406 & n4186 ;
  assign n4188 = ~n4185 & ~n4187 ;
  assign n4189 = \wb0_addr_i[29]_pad  & \wb0_cyc_i_pad  ;
  assign n4190 = ~\u2_mast1_adr_reg[29]/P0001  & ~n4189 ;
  assign n4191 = \wb0_cyc_i_pad  & ~n4189 ;
  assign n4192 = ~n3406 & n4191 ;
  assign n4193 = ~n4190 & ~n4192 ;
  assign n4194 = \u2_mast1_adr_reg[2]/P0001  & ~n3474 ;
  assign n4195 = \wb0_addr_i[2]_pad  & \wb0_cyc_i_pad  ;
  assign n4196 = ~n3406 & n4195 ;
  assign n4197 = ~n4194 & ~n4196 ;
  assign n4198 = \wb0_addr_i[30]_pad  & \wb0_cyc_i_pad  ;
  assign n4199 = ~\u2_mast1_adr_reg[30]/P0001  & ~n4198 ;
  assign n4200 = \wb0_cyc_i_pad  & ~n4198 ;
  assign n4201 = ~n3406 & n4200 ;
  assign n4202 = ~n4199 & ~n4201 ;
  assign n4203 = \wb0_addr_i[31]_pad  & \wb0_cyc_i_pad  ;
  assign n4204 = ~\u2_mast1_adr_reg[31]/P0001  & ~n4203 ;
  assign n4205 = \wb0_cyc_i_pad  & ~n4203 ;
  assign n4206 = ~n3406 & n4205 ;
  assign n4207 = ~n4204 & ~n4206 ;
  assign n4208 = \u2_mast1_adr_reg[3]/P0001  & ~n3474 ;
  assign n4209 = \wb0_addr_i[3]_pad  & \wb0_cyc_i_pad  ;
  assign n4210 = ~n3406 & n4209 ;
  assign n4211 = ~n4208 & ~n4210 ;
  assign n4212 = \u2_mast1_adr_reg[4]/P0001  & ~n3474 ;
  assign n4213 = \wb0_addr_i[4]_pad  & \wb0_cyc_i_pad  ;
  assign n4214 = ~n3406 & n4213 ;
  assign n4215 = ~n4212 & ~n4214 ;
  assign n4216 = \u2_mast1_adr_reg[5]/P0001  & ~n3474 ;
  assign n4217 = \wb0_addr_i[5]_pad  & \wb0_cyc_i_pad  ;
  assign n4218 = ~n3406 & n4217 ;
  assign n4219 = ~n4216 & ~n4218 ;
  assign n4220 = \u2_mast1_adr_reg[6]/P0001  & ~n3474 ;
  assign n4221 = \wb0_addr_i[6]_pad  & \wb0_cyc_i_pad  ;
  assign n4222 = ~n3406 & n4221 ;
  assign n4223 = ~n4220 & ~n4222 ;
  assign n4224 = \u2_mast1_adr_reg[7]/P0001  & ~n3474 ;
  assign n4225 = \wb0_addr_i[7]_pad  & \wb0_cyc_i_pad  ;
  assign n4226 = ~n3406 & n4225 ;
  assign n4227 = ~n4224 & ~n4226 ;
  assign n4228 = \u2_mast1_adr_reg[8]/P0001  & ~n3474 ;
  assign n4229 = \wb0_addr_i[8]_pad  & \wb0_cyc_i_pad  ;
  assign n4230 = ~n3406 & n4229 ;
  assign n4231 = ~n4228 & ~n4230 ;
  assign n4232 = \u2_mast1_adr_reg[9]/P0001  & ~n3474 ;
  assign n4233 = \wb0_addr_i[9]_pad  & \wb0_cyc_i_pad  ;
  assign n4234 = ~n3406 & n4233 ;
  assign n4235 = ~n4232 & ~n4234 ;
  assign n4236 = ~\u4_u0_mast_cyc_reg/P0001  & ~n3474 ;
  assign n4237 = \wb0_err_i_pad  & \wb1_cyc_i_pad  ;
  assign n4238 = ~n3399 & n4237 ;
  assign n4239 = \wb0_rty_i_pad  & \wb1_cyc_i_pad  ;
  assign n4240 = ~n3399 & n4239 ;
  assign n4241 = \wb0_cyc_i_pad  & ~\wb0_sel_i[0]_pad  ;
  assign n4242 = ~n3406 & n4241 ;
  assign n4243 = \wb0_cyc_i_pad  & ~\wb0_sel_i[1]_pad  ;
  assign n4244 = ~n3406 & n4243 ;
  assign n4245 = \wb0_cyc_i_pad  & ~\wb0_sel_i[2]_pad  ;
  assign n4246 = ~n3406 & n4245 ;
  assign n4247 = \wb0_cyc_i_pad  & ~\wb0_sel_i[3]_pad  ;
  assign n4248 = ~n3406 & n4247 ;
  assign n4249 = \u4_u0_mast_stb_reg/P0001  & ~n3474 ;
  assign n4250 = \wb0_cyc_i_pad  & \wb0_stb_i_pad  ;
  assign n4251 = ~n3406 & n4250 ;
  assign n4252 = ~n4249 & ~n4251 ;
  assign n4253 = \u4_u0_mast_we_r_reg/P0001  & ~n3474 ;
  assign n4254 = \wb0_cyc_i_pad  & \wb0_we_i_pad  ;
  assign n4255 = ~n3406 & n4254 ;
  assign n4256 = ~n4253 & ~n4255 ;
  assign n4257 = \wb0s_data_i[0]_pad  & \wb1_cyc_i_pad  ;
  assign n4258 = ~n3399 & n4257 ;
  assign n4259 = \wb0s_data_i[10]_pad  & \wb1_cyc_i_pad  ;
  assign n4260 = ~n3399 & n4259 ;
  assign n4261 = \wb0s_data_i[11]_pad  & \wb1_cyc_i_pad  ;
  assign n4262 = ~n3399 & n4261 ;
  assign n4263 = \wb0s_data_i[12]_pad  & \wb1_cyc_i_pad  ;
  assign n4264 = ~n3399 & n4263 ;
  assign n4265 = \wb0s_data_i[13]_pad  & \wb1_cyc_i_pad  ;
  assign n4266 = ~n3399 & n4265 ;
  assign n4267 = \wb0s_data_i[14]_pad  & \wb1_cyc_i_pad  ;
  assign n4268 = ~n3399 & n4267 ;
  assign n4269 = \wb0s_data_i[15]_pad  & \wb1_cyc_i_pad  ;
  assign n4270 = ~n3399 & n4269 ;
  assign n4271 = \wb0s_data_i[16]_pad  & \wb1_cyc_i_pad  ;
  assign n4272 = ~n3399 & n4271 ;
  assign n4273 = \wb0s_data_i[17]_pad  & \wb1_cyc_i_pad  ;
  assign n4274 = ~n3399 & n4273 ;
  assign n4275 = \wb0s_data_i[18]_pad  & \wb1_cyc_i_pad  ;
  assign n4276 = ~n3399 & n4275 ;
  assign n4277 = \wb0s_data_i[19]_pad  & \wb1_cyc_i_pad  ;
  assign n4278 = ~n3399 & n4277 ;
  assign n4279 = \wb0s_data_i[1]_pad  & \wb1_cyc_i_pad  ;
  assign n4280 = ~n3399 & n4279 ;
  assign n4281 = \wb0s_data_i[20]_pad  & \wb1_cyc_i_pad  ;
  assign n4282 = ~n3399 & n4281 ;
  assign n4283 = \wb0s_data_i[21]_pad  & \wb1_cyc_i_pad  ;
  assign n4284 = ~n3399 & n4283 ;
  assign n4285 = \wb0s_data_i[22]_pad  & \wb1_cyc_i_pad  ;
  assign n4286 = ~n3399 & n4285 ;
  assign n4287 = \wb0s_data_i[23]_pad  & \wb1_cyc_i_pad  ;
  assign n4288 = ~n3399 & n4287 ;
  assign n4289 = \wb0s_data_i[24]_pad  & \wb1_cyc_i_pad  ;
  assign n4290 = ~n3399 & n4289 ;
  assign n4291 = \wb0s_data_i[25]_pad  & \wb1_cyc_i_pad  ;
  assign n4292 = ~n3399 & n4291 ;
  assign n4293 = \wb0s_data_i[26]_pad  & \wb1_cyc_i_pad  ;
  assign n4294 = ~n3399 & n4293 ;
  assign n4295 = \wb0s_data_i[27]_pad  & \wb1_cyc_i_pad  ;
  assign n4296 = ~n3399 & n4295 ;
  assign n4297 = \wb0s_data_i[28]_pad  & \wb1_cyc_i_pad  ;
  assign n4298 = ~n3399 & n4297 ;
  assign n4299 = \wb0s_data_i[29]_pad  & \wb1_cyc_i_pad  ;
  assign n4300 = ~n3399 & n4299 ;
  assign n4301 = \wb0s_data_i[2]_pad  & \wb1_cyc_i_pad  ;
  assign n4302 = ~n3399 & n4301 ;
  assign n4303 = \wb0s_data_i[30]_pad  & \wb1_cyc_i_pad  ;
  assign n4304 = ~n3399 & n4303 ;
  assign n4305 = \wb0s_data_i[31]_pad  & \wb1_cyc_i_pad  ;
  assign n4306 = ~n3399 & n4305 ;
  assign n4307 = \wb0s_data_i[3]_pad  & \wb1_cyc_i_pad  ;
  assign n4308 = ~n3399 & n4307 ;
  assign n4309 = \wb0s_data_i[4]_pad  & \wb1_cyc_i_pad  ;
  assign n4310 = ~n3399 & n4309 ;
  assign n4311 = \wb0s_data_i[5]_pad  & \wb1_cyc_i_pad  ;
  assign n4312 = ~n3399 & n4311 ;
  assign n4313 = \wb0s_data_i[6]_pad  & \wb1_cyc_i_pad  ;
  assign n4314 = ~n3399 & n4313 ;
  assign n4315 = \wb0s_data_i[7]_pad  & \wb1_cyc_i_pad  ;
  assign n4316 = ~n3399 & n4315 ;
  assign n4317 = \wb0s_data_i[8]_pad  & \wb1_cyc_i_pad  ;
  assign n4318 = ~n3399 & n4317 ;
  assign n4319 = \wb0s_data_i[9]_pad  & \wb1_cyc_i_pad  ;
  assign n4320 = ~n3399 & n4319 ;
  assign n4321 = ~n3474 & n3760 ;
  assign n4322 = \wb0_cyc_i_pad  & ~\wb0m_data_i[0]_pad  ;
  assign n4323 = ~n3406 & n4322 ;
  assign n4324 = ~n4321 & ~n4323 ;
  assign n4325 = ~n3474 & n3774 ;
  assign n4326 = \wb0_cyc_i_pad  & ~\wb0m_data_i[10]_pad  ;
  assign n4327 = ~n3406 & n4326 ;
  assign n4328 = ~n4325 & ~n4327 ;
  assign n4329 = ~n3474 & n3788 ;
  assign n4330 = \wb0_cyc_i_pad  & ~\wb0m_data_i[11]_pad  ;
  assign n4331 = ~n3406 & n4330 ;
  assign n4332 = ~n4329 & ~n4331 ;
  assign n4333 = ~n3474 & n3802 ;
  assign n4334 = \wb0_cyc_i_pad  & ~\wb0m_data_i[12]_pad  ;
  assign n4335 = ~n3406 & n4334 ;
  assign n4336 = ~n4333 & ~n4335 ;
  assign n4337 = ~n3474 & n3811 ;
  assign n4338 = \wb0_cyc_i_pad  & ~\wb0m_data_i[13]_pad  ;
  assign n4339 = ~n3406 & n4338 ;
  assign n4340 = ~n4337 & ~n4339 ;
  assign n4341 = ~n3474 & n3820 ;
  assign n4342 = \wb0_cyc_i_pad  & ~\wb0m_data_i[14]_pad  ;
  assign n4343 = ~n3406 & n4342 ;
  assign n4344 = ~n4341 & ~n4343 ;
  assign n4345 = ~n3474 & n3829 ;
  assign n4346 = \wb0_cyc_i_pad  & ~\wb0m_data_i[15]_pad  ;
  assign n4347 = ~n3406 & n4346 ;
  assign n4348 = ~n4345 & ~n4347 ;
  assign n4349 = ~n3474 & n3838 ;
  assign n4350 = \wb0_cyc_i_pad  & ~\wb0m_data_i[16]_pad  ;
  assign n4351 = ~n3406 & n4350 ;
  assign n4352 = ~n4349 & ~n4351 ;
  assign n4353 = ~n3474 & n3847 ;
  assign n4354 = \wb0_cyc_i_pad  & ~\wb0m_data_i[17]_pad  ;
  assign n4355 = ~n3406 & n4354 ;
  assign n4356 = ~n4353 & ~n4355 ;
  assign n4357 = ~n3474 & n3856 ;
  assign n4358 = \wb0_cyc_i_pad  & ~\wb0m_data_i[18]_pad  ;
  assign n4359 = ~n3406 & n4358 ;
  assign n4360 = ~n4357 & ~n4359 ;
  assign n4361 = ~n3474 & n3865 ;
  assign n4362 = \wb0_cyc_i_pad  & ~\wb0m_data_i[19]_pad  ;
  assign n4363 = ~n3406 & n4362 ;
  assign n4364 = ~n4361 & ~n4363 ;
  assign n4365 = ~n3474 & n3874 ;
  assign n4366 = \wb0_cyc_i_pad  & ~\wb0m_data_i[1]_pad  ;
  assign n4367 = ~n3406 & n4366 ;
  assign n4368 = ~n4365 & ~n4367 ;
  assign n4369 = ~n3474 & n3888 ;
  assign n4370 = \wb0_cyc_i_pad  & ~\wb0m_data_i[20]_pad  ;
  assign n4371 = ~n3406 & n4370 ;
  assign n4372 = ~n4369 & ~n4371 ;
  assign n4373 = ~n3474 & n3897 ;
  assign n4374 = \wb0_cyc_i_pad  & ~\wb0m_data_i[21]_pad  ;
  assign n4375 = ~n3406 & n4374 ;
  assign n4376 = ~n4373 & ~n4375 ;
  assign n4377 = ~n3474 & n3906 ;
  assign n4378 = \wb0_cyc_i_pad  & ~\wb0m_data_i[22]_pad  ;
  assign n4379 = ~n3406 & n4378 ;
  assign n4380 = ~n4377 & ~n4379 ;
  assign n4381 = ~n3474 & n3915 ;
  assign n4382 = \wb0_cyc_i_pad  & ~\wb0m_data_i[23]_pad  ;
  assign n4383 = ~n3406 & n4382 ;
  assign n4384 = ~n4381 & ~n4383 ;
  assign n4385 = ~n3474 & n3924 ;
  assign n4386 = \wb0_cyc_i_pad  & ~\wb0m_data_i[24]_pad  ;
  assign n4387 = ~n3406 & n4386 ;
  assign n4388 = ~n4385 & ~n4387 ;
  assign n4389 = ~n3474 & n3933 ;
  assign n4390 = \wb0_cyc_i_pad  & ~\wb0m_data_i[25]_pad  ;
  assign n4391 = ~n3406 & n4390 ;
  assign n4392 = ~n4389 & ~n4391 ;
  assign n4393 = ~n3474 & n3942 ;
  assign n4394 = \wb0_cyc_i_pad  & ~\wb0m_data_i[26]_pad  ;
  assign n4395 = ~n3406 & n4394 ;
  assign n4396 = ~n4393 & ~n4395 ;
  assign n4397 = ~n3474 & n3951 ;
  assign n4398 = \wb0_cyc_i_pad  & ~\wb0m_data_i[27]_pad  ;
  assign n4399 = ~n3406 & n4398 ;
  assign n4400 = ~n4397 & ~n4399 ;
  assign n4401 = ~n3474 & n3960 ;
  assign n4402 = \wb0_cyc_i_pad  & ~\wb0m_data_i[28]_pad  ;
  assign n4403 = ~n3406 & n4402 ;
  assign n4404 = ~n4401 & ~n4403 ;
  assign n4405 = ~n3474 & n3969 ;
  assign n4406 = \wb0_cyc_i_pad  & ~\wb0m_data_i[29]_pad  ;
  assign n4407 = ~n3406 & n4406 ;
  assign n4408 = ~n4405 & ~n4407 ;
  assign n4409 = ~n3474 & n3978 ;
  assign n4410 = \wb0_cyc_i_pad  & ~\wb0m_data_i[2]_pad  ;
  assign n4411 = ~n3406 & n4410 ;
  assign n4412 = ~n4409 & ~n4411 ;
  assign n4413 = ~n3474 & n3992 ;
  assign n4414 = \wb0_cyc_i_pad  & ~\wb0m_data_i[30]_pad  ;
  assign n4415 = ~n3406 & n4414 ;
  assign n4416 = ~n4413 & ~n4415 ;
  assign n4417 = ~n3474 & n4001 ;
  assign n4418 = \wb0_cyc_i_pad  & ~\wb0m_data_i[31]_pad  ;
  assign n4419 = ~n3406 & n4418 ;
  assign n4420 = ~n4417 & ~n4419 ;
  assign n4421 = ~n3474 & n4010 ;
  assign n4422 = \wb0_cyc_i_pad  & ~\wb0m_data_i[3]_pad  ;
  assign n4423 = ~n3406 & n4422 ;
  assign n4424 = ~n4421 & ~n4423 ;
  assign n4425 = ~n3474 & n4024 ;
  assign n4426 = \wb0_cyc_i_pad  & ~\wb0m_data_i[4]_pad  ;
  assign n4427 = ~n3406 & n4426 ;
  assign n4428 = ~n4425 & ~n4427 ;
  assign n4429 = ~n3474 & n4038 ;
  assign n4430 = \wb0_cyc_i_pad  & ~\wb0m_data_i[5]_pad  ;
  assign n4431 = ~n3406 & n4430 ;
  assign n4432 = ~n4429 & ~n4431 ;
  assign n4433 = ~n3474 & n4052 ;
  assign n4434 = \wb0_cyc_i_pad  & ~\wb0m_data_i[6]_pad  ;
  assign n4435 = ~n3406 & n4434 ;
  assign n4436 = ~n4433 & ~n4435 ;
  assign n4437 = ~n3474 & n4066 ;
  assign n4438 = \wb0_cyc_i_pad  & ~\wb0m_data_i[7]_pad  ;
  assign n4439 = ~n3406 & n4438 ;
  assign n4440 = ~n4437 & ~n4439 ;
  assign n4441 = ~n3474 & n4080 ;
  assign n4442 = \wb0_cyc_i_pad  & ~\wb0m_data_i[8]_pad  ;
  assign n4443 = ~n3406 & n4442 ;
  assign n4444 = ~n4441 & ~n4443 ;
  assign n4445 = ~n3474 & n4094 ;
  assign n4446 = \wb0_cyc_i_pad  & ~\wb0m_data_i[9]_pad  ;
  assign n4447 = ~n3406 & n4446 ;
  assign n4448 = ~n4445 & ~n4447 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g22594/_0_  = ~n764 ;
  assign \g22595/_0_  = ~n789 ;
  assign \g22599/_0_  = ~n796 ;
  assign \g22600/_0_  = ~n804 ;
  assign \g22606/_0_  = ~n811 ;
  assign \g22607/_0_  = ~n818 ;
  assign \g22610/_0_  = ~n826 ;
  assign \g22614/_0_  = ~n835 ;
  assign \g22615/_0_  = ~n844 ;
  assign \g22616/_0_  = ~n850 ;
  assign \g22619/_0_  = ~n855 ;
  assign \g22620/_0_  = ~n861 ;
  assign \g22626/_0_  = ~n867 ;
  assign \g22635/_0_  = ~n875 ;
  assign \g22650/_0_  = ~n885 ;
  assign \g22651/_0_  = ~n892 ;
  assign \g22692/_0_  = ~n898 ;
  assign \g22727/_0_  = ~n904 ;
  assign \g22729/_3_  = n912 ;
  assign \g22774/_0_  = n982 ;
  assign \g22775/_0_  = n993 ;
  assign \g22776/_0_  = ~n1022 ;
  assign \g22777/_0_  = ~n1035 ;
  assign \g22779/_3_  = ~n1043 ;
  assign \g22780/_0_  = ~n1050 ;
  assign \g22781/_0_  = ~n1057 ;
  assign \g22782/_0_  = ~n1064 ;
  assign \g22784/_0_  = ~n1071 ;
  assign \g22785/_0_  = ~n1078 ;
  assign \g22786/_0_  = ~n1083 ;
  assign \g22787/_0_  = ~n1088 ;
  assign \g22789/_3_  = ~n1095 ;
  assign \g22790/_0_  = ~n1100 ;
  assign \g22791/_0_  = ~n1105 ;
  assign \g22792/_0_  = ~n1112 ;
  assign \g22793/_0_  = ~n1119 ;
  assign \g22794/_0_  = ~n1126 ;
  assign \g22795/_0_  = ~n1133 ;
  assign \g22796/_0_  = ~n1140 ;
  assign \g22797/_0_  = ~n1147 ;
  assign \g22798/_0_  = ~n1154 ;
  assign \g22799/_0_  = ~n1161 ;
  assign \g22838/_0_  = ~n981 ;
  assign \g22839/_0_  = n1172 ;
  assign \g22841/_0_  = ~n1179 ;
  assign \g22842/_0_  = ~n1184 ;
  assign \g22847/_0_  = ~n1190 ;
  assign \g22848/_0_  = ~n1196 ;
  assign \g22849/_0_  = ~n1202 ;
  assign \g22850/_0_  = ~n1208 ;
  assign \g22851/_0_  = ~n1214 ;
  assign \g22852/_0_  = ~n1220 ;
  assign \g22853/_0_  = ~n1226 ;
  assign \g22854/_0_  = ~n1232 ;
  assign \g22855/_0_  = ~n1238 ;
  assign \g22856/_0_  = ~n1244 ;
  assign \g22857/_0_  = ~n1250 ;
  assign \g22858/_0_  = ~n1256 ;
  assign \g22859/_0_  = ~n1262 ;
  assign \g22860/_0_  = ~n1268 ;
  assign \g22861/_0_  = ~n1274 ;
  assign \g22862/_0_  = ~n1280 ;
  assign \g22863/_0_  = ~n1286 ;
  assign \g22864/_0_  = ~n1292 ;
  assign \g22865/_0_  = ~n1298 ;
  assign \g22867/_0_  = ~n1304 ;
  assign \g22868/_0_  = ~n1310 ;
  assign \g22869/_0_  = ~n1316 ;
  assign \g22871/_0_  = ~n1322 ;
  assign \g22872/_0_  = ~n1328 ;
  assign \g22873/_0_  = ~n1334 ;
  assign \g22874/_0_  = ~n1340 ;
  assign \g22875/_0_  = ~n1346 ;
  assign \g22876/_0_  = ~n1352 ;
  assign \g22878/_0_  = n1374 ;
  assign \g22882/_2_  = ~n1171 ;
  assign \g22995/_0_  = ~n1402 ;
  assign \g23030/_0_  = ~n1420 ;
  assign \g23046/_0_  = ~n1428 ;
  assign \g23077/_0_  = ~n1435 ;
  assign \g23111/_0_  = n1436 ;
  assign \g23115/_1_  = ~n1449 ;
  assign \g23124/_2_  = ~n1451 ;
  assign \g23126/_2_  = ~n1453 ;
  assign \g23128/_2_  = ~n1455 ;
  assign \g23130/_2_  = ~n1457 ;
  assign \g23132/_2_  = ~n1459 ;
  assign \g23134/_2_  = ~n1461 ;
  assign \g23136/_2_  = ~n1463 ;
  assign \g23137/_0_  = ~n1465 ;
  assign \g23140/_2_  = ~n1467 ;
  assign \g23142/_2_  = ~n1469 ;
  assign \g23144/_2_  = ~n1471 ;
  assign \g23146/_2_  = ~n1473 ;
  assign \g23148/_2_  = ~n1475 ;
  assign \g23150/_2_  = ~n1477 ;
  assign \g23152/_2_  = ~n1479 ;
  assign \g23154/_2_  = ~n1481 ;
  assign \g23156/_2_  = ~n1483 ;
  assign \g23158/_2_  = ~n1485 ;
  assign \g23160/_2_  = ~n1487 ;
  assign \g23162/_2_  = ~n1489 ;
  assign \g23163/_3_  = ~n1491 ;
  assign \g23164/_0_  = ~n1493 ;
  assign \g23166/_0_  = ~n1495 ;
  assign \g23168/_0_  = ~n1497 ;
  assign \g23170/_2_  = ~n1499 ;
  assign \g23172/_2_  = ~n1501 ;
  assign \g23174/_2_  = ~n1503 ;
  assign \g23175/_0_  = ~n1505 ;
  assign \g23177/_0_  = ~n1507 ;
  assign \g23180/_2_  = ~n1509 ;
  assign \g23220/_0_  = ~n1518 ;
  assign \g23238/_0_  = ~n1525 ;
  assign \g23239/_0_  = ~n1532 ;
  assign \g23240/_0_  = ~n1539 ;
  assign \g23241/_0_  = ~n1546 ;
  assign \g23242/_0_  = ~n1553 ;
  assign \g23243/_0_  = ~n1560 ;
  assign \g23244/_0_  = ~n1567 ;
  assign \g23245/_0_  = ~n1574 ;
  assign \g23247/_3_  = ~n1581 ;
  assign \g23248/_0_  = ~n1588 ;
  assign \g23249/_0_  = ~n1595 ;
  assign \g23250/_0_  = ~n1602 ;
  assign \g23251/_0_  = ~n1609 ;
  assign \g23252/_0_  = ~n1616 ;
  assign \g23253/_0_  = ~n1623 ;
  assign \g23255/_3_  = ~n1630 ;
  assign \g23260/_0_  = n1632 ;
  assign \g23284/_3_  = n1634 ;
  assign \g23285/_0_  = ~n1637 ;
  assign \g23334/_0_  = ~n1646 ;
  assign \g23343/_0_  = n1635 ;
  assign \g23366/_0_  = ~n1659 ;
  assign \g23402/_0_  = n1660 ;
  assign \g23403/_0_  = ~n1674 ;
  assign \g23404/_0_  = n1681 ;
  assign \g23405/_0_  = ~n1687 ;
  assign \g23407/_0_  = ~n1695 ;
  assign \g23408/_0_  = n1702 ;
  assign \g23409/_0_  = ~n1708 ;
  assign \g23410/_0_  = ~n1714 ;
  assign \g23411/_0_  = ~n1722 ;
  assign \g23413/_2_  = ~n1727 ;
  assign \g23415/_2_  = ~n1732 ;
  assign \g23417/_2_  = n1737 ;
  assign \g23542/_0_  = n1162 ;
  assign \g23607/_0_  = ~n1753 ;
  assign \g23608/_0_  = ~n1774 ;
  assign \g23609/_3_  = ~n1786 ;
  assign \g23707/_0_  = ~n1797 ;
  assign \g23708/_0_  = ~n1808 ;
  assign \g23709/_0_  = ~n1819 ;
  assign \g23710/_0_  = ~n1830 ;
  assign \g23711/_0_  = ~n1841 ;
  assign \g23712/_0_  = ~n1852 ;
  assign \g23713/_0_  = ~n1863 ;
  assign \g23714/_0_  = ~n1874 ;
  assign \g23715/_0_  = ~n1885 ;
  assign \g23716/_0_  = ~n1896 ;
  assign \g23754/_0_  = ~n1902 ;
  assign \g23755/_0_  = ~n1907 ;
  assign \g23756/_0_  = ~n1913 ;
  assign \g23757/_0_  = ~n1919 ;
  assign \g23758/_0_  = ~n1924 ;
  assign \g23759/_0_  = ~n1930 ;
  assign \g23760/_0_  = ~n1939 ;
  assign \g23761/_0_  = n1946 ;
  assign \g23763/_3_  = n1954 ;
  assign \g23767/_0_  = n1970 ;
  assign \g23768/_0_  = n1986 ;
  assign \g23833/_0_  = ~n2031 ;
  assign \g23837/_0_  = ~n2046 ;
  assign \g23838/_0_  = ~n2060 ;
  assign \g23839/_0_  = ~n2074 ;
  assign \g23840/_0_  = ~n2088 ;
  assign \g23841/_0_  = ~n2102 ;
  assign \g23842/_0_  = ~n2116 ;
  assign \g23843/_0_  = ~n2130 ;
  assign \g23844/_0_  = ~n2145 ;
  assign \g23845/_0_  = ~n2160 ;
  assign \g23849/_3_  = n2164 ;
  assign \g23851/_3_  = n2168 ;
  assign \g23858/_0_  = ~n2192 ;
  assign \g23870/_0_  = n2197 ;
  assign \g23871/_0_  = n2202 ;
  assign \g23872/_3_  = n2218 ;
  assign \g23873/_3_  = n2230 ;
  assign \g23874/_3_  = n2242 ;
  assign \g23875/_3_  = n2254 ;
  assign \g23876/_3_  = n2266 ;
  assign \g23877/_3_  = n2278 ;
  assign \g23878/_3_  = n2290 ;
  assign \g23879/_3_  = n2302 ;
  assign \g23880/_3_  = n2314 ;
  assign \g23881/_3_  = n2326 ;
  assign \g23882/_3_  = n2338 ;
  assign \g23883/_3_  = n2350 ;
  assign \g23884/_3_  = n2362 ;
  assign \g23885/_3_  = n2374 ;
  assign \g23886/_3_  = n2386 ;
  assign \g23887/_3_  = n2398 ;
  assign \g23888/_3_  = n2410 ;
  assign \g23889/_3_  = n2422 ;
  assign \g23890/_3_  = n2434 ;
  assign \g23891/_3_  = n2446 ;
  assign \g23892/_3_  = n2463 ;
  assign \g23893/_3_  = n2476 ;
  assign \g23894/_3_  = n2489 ;
  assign \g23895/_3_  = n2502 ;
  assign \g23896/_3_  = n2515 ;
  assign \g23897/_3_  = n2528 ;
  assign \g23898/_3_  = n2541 ;
  assign \g23899/_3_  = n2554 ;
  assign \g23900/_3_  = n2567 ;
  assign \g23901/_3_  = n2580 ;
  assign \g23902/_3_  = n2593 ;
  assign \g23903/_3_  = n2606 ;
  assign \g23904/_3_  = n2619 ;
  assign \g23905/_3_  = n2632 ;
  assign \g23906/_3_  = n2645 ;
  assign \g23907/_3_  = n2658 ;
  assign \g23908/_3_  = n2671 ;
  assign \g23909/_3_  = n2684 ;
  assign \g23910/_3_  = n2697 ;
  assign \g23911/_3_  = n2710 ;
  assign \g23912/_3_  = ~n2724 ;
  assign \g23913/_3_  = ~n2733 ;
  assign \g23914/_3_  = ~n2742 ;
  assign \g23915/_3_  = ~n2751 ;
  assign \g23959/_0_  = ~n2763 ;
  assign \g23961/_0_  = ~n2772 ;
  assign \g23962/_0_  = ~n2781 ;
  assign \g23966/_0_  = ~n2790 ;
  assign \g23967/_0_  = ~n2799 ;
  assign \g23969/_0_  = ~n2808 ;
  assign \g23970/_0_  = ~n2817 ;
  assign \g23971/_0_  = ~n2826 ;
  assign \g23972/_0_  = ~n2835 ;
  assign \g23979/_0_  = ~n2844 ;
  assign \g23987/_0_  = ~n2856 ;
  assign \g23988/_0_  = ~n2868 ;
  assign \g23989/_0_  = ~n2880 ;
  assign \g23990/_0_  = ~n2892 ;
  assign \g24005/_0_  = ~n2902 ;
  assign \g24010/_0_  = n933 ;
  assign \g24012/_0_  = ~n2912 ;
  assign \g24013/_0_  = ~n2922 ;
  assign \g24014/_0_  = ~n2932 ;
  assign \g24015/_0_  = ~n2942 ;
  assign \g24016/_0_  = ~n2952 ;
  assign \g24017/_0_  = ~n2962 ;
  assign \g24018/_0_  = ~n2972 ;
  assign \g24019/_0_  = ~n2982 ;
  assign \g24020/_0_  = ~n2992 ;
  assign \g24026/_0_  = ~n3008 ;
  assign \g24027/_0_  = ~n3024 ;
  assign \g24028/_0_  = ~n3040 ;
  assign \g24029/_0_  = ~n3056 ;
  assign \g24030/_0_  = ~n3072 ;
  assign \g24031/_0_  = ~n3088 ;
  assign \g24032/_0_  = ~n3102 ;
  assign \g24033/_0_  = ~n3118 ;
  assign \g24034/_0_  = ~n3134 ;
  assign \g24035/_0_  = ~n3150 ;
  assign \g24036/_0_  = ~n3166 ;
  assign \g24037/_0_  = ~n3182 ;
  assign \g24038/_0_  = ~n3198 ;
  assign \g24039/_0_  = ~n3214 ;
  assign \g24042/_0_  = ~n3222 ;
  assign \g24049/_0_  = ~n3229 ;
  assign \g24063/_0_  = n3233 ;
  assign \g24119/_0_  = n3235 ;
  assign \g24120/_0_  = n3237 ;
  assign \g24357/_0_  = ~n1638 ;
  assign \g24432/_0_  = n3240 ;
  assign \g24433/_0_  = n3243 ;
  assign \g24437/_0_  = n3246 ;
  assign \g24438/_0_  = n3249 ;
  assign \g24477/_0_  = ~n3251 ;
  assign \g24491/_0_  = ~n3259 ;
  assign \g24530/_2_  = n3266 ;
  assign \g24532/_0_  = n3268 ;
  assign \g24534/_0_  = ~n3275 ;
  assign \g24537/_0_  = n3280 ;
  assign \g24538/_0_  = n3285 ;
  assign \g24539/_0_  = n3287 ;
  assign \g24540/_0_  = n3289 ;
  assign \g24606/_2_  = n3293 ;
  assign \g24612/_0_  = n3294 ;
  assign \g24677/_0_  = ~n3298 ;
  assign \g24678/_0_  = ~n3302 ;
  assign \g24679/_0_  = ~n3306 ;
  assign \g24688/_0_  = ~n3310 ;
  assign \g24743/_0_  = n3312 ;
  assign \g24847/_0_  = n3315 ;
  assign \g24849/_0_  = ~n3321 ;
  assign \g24850/_0_  = ~n3324 ;
  assign \g24854/_0_  = ~n3327 ;
  assign \g24862/_0_  = ~n3330 ;
  assign \g24872/_0_  = ~n3333 ;
  assign \g24873/_0_  = ~n3336 ;
  assign \g24874/_0_  = ~n3339 ;
  assign \g24876/_0_  = ~n3342 ;
  assign \g24879/_0_  = ~n3347 ;
  assign \g24880/_0_  = n3350 ;
  assign \g24881/_0_  = n3352 ;
  assign \g24882/_0_  = n3354 ;
  assign \g24952/_2_  = n1362 ;
  assign \g24976/_1_  = n1757 ;
  assign \g25003/_0_  = n3358 ;
  assign \g25004/_0_  = n3360 ;
  assign \g25005/_0_  = n3362 ;
  assign \g25006/_0_  = n3366 ;
  assign \g25011/_0_  = ~n3370 ;
  assign \g25012/_0_  = ~n3373 ;
  assign \g25013/_0_  = ~n3377 ;
  assign \g25031/_0_  = ~n3380 ;
  assign \g25032/_0_  = ~n3383 ;
  assign \g25033/_0_  = ~n3386 ;
  assign \g25034/_0_  = ~n3389 ;
  assign \g25035/_0_  = ~n3392 ;
  assign \g25153/_2_  = n3318 ;
  assign \g25183/_0_  = n3394 ;
  assign \g25184/_0_  = n3396 ;
  assign \g25224/_0_  = n3403 ;
  assign \g25232/_0_  = n3411 ;
  assign \g25237/_0_  = n3414 ;
  assign \g25241/_2_  = n2178 ;
  assign \g25243/_2_  = n2180 ;
  assign \g25248/_3_  = n3367 ;
  assign \g25261/_0_  = n3416 ;
  assign \g25262/_0_  = n3418 ;
  assign \g25266/_3_  = n3421 ;
  assign \g25267/_0_  = n3423 ;
  assign \g25269/_0_  = n3425 ;
  assign \g25543/_1_  = n3426 ;
  assign \g25602/_3_  = n3428 ;
  assign \g25610/_0_  = n3430 ;
  assign \g25611/_0_  = n3432 ;
  assign \g25841/_0_  = n3433 ;
  assign \g25843/_0_  = n3434 ;
  assign \g25893/_0_  = n3435 ;
  assign \g27013/_0_  = ~n3440 ;
  assign \g27060/_0_  = ~n3445 ;
  assign \g27073/_0_  = ~n3452 ;
  assign \g27184/_0_  = ~n973 ;
  assign \g27186/_0_  = ~n942 ;
  assign \g27189/_2_  = ~n946 ;
  assign \g47/_0_  = ~n3468 ;
  assign \u0_u0_ch_done_reg/_05_  = ~n3471 ;
  assign \u2_adr0_cnt_reg[0]/P0000  = ~\u2_adr0_cnt_reg[0]/P0001  ;
  assign \u2_adr1_cnt_reg[0]/P0000  = ~\u2_adr1_cnt_reg[0]/P0001  ;
  assign \u3_u0_mast_we_r_reg/_05_  = n3473 ;
  assign \wb0_ack_o_pad  = ~n3478 ;
  assign \wb0_addr_o[0]_pad  = n3480 ;
  assign \wb0_addr_o[10]_pad  = ~n3485 ;
  assign \wb0_addr_o[11]_pad  = ~n3489 ;
  assign \wb0_addr_o[12]_pad  = ~n3493 ;
  assign \wb0_addr_o[13]_pad  = ~n3497 ;
  assign \wb0_addr_o[14]_pad  = ~n3501 ;
  assign \wb0_addr_o[15]_pad  = ~n3505 ;
  assign \wb0_addr_o[16]_pad  = ~n3509 ;
  assign \wb0_addr_o[17]_pad  = ~n3513 ;
  assign \wb0_addr_o[18]_pad  = ~n3517 ;
  assign \wb0_addr_o[19]_pad  = ~n3521 ;
  assign \wb0_addr_o[1]_pad  = n3523 ;
  assign \wb0_addr_o[20]_pad  = ~n3527 ;
  assign \wb0_addr_o[21]_pad  = ~n3531 ;
  assign \wb0_addr_o[22]_pad  = ~n3535 ;
  assign \wb0_addr_o[23]_pad  = ~n3539 ;
  assign \wb0_addr_o[24]_pad  = ~n3543 ;
  assign \wb0_addr_o[25]_pad  = ~n3547 ;
  assign \wb0_addr_o[26]_pad  = ~n3551 ;
  assign \wb0_addr_o[27]_pad  = ~n3555 ;
  assign \wb0_addr_o[28]_pad  = n3560 ;
  assign \wb0_addr_o[29]_pad  = n3565 ;
  assign \wb0_addr_o[2]_pad  = ~n3569 ;
  assign \wb0_addr_o[30]_pad  = n3574 ;
  assign \wb0_addr_o[31]_pad  = n3579 ;
  assign \wb0_addr_o[3]_pad  = ~n3583 ;
  assign \wb0_addr_o[4]_pad  = ~n3587 ;
  assign \wb0_addr_o[5]_pad  = ~n3591 ;
  assign \wb0_addr_o[6]_pad  = ~n3595 ;
  assign \wb0_addr_o[7]_pad  = ~n3599 ;
  assign \wb0_addr_o[8]_pad  = ~n3603 ;
  assign \wb0_addr_o[9]_pad  = ~n3607 ;
  assign \wb0_cyc_o_pad  = ~n3608 ;
  assign \wb0_err_o_pad  = n3610 ;
  assign \wb0_rty_o_pad  = n3612 ;
  assign \wb0_sel_o[0]_pad  = ~n3614 ;
  assign \wb0_sel_o[1]_pad  = ~n3616 ;
  assign \wb0_sel_o[2]_pad  = ~n3618 ;
  assign \wb0_sel_o[3]_pad  = ~n3620 ;
  assign \wb0_stb_o_pad  = ~n3624 ;
  assign \wb0_we_o_pad  = ~n3627 ;
  assign \wb0m_data_o[0]_pad  = ~n3631 ;
  assign \wb0m_data_o[10]_pad  = ~n3635 ;
  assign \wb0m_data_o[11]_pad  = ~n3639 ;
  assign \wb0m_data_o[12]_pad  = ~n3643 ;
  assign \wb0m_data_o[13]_pad  = ~n3647 ;
  assign \wb0m_data_o[14]_pad  = ~n3651 ;
  assign \wb0m_data_o[15]_pad  = ~n3655 ;
  assign \wb0m_data_o[16]_pad  = ~n3659 ;
  assign \wb0m_data_o[17]_pad  = ~n3663 ;
  assign \wb0m_data_o[18]_pad  = ~n3667 ;
  assign \wb0m_data_o[19]_pad  = ~n3671 ;
  assign \wb0m_data_o[1]_pad  = ~n3675 ;
  assign \wb0m_data_o[20]_pad  = ~n3679 ;
  assign \wb0m_data_o[21]_pad  = ~n3683 ;
  assign \wb0m_data_o[22]_pad  = ~n3687 ;
  assign \wb0m_data_o[23]_pad  = ~n3691 ;
  assign \wb0m_data_o[24]_pad  = ~n3695 ;
  assign \wb0m_data_o[25]_pad  = ~n3699 ;
  assign \wb0m_data_o[26]_pad  = ~n3703 ;
  assign \wb0m_data_o[27]_pad  = ~n3707 ;
  assign \wb0m_data_o[28]_pad  = ~n3711 ;
  assign \wb0m_data_o[29]_pad  = ~n3715 ;
  assign \wb0m_data_o[2]_pad  = ~n3719 ;
  assign \wb0m_data_o[30]_pad  = ~n3723 ;
  assign \wb0m_data_o[31]_pad  = ~n3727 ;
  assign \wb0m_data_o[3]_pad  = ~n3731 ;
  assign \wb0m_data_o[4]_pad  = ~n3735 ;
  assign \wb0m_data_o[5]_pad  = ~n3739 ;
  assign \wb0m_data_o[6]_pad  = ~n3743 ;
  assign \wb0m_data_o[7]_pad  = ~n3747 ;
  assign \wb0m_data_o[8]_pad  = ~n3751 ;
  assign \wb0m_data_o[9]_pad  = ~n3755 ;
  assign \wb0s_data_o[0]_pad  = ~n3769 ;
  assign \wb0s_data_o[10]_pad  = ~n3783 ;
  assign \wb0s_data_o[11]_pad  = ~n3797 ;
  assign \wb0s_data_o[12]_pad  = ~n3806 ;
  assign \wb0s_data_o[13]_pad  = ~n3815 ;
  assign \wb0s_data_o[14]_pad  = ~n3824 ;
  assign \wb0s_data_o[15]_pad  = ~n3833 ;
  assign \wb0s_data_o[16]_pad  = ~n3842 ;
  assign \wb0s_data_o[17]_pad  = ~n3851 ;
  assign \wb0s_data_o[18]_pad  = ~n3860 ;
  assign \wb0s_data_o[19]_pad  = ~n3869 ;
  assign \wb0s_data_o[1]_pad  = ~n3883 ;
  assign \wb0s_data_o[20]_pad  = ~n3892 ;
  assign \wb0s_data_o[21]_pad  = ~n3901 ;
  assign \wb0s_data_o[22]_pad  = ~n3910 ;
  assign \wb0s_data_o[23]_pad  = ~n3919 ;
  assign \wb0s_data_o[24]_pad  = ~n3928 ;
  assign \wb0s_data_o[25]_pad  = ~n3937 ;
  assign \wb0s_data_o[26]_pad  = ~n3946 ;
  assign \wb0s_data_o[27]_pad  = ~n3955 ;
  assign \wb0s_data_o[28]_pad  = ~n3964 ;
  assign \wb0s_data_o[29]_pad  = ~n3973 ;
  assign \wb0s_data_o[2]_pad  = ~n3987 ;
  assign \wb0s_data_o[30]_pad  = ~n3996 ;
  assign \wb0s_data_o[31]_pad  = ~n4005 ;
  assign \wb0s_data_o[3]_pad  = ~n4019 ;
  assign \wb0s_data_o[4]_pad  = ~n4033 ;
  assign \wb0s_data_o[5]_pad  = ~n4047 ;
  assign \wb0s_data_o[6]_pad  = ~n4061 ;
  assign \wb0s_data_o[7]_pad  = ~n4075 ;
  assign \wb0s_data_o[8]_pad  = ~n4089 ;
  assign \wb0s_data_o[9]_pad  = ~n4103 ;
  assign \wb1_ack_o_pad  = ~n4107 ;
  assign \wb1_addr_o[0]_pad  = n4109 ;
  assign \wb1_addr_o[10]_pad  = ~n4113 ;
  assign \wb1_addr_o[11]_pad  = ~n4117 ;
  assign \wb1_addr_o[12]_pad  = ~n4121 ;
  assign \wb1_addr_o[13]_pad  = ~n4125 ;
  assign \wb1_addr_o[14]_pad  = ~n4129 ;
  assign \wb1_addr_o[15]_pad  = ~n4133 ;
  assign \wb1_addr_o[16]_pad  = ~n4137 ;
  assign \wb1_addr_o[17]_pad  = ~n4141 ;
  assign \wb1_addr_o[18]_pad  = ~n4145 ;
  assign \wb1_addr_o[19]_pad  = ~n4149 ;
  assign \wb1_addr_o[1]_pad  = n4151 ;
  assign \wb1_addr_o[20]_pad  = ~n4155 ;
  assign \wb1_addr_o[21]_pad  = ~n4159 ;
  assign \wb1_addr_o[22]_pad  = ~n4163 ;
  assign \wb1_addr_o[23]_pad  = ~n4167 ;
  assign \wb1_addr_o[24]_pad  = ~n4171 ;
  assign \wb1_addr_o[25]_pad  = ~n4175 ;
  assign \wb1_addr_o[26]_pad  = ~n4179 ;
  assign \wb1_addr_o[27]_pad  = ~n4183 ;
  assign \wb1_addr_o[28]_pad  = n4188 ;
  assign \wb1_addr_o[29]_pad  = n4193 ;
  assign \wb1_addr_o[2]_pad  = ~n4197 ;
  assign \wb1_addr_o[30]_pad  = n4202 ;
  assign \wb1_addr_o[31]_pad  = n4207 ;
  assign \wb1_addr_o[3]_pad  = ~n4211 ;
  assign \wb1_addr_o[4]_pad  = ~n4215 ;
  assign \wb1_addr_o[5]_pad  = ~n4219 ;
  assign \wb1_addr_o[6]_pad  = ~n4223 ;
  assign \wb1_addr_o[7]_pad  = ~n4227 ;
  assign \wb1_addr_o[8]_pad  = ~n4231 ;
  assign \wb1_addr_o[9]_pad  = ~n4235 ;
  assign \wb1_cyc_o_pad  = ~n4236 ;
  assign \wb1_err_o_pad  = n4238 ;
  assign \wb1_rty_o_pad  = n4240 ;
  assign \wb1_sel_o[0]_pad  = ~n4242 ;
  assign \wb1_sel_o[1]_pad  = ~n4244 ;
  assign \wb1_sel_o[2]_pad  = ~n4246 ;
  assign \wb1_sel_o[3]_pad  = ~n4248 ;
  assign \wb1_stb_o_pad  = ~n4252 ;
  assign \wb1_we_o_pad  = ~n4256 ;
  assign \wb1m_data_o[0]_pad  = n4258 ;
  assign \wb1m_data_o[10]_pad  = n4260 ;
  assign \wb1m_data_o[11]_pad  = n4262 ;
  assign \wb1m_data_o[12]_pad  = n4264 ;
  assign \wb1m_data_o[13]_pad  = n4266 ;
  assign \wb1m_data_o[14]_pad  = n4268 ;
  assign \wb1m_data_o[15]_pad  = n4270 ;
  assign \wb1m_data_o[16]_pad  = n4272 ;
  assign \wb1m_data_o[17]_pad  = n4274 ;
  assign \wb1m_data_o[18]_pad  = n4276 ;
  assign \wb1m_data_o[19]_pad  = n4278 ;
  assign \wb1m_data_o[1]_pad  = n4280 ;
  assign \wb1m_data_o[20]_pad  = n4282 ;
  assign \wb1m_data_o[21]_pad  = n4284 ;
  assign \wb1m_data_o[22]_pad  = n4286 ;
  assign \wb1m_data_o[23]_pad  = n4288 ;
  assign \wb1m_data_o[24]_pad  = n4290 ;
  assign \wb1m_data_o[25]_pad  = n4292 ;
  assign \wb1m_data_o[26]_pad  = n4294 ;
  assign \wb1m_data_o[27]_pad  = n4296 ;
  assign \wb1m_data_o[28]_pad  = n4298 ;
  assign \wb1m_data_o[29]_pad  = n4300 ;
  assign \wb1m_data_o[2]_pad  = n4302 ;
  assign \wb1m_data_o[30]_pad  = n4304 ;
  assign \wb1m_data_o[31]_pad  = n4306 ;
  assign \wb1m_data_o[3]_pad  = n4308 ;
  assign \wb1m_data_o[4]_pad  = n4310 ;
  assign \wb1m_data_o[5]_pad  = n4312 ;
  assign \wb1m_data_o[6]_pad  = n4314 ;
  assign \wb1m_data_o[7]_pad  = n4316 ;
  assign \wb1m_data_o[8]_pad  = n4318 ;
  assign \wb1m_data_o[9]_pad  = n4320 ;
  assign \wb1s_data_o[0]_pad  = n4324 ;
  assign \wb1s_data_o[10]_pad  = n4328 ;
  assign \wb1s_data_o[11]_pad  = n4332 ;
  assign \wb1s_data_o[12]_pad  = n4336 ;
  assign \wb1s_data_o[13]_pad  = n4340 ;
  assign \wb1s_data_o[14]_pad  = n4344 ;
  assign \wb1s_data_o[15]_pad  = n4348 ;
  assign \wb1s_data_o[16]_pad  = n4352 ;
  assign \wb1s_data_o[17]_pad  = n4356 ;
  assign \wb1s_data_o[18]_pad  = n4360 ;
  assign \wb1s_data_o[19]_pad  = n4364 ;
  assign \wb1s_data_o[1]_pad  = n4368 ;
  assign \wb1s_data_o[20]_pad  = n4372 ;
  assign \wb1s_data_o[21]_pad  = n4376 ;
  assign \wb1s_data_o[22]_pad  = n4380 ;
  assign \wb1s_data_o[23]_pad  = n4384 ;
  assign \wb1s_data_o[24]_pad  = n4388 ;
  assign \wb1s_data_o[25]_pad  = n4392 ;
  assign \wb1s_data_o[26]_pad  = n4396 ;
  assign \wb1s_data_o[27]_pad  = n4400 ;
  assign \wb1s_data_o[28]_pad  = n4404 ;
  assign \wb1s_data_o[29]_pad  = n4408 ;
  assign \wb1s_data_o[2]_pad  = n4412 ;
  assign \wb1s_data_o[30]_pad  = n4416 ;
  assign \wb1s_data_o[31]_pad  = n4420 ;
  assign \wb1s_data_o[3]_pad  = n4424 ;
  assign \wb1s_data_o[4]_pad  = n4428 ;
  assign \wb1s_data_o[5]_pad  = n4432 ;
  assign \wb1s_data_o[6]_pad  = n4436 ;
  assign \wb1s_data_o[7]_pad  = n4440 ;
  assign \wb1s_data_o[8]_pad  = n4444 ;
  assign \wb1s_data_o[9]_pad  = n4448 ;
endmodule
