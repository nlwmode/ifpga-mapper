module top( \a0_pad  , a_pad , b_pad , c_pad , \d0_pad  , d_pad , e_pad , f_pad , g_pad , h_pad , j_pad , k_pad , l_pad , m_pad , n_pad , o_pad , p_pad , q_pad , s_pad , t_pad , u_pad , v_pad , w_pad , x_pad , y_pad , z_pad , \b0_pad  , \c0_pad  , \e0_pad  , \f0_pad  , \g0_pad  , \h0_pad  , \i0_pad  , \j0_pad  , \k0_pad  , \l0_pad  , \m0_pad  , \n0_pad  , \o0_pad  , \p0_pad  , \q0_pad  , \r0_pad  , \s0_pad  , \t0_pad  );
  input \a0_pad  ;
  input a_pad ;
  input b_pad ;
  input c_pad ;
  input \d0_pad  ;
  input d_pad ;
  input e_pad ;
  input f_pad ;
  input g_pad ;
  input h_pad ;
  input j_pad ;
  input k_pad ;
  input l_pad ;
  input m_pad ;
  input n_pad ;
  input o_pad ;
  input p_pad ;
  input q_pad ;
  input s_pad ;
  input t_pad ;
  input u_pad ;
  input v_pad ;
  input w_pad ;
  input x_pad ;
  input y_pad ;
  input z_pad ;
  output \b0_pad  ;
  output \c0_pad  ;
  output \e0_pad  ;
  output \f0_pad  ;
  output \g0_pad  ;
  output \h0_pad  ;
  output \i0_pad  ;
  output \j0_pad  ;
  output \k0_pad  ;
  output \l0_pad  ;
  output \m0_pad  ;
  output \n0_pad  ;
  output \o0_pad  ;
  output \p0_pad  ;
  output \q0_pad  ;
  output \r0_pad  ;
  output \s0_pad  ;
  output \t0_pad  ;
  wire n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 ;
  assign n27 = ~\d0_pad  & j_pad ;
  assign n28 = ~s_pad & ~t_pad ;
  assign n29 = ~u_pad & n28 ;
  assign n30 = ~v_pad & ~n29 ;
  assign n31 = w_pad & x_pad ;
  assign n32 = ~n30 & n31 ;
  assign n33 = ~y_pad & ~n32 ;
  assign n34 = ~\a0_pad  & n33 ;
  assign n36 = ~\a0_pad  & ~z_pad ;
  assign n35 = e_pad & f_pad ;
  assign n37 = ~h_pad & ~n35 ;
  assign n38 = ~n36 & n37 ;
  assign n39 = ~n34 & n38 ;
  assign n40 = z_pad & ~n33 ;
  assign n41 = ~\a0_pad  & ~n40 ;
  assign n44 = c_pad & ~m_pad ;
  assign n45 = ~c_pad & m_pad ;
  assign n52 = ~n44 & ~n45 ;
  assign n49 = a_pad & ~k_pad ;
  assign n50 = ~a_pad & k_pad ;
  assign n53 = ~n49 & ~n50 ;
  assign n54 = n52 & n53 ;
  assign n46 = ~d_pad & ~n_pad ;
  assign n47 = d_pad & n_pad ;
  assign n48 = ~n46 & ~n47 ;
  assign n42 = b_pad & ~l_pad ;
  assign n43 = ~b_pad & l_pad ;
  assign n51 = ~n42 & ~n43 ;
  assign n55 = ~n48 & n51 ;
  assign n56 = n54 & n55 ;
  assign n57 = ~j_pad & ~n56 ;
  assign n58 = ~j_pad & ~o_pad ;
  assign n59 = ~j_pad & p_pad ;
  assign n60 = g_pad & ~j_pad ;
  assign n61 = ~h_pad & ~q_pad ;
  assign n62 = n35 & n61 ;
  assign n63 = ~n35 & n61 ;
  assign n64 = ~s_pad & n63 ;
  assign n65 = s_pad & t_pad ;
  assign n66 = ~n28 & ~n65 ;
  assign n67 = n63 & n66 ;
  assign n68 = ~u_pad & ~n65 ;
  assign n69 = u_pad & n65 ;
  assign n70 = n63 & ~n69 ;
  assign n71 = ~n68 & n70 ;
  assign n74 = v_pad & n70 ;
  assign n72 = u_pad & ~v_pad ;
  assign n73 = n65 & n72 ;
  assign n75 = n63 & ~n73 ;
  assign n76 = ~n74 & n75 ;
  assign n78 = ~w_pad & n73 ;
  assign n77 = w_pad & ~n73 ;
  assign n79 = n63 & ~n77 ;
  assign n80 = ~n78 & n79 ;
  assign n83 = x_pad & ~n78 ;
  assign n81 = ~w_pad & ~x_pad ;
  assign n82 = n73 & n81 ;
  assign n84 = n63 & ~n82 ;
  assign n85 = ~n83 & n84 ;
  assign n87 = ~y_pad & n82 ;
  assign n86 = y_pad & ~n82 ;
  assign n88 = n63 & ~n86 ;
  assign n89 = ~n87 & n88 ;
  assign n91 = ~z_pad & n87 ;
  assign n90 = z_pad & ~n87 ;
  assign n92 = n63 & ~n90 ;
  assign n93 = ~n91 & n92 ;
  assign n94 = \a0_pad  & ~n91 ;
  assign n95 = n36 & n87 ;
  assign n96 = n63 & ~n95 ;
  assign n97 = ~n94 & n96 ;
  assign \b0_pad  = n27 ;
  assign \c0_pad  = ~n39 ;
  assign \e0_pad  = n41 ;
  assign \f0_pad  = n57 ;
  assign \g0_pad  = n58 ;
  assign \h0_pad  = n59 ;
  assign \i0_pad  = ~n60 ;
  assign \j0_pad  = ~n41 ;
  assign \k0_pad  = n62 ;
  assign \l0_pad  = n64 ;
  assign \m0_pad  = n67 ;
  assign \n0_pad  = n71 ;
  assign \o0_pad  = ~n76 ;
  assign \p0_pad  = ~n80 ;
  assign \q0_pad  = ~n85 ;
  assign \r0_pad  = ~n89 ;
  assign \s0_pad  = ~n93 ;
  assign \t0_pad  = ~n97 ;
endmodule
