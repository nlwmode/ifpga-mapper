module top (\1_pad , \2_pad , \3_pad , \4_pad , \5_pad , \6_pad , \7_pad , \8_pad , \44_pad , \45_pad , \46_pad , \47_pad , \48_pad , \49_pad , \50_pad , \51_pad );
	input \1_pad  ;
	input \2_pad  ;
	input \3_pad  ;
	input \4_pad  ;
	input \5_pad  ;
	input \6_pad  ;
	input \7_pad  ;
	input \8_pad  ;
	output \44_pad  ;
	output \45_pad  ;
	output \46_pad  ;
	output \47_pad  ;
	output \48_pad  ;
	output \49_pad  ;
	output \50_pad  ;
	output \51_pad  ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w56_ ;
	wire _w55_ ;
	wire _w54_ ;
	wire _w53_ ;
	wire _w52_ ;
	wire _w51_ ;
	wire _w50_ ;
	wire _w49_ ;
	wire _w48_ ;
	wire _w47_ ;
	wire _w46_ ;
	wire _w45_ ;
	wire _w44_ ;
	wire _w43_ ;
	wire _w42_ ;
	wire _w41_ ;
	wire _w40_ ;
	wire _w39_ ;
	wire _w22_ ;
	wire _w21_ ;
	wire _w20_ ;
	wire _w19_ ;
	wire _w18_ ;
	wire _w17_ ;
	wire _w16_ ;
	wire _w15_ ;
	wire _w14_ ;
	wire _w13_ ;
	wire _w12_ ;
	wire _w11_ ;
	wire _w10_ ;
	wire _w23_ ;
	wire _w24_ ;
	wire _w25_ ;
	wire _w26_ ;
	wire _w27_ ;
	wire _w28_ ;
	wire _w29_ ;
	wire _w30_ ;
	wire _w31_ ;
	wire _w32_ ;
	wire _w33_ ;
	wire _w34_ ;
	wire _w35_ ;
	wire _w36_ ;
	wire _w37_ ;
	wire _w38_ ;
	LUT1 #(
		.INIT('h1)
	) name0 (
		\8_pad ,
		_w10_
	);
	LUT2 #(
		.INIT('h8)
	) name1 (
		\7_pad ,
		\8_pad ,
		_w11_
	);
	LUT3 #(
		.INIT('h06)
	) name2 (
		\1_pad ,
		\3_pad ,
		\4_pad ,
		_w12_
	);
	LUT4 #(
		.INIT('h009a)
	) name3 (
		\1_pad ,
		\2_pad ,
		\3_pad ,
		\4_pad ,
		_w13_
	);
	LUT4 #(
		.INIT('hb830)
	) name4 (
		\6_pad ,
		_w11_,
		_w12_,
		_w13_,
		_w14_
	);
	LUT4 #(
		.INIT('ha600)
	) name5 (
		\1_pad ,
		\2_pad ,
		\3_pad ,
		\4_pad ,
		_w15_
	);
	LUT4 #(
		.INIT('h00ae)
	) name6 (
		\6_pad ,
		_w11_,
		_w12_,
		_w15_,
		_w16_
	);
	LUT4 #(
		.INIT('h9600)
	) name7 (
		\1_pad ,
		\2_pad ,
		\3_pad ,
		\4_pad ,
		_w17_
	);
	LUT4 #(
		.INIT('h0001)
	) name8 (
		\6_pad ,
		_w11_,
		_w12_,
		_w17_,
		_w18_
	);
	LUT4 #(
		.INIT('h5510)
	) name9 (
		\5_pad ,
		_w14_,
		_w16_,
		_w18_,
		_w19_
	);
	LUT3 #(
		.INIT('h90)
	) name10 (
		\1_pad ,
		\3_pad ,
		\4_pad ,
		_w20_
	);
	LUT4 #(
		.INIT('h0096)
	) name11 (
		\1_pad ,
		\2_pad ,
		\3_pad ,
		\4_pad ,
		_w21_
	);
	LUT2 #(
		.INIT('h8)
	) name12 (
		\8_pad ,
		_w21_,
		_w22_
	);
	LUT4 #(
		.INIT('ha0a2)
	) name13 (
		\6_pad ,
		\7_pad ,
		\8_pad ,
		_w13_,
		_w23_
	);
	LUT4 #(
		.INIT('h048c)
	) name14 (
		\6_pad ,
		\7_pad ,
		_w13_,
		_w21_,
		_w24_
	);
	LUT4 #(
		.INIT('h5510)
	) name15 (
		_w20_,
		_w22_,
		_w23_,
		_w24_,
		_w25_
	);
	LUT4 #(
		.INIT('h0001)
	) name16 (
		\6_pad ,
		\7_pad ,
		_w13_,
		_w15_,
		_w26_
	);
	LUT4 #(
		.INIT('h1113)
	) name17 (
		\5_pad ,
		_w19_,
		_w25_,
		_w26_,
		_w27_
	);
	LUT4 #(
		.INIT('he0c0)
	) name18 (
		\3_pad ,
		\5_pad ,
		\7_pad ,
		\8_pad ,
		_w28_
	);
	LUT4 #(
		.INIT('h1737)
	) name19 (
		\3_pad ,
		\5_pad ,
		\7_pad ,
		\8_pad ,
		_w29_
	);
	LUT2 #(
		.INIT('h2)
	) name20 (
		\4_pad ,
		_w29_,
		_w30_
	);
	LUT4 #(
		.INIT('h0026)
	) name21 (
		\3_pad ,
		\5_pad ,
		\7_pad ,
		\8_pad ,
		_w31_
	);
	LUT4 #(
		.INIT('h3f35)
	) name22 (
		\3_pad ,
		\4_pad ,
		\5_pad ,
		\7_pad ,
		_w32_
	);
	LUT3 #(
		.INIT('h8a)
	) name23 (
		\6_pad ,
		_w31_,
		_w32_,
		_w33_
	);
	LUT3 #(
		.INIT('h54)
	) name24 (
		\2_pad ,
		_w30_,
		_w33_,
		_w34_
	);
	LUT3 #(
		.INIT('h07)
	) name25 (
		\3_pad ,
		\5_pad ,
		\6_pad ,
		_w35_
	);
	LUT3 #(
		.INIT('he8)
	) name26 (
		\3_pad ,
		\5_pad ,
		\6_pad ,
		_w36_
	);
	LUT2 #(
		.INIT('h2)
	) name27 (
		\2_pad ,
		\4_pad ,
		_w37_
	);
	LUT4 #(
		.INIT('h0109)
	) name28 (
		\2_pad ,
		\4_pad ,
		_w36_,
		_w28_,
		_w38_
	);
	LUT4 #(
		.INIT('h1337)
	) name29 (
		\3_pad ,
		\5_pad ,
		\7_pad ,
		\8_pad ,
		_w39_
	);
	LUT3 #(
		.INIT('h04)
	) name30 (
		_w35_,
		_w37_,
		_w39_,
		_w40_
	);
	LUT2 #(
		.INIT('h1)
	) name31 (
		_w38_,
		_w40_,
		_w41_
	);
	LUT2 #(
		.INIT('h4)
	) name32 (
		_w34_,
		_w41_,
		_w42_
	);
	LUT4 #(
		.INIT('h7277)
	) name33 (
		\4_pad ,
		\5_pad ,
		\7_pad ,
		\8_pad ,
		_w43_
	);
	LUT3 #(
		.INIT('h08)
	) name34 (
		\3_pad ,
		\4_pad ,
		\5_pad ,
		_w44_
	);
	LUT4 #(
		.INIT('hcc04)
	) name35 (
		\3_pad ,
		\6_pad ,
		_w43_,
		_w44_,
		_w45_
	);
	LUT3 #(
		.INIT('hc8)
	) name36 (
		\4_pad ,
		\6_pad ,
		\8_pad ,
		_w46_
	);
	LUT3 #(
		.INIT('h80)
	) name37 (
		\4_pad ,
		\7_pad ,
		\8_pad ,
		_w47_
	);
	LUT3 #(
		.INIT('he0)
	) name38 (
		\4_pad ,
		\6_pad ,
		\7_pad ,
		_w48_
	);
	LUT4 #(
		.INIT('hfe76)
	) name39 (
		\3_pad ,
		\5_pad ,
		_w47_,
		_w48_,
		_w49_
	);
	LUT4 #(
		.INIT('h5f4c)
	) name40 (
		\3_pad ,
		\4_pad ,
		\5_pad ,
		\6_pad ,
		_w50_
	);
	LUT2 #(
		.INIT('h8)
	) name41 (
		_w28_,
		_w50_,
		_w51_
	);
	LUT4 #(
		.INIT('h000e)
	) name42 (
		_w46_,
		_w49_,
		_w45_,
		_w51_,
		_w52_
	);
	LUT4 #(
		.INIT('h69a5)
	) name43 (
		\4_pad ,
		\5_pad ,
		\6_pad ,
		\7_pad ,
		_w53_
	);
	LUT4 #(
		.INIT('h5a65)
	) name44 (
		\4_pad ,
		\5_pad ,
		\6_pad ,
		\7_pad ,
		_w54_
	);
	LUT3 #(
		.INIT('h1b)
	) name45 (
		\8_pad ,
		_w53_,
		_w54_,
		_w55_
	);
	LUT4 #(
		.INIT('ha65a)
	) name46 (
		\5_pad ,
		\6_pad ,
		\7_pad ,
		\8_pad ,
		_w56_
	);
	LUT3 #(
		.INIT('h9a)
	) name47 (
		\6_pad ,
		\7_pad ,
		\8_pad ,
		_w57_
	);
	LUT2 #(
		.INIT('h6)
	) name48 (
		\7_pad ,
		\8_pad ,
		_w58_
	);
	assign \44_pad  = _w27_ ;
	assign \45_pad  = _w42_ ;
	assign \46_pad  = _w52_ ;
	assign \47_pad  = _w55_ ;
	assign \48_pad  = _w56_ ;
	assign \49_pad  = _w57_ ;
	assign \50_pad  = _w58_ ;
	assign \51_pad  = _w10_ ;
endmodule;